module real_aes_8183_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g524 ( .A1(n_0), .A2(n_171), .B(n_525), .C(n_528), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_1), .B(n_513), .Y(n_529) );
INVx1_ASAP7_75t_L g416 ( .A(n_2), .Y(n_416) );
INVx1_ASAP7_75t_L g189 ( .A(n_3), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_4), .B(n_160), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_5), .A2(n_428), .B(n_507), .Y(n_506) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_6), .A2(n_136), .B(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_7), .A2(n_35), .B1(n_116), .B2(n_125), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_8), .B(n_136), .Y(n_200) );
AND2x6_ASAP7_75t_L g134 ( .A(n_9), .B(n_135), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_10), .A2(n_134), .B(n_431), .C(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_11), .B(n_36), .Y(n_417) );
INVx1_ASAP7_75t_L g744 ( .A(n_11), .Y(n_744) );
INVx1_ASAP7_75t_L g132 ( .A(n_12), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_13), .B(n_123), .Y(n_143) );
INVx1_ASAP7_75t_L g181 ( .A(n_14), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_15), .B(n_160), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_16), .B(n_137), .Y(n_205) );
AO32x2_ASAP7_75t_L g168 ( .A1(n_17), .A2(n_133), .A3(n_136), .B1(n_169), .B2(n_173), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_18), .B(n_125), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_19), .B(n_137), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_20), .A2(n_51), .B1(n_116), .B2(n_125), .Y(n_172) );
AOI22xp33_ASAP7_75t_SL g122 ( .A1(n_21), .A2(n_79), .B1(n_123), .B2(n_125), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_22), .B(n_125), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_23), .A2(n_133), .B(n_431), .C(n_433), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_24), .A2(n_133), .B(n_431), .C(n_478), .Y(n_477) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_25), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_26), .B(n_128), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_27), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_28), .A2(n_428), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_29), .B(n_128), .Y(n_166) );
INVx2_ASAP7_75t_L g118 ( .A(n_30), .Y(n_118) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_31), .A2(n_452), .B(n_461), .C(n_463), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_32), .B(n_125), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_33), .B(n_128), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_34), .B(n_145), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_36), .B(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_37), .B(n_427), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_38), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_39), .B(n_160), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_40), .B(n_428), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_41), .A2(n_452), .B(n_461), .C(n_498), .Y(n_497) );
OAI22xp5_ASAP7_75t_SL g105 ( .A1(n_42), .A2(n_106), .B1(n_410), .B2(n_411), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_42), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_42), .A2(n_77), .B1(n_410), .B2(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_43), .B(n_125), .Y(n_195) );
INVx1_ASAP7_75t_L g526 ( .A(n_44), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_45), .A2(n_88), .B1(n_116), .B2(n_119), .Y(n_115) );
INVx1_ASAP7_75t_L g499 ( .A(n_46), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_47), .B(n_125), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_48), .B(n_125), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_49), .B(n_428), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_50), .B(n_187), .Y(n_199) );
AOI22xp33_ASAP7_75t_SL g209 ( .A1(n_52), .A2(n_56), .B1(n_123), .B2(n_125), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_53), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_54), .B(n_125), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_55), .B(n_125), .Y(n_224) );
INVx1_ASAP7_75t_L g135 ( .A(n_57), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_58), .B(n_428), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_59), .B(n_513), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_60), .A2(n_184), .B(n_187), .C(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_61), .B(n_125), .Y(n_190) );
INVx1_ASAP7_75t_L g131 ( .A(n_62), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_63), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_64), .B(n_160), .Y(n_465) );
AO32x2_ASAP7_75t_L g113 ( .A1(n_65), .A2(n_114), .A3(n_127), .B1(n_133), .B2(n_136), .Y(n_113) );
AOI22xp33_ASAP7_75t_SL g100 ( .A1(n_66), .A2(n_101), .B1(n_739), .B2(n_749), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_67), .B(n_126), .Y(n_489) );
INVx1_ASAP7_75t_L g223 ( .A(n_68), .Y(n_223) );
INVx1_ASAP7_75t_L g158 ( .A(n_69), .Y(n_158) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_70), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_71), .B(n_435), .Y(n_434) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_72), .A2(n_431), .B(n_448), .C(n_452), .Y(n_447) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_73), .A2(n_81), .B1(n_103), .B2(n_715), .C1(n_716), .C2(n_720), .Y(n_102) );
INVx1_ASAP7_75t_L g715 ( .A(n_73), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_74), .B(n_123), .Y(n_159) );
CKINVDCx16_ASAP7_75t_R g508 ( .A(n_75), .Y(n_508) );
INVx1_ASAP7_75t_L g748 ( .A(n_76), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_77), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_78), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_80), .B(n_116), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_82), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_83), .B(n_123), .Y(n_163) );
INVx2_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_85), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_86), .B(n_120), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_87), .B(n_123), .Y(n_196) );
OR2x2_ASAP7_75t_L g414 ( .A(n_89), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g714 ( .A(n_89), .Y(n_714) );
OR2x2_ASAP7_75t_L g732 ( .A(n_89), .B(n_719), .Y(n_732) );
NAND3xp33_ASAP7_75t_SL g745 ( .A(n_89), .B(n_416), .C(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_90), .A2(n_99), .B1(n_123), .B2(n_124), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_91), .B(n_428), .Y(n_459) );
INVx1_ASAP7_75t_L g464 ( .A(n_92), .Y(n_464) );
INVxp67_ASAP7_75t_L g511 ( .A(n_93), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_94), .B(n_123), .Y(n_221) );
INVx1_ASAP7_75t_L g449 ( .A(n_95), .Y(n_449) );
INVx1_ASAP7_75t_L g485 ( .A(n_96), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_97), .B(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g501 ( .A(n_98), .B(n_128), .Y(n_501) );
AOI22x1_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_724), .B1(n_733), .B2(n_734), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_412), .B1(n_418), .B2(n_711), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_105), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_720) );
INVx2_ASAP7_75t_L g411 ( .A(n_106), .Y(n_411) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
XOR2x2_ASAP7_75t_L g735 ( .A(n_107), .B(n_736), .Y(n_735) );
AND3x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_330), .C(n_378), .Y(n_107) );
NOR4xp25_ASAP7_75t_L g108 ( .A(n_109), .B(n_258), .C(n_303), .D(n_317), .Y(n_108) );
OAI311xp33_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_174), .A3(n_201), .B1(n_211), .C1(n_226), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_138), .Y(n_110) );
OAI21xp33_ASAP7_75t_L g211 ( .A1(n_111), .A2(n_212), .B(n_214), .Y(n_211) );
AND2x2_ASAP7_75t_L g319 ( .A(n_111), .B(n_246), .Y(n_319) );
AND2x2_ASAP7_75t_L g376 ( .A(n_111), .B(n_262), .Y(n_376) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g269 ( .A(n_112), .B(n_167), .Y(n_269) );
AND2x2_ASAP7_75t_L g326 ( .A(n_112), .B(n_274), .Y(n_326) );
INVx1_ASAP7_75t_L g367 ( .A(n_112), .Y(n_367) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_113), .Y(n_235) );
AND2x2_ASAP7_75t_L g276 ( .A(n_113), .B(n_167), .Y(n_276) );
AND2x2_ASAP7_75t_L g280 ( .A(n_113), .B(n_168), .Y(n_280) );
INVx1_ASAP7_75t_L g292 ( .A(n_113), .Y(n_292) );
OAI22xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_120), .B1(n_122), .B2(n_126), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g119 ( .A(n_117), .Y(n_119) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_117), .Y(n_125) );
AND2x6_ASAP7_75t_L g431 ( .A(n_117), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g124 ( .A(n_118), .Y(n_124) );
INVx1_ASAP7_75t_L g188 ( .A(n_118), .Y(n_188) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_119), .Y(n_466) );
INVx2_ASAP7_75t_L g528 ( .A(n_119), .Y(n_528) );
INVx2_ASAP7_75t_L g149 ( .A(n_120), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g169 ( .A1(n_120), .A2(n_170), .B1(n_171), .B2(n_172), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_120), .A2(n_171), .B1(n_208), .B2(n_209), .Y(n_207) );
INVx4_ASAP7_75t_L g527 ( .A(n_120), .Y(n_527) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g126 ( .A(n_121), .Y(n_126) );
INVx1_ASAP7_75t_L g145 ( .A(n_121), .Y(n_145) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_121), .Y(n_165) );
AND2x2_ASAP7_75t_L g429 ( .A(n_121), .B(n_188), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_121), .Y(n_432) );
INVx2_ASAP7_75t_L g182 ( .A(n_123), .Y(n_182) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx3_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_125), .Y(n_451) );
INVx5_ASAP7_75t_L g160 ( .A(n_126), .Y(n_160) );
INVx1_ASAP7_75t_L g438 ( .A(n_127), .Y(n_438) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_128), .A2(n_140), .B(n_150), .Y(n_139) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_128), .A2(n_155), .B(n_166), .Y(n_154) );
INVx1_ASAP7_75t_L g441 ( .A(n_128), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_128), .A2(n_459), .B(n_460), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_128), .A2(n_496), .B(n_497), .Y(n_495) );
AND2x2_ASAP7_75t_SL g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_L g137 ( .A(n_129), .B(n_130), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
NAND3xp33_ASAP7_75t_L g206 ( .A(n_133), .B(n_207), .C(n_210), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_133), .A2(n_219), .B(n_222), .Y(n_218) );
BUFx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_134), .A2(n_141), .B(n_146), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g155 ( .A1(n_134), .A2(n_156), .B(n_161), .Y(n_155) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_134), .A2(n_180), .B(n_185), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g193 ( .A1(n_134), .A2(n_194), .B(n_197), .Y(n_193) );
AND2x4_ASAP7_75t_L g428 ( .A(n_134), .B(n_429), .Y(n_428) );
INVx4_ASAP7_75t_SL g453 ( .A(n_134), .Y(n_453) );
NAND2x1p5_ASAP7_75t_L g486 ( .A(n_134), .B(n_429), .Y(n_486) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_136), .A2(n_193), .B(n_200), .Y(n_192) );
INVx4_ASAP7_75t_L g210 ( .A(n_136), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_136), .A2(n_476), .B(n_477), .Y(n_475) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_136), .Y(n_505) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g173 ( .A(n_137), .Y(n_173) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_151), .Y(n_138) );
AND2x2_ASAP7_75t_L g213 ( .A(n_139), .B(n_167), .Y(n_213) );
INVx2_ASAP7_75t_L g247 ( .A(n_139), .Y(n_247) );
AND2x2_ASAP7_75t_L g262 ( .A(n_139), .B(n_168), .Y(n_262) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_139), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_139), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g282 ( .A(n_139), .B(n_245), .Y(n_282) );
INVx1_ASAP7_75t_L g294 ( .A(n_139), .Y(n_294) );
INVx1_ASAP7_75t_L g335 ( .A(n_139), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_139), .B(n_235), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_149), .Y(n_146) );
O2A1O1Ixp5_ASAP7_75t_L g222 ( .A1(n_149), .A2(n_186), .B(n_223), .C(n_224), .Y(n_222) );
NOR2xp67_ASAP7_75t_L g151 ( .A(n_152), .B(n_167), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g212 ( .A(n_153), .B(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_153), .Y(n_240) );
AND2x2_ASAP7_75t_SL g293 ( .A(n_153), .B(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g297 ( .A(n_153), .B(n_167), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_153), .B(n_292), .Y(n_355) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g245 ( .A(n_154), .Y(n_245) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_154), .Y(n_261) );
OR2x2_ASAP7_75t_L g334 ( .A(n_154), .B(n_335), .Y(n_334) );
O2A1O1Ixp5_ASAP7_75t_SL g156 ( .A1(n_157), .A2(n_158), .B(n_159), .C(n_160), .Y(n_156) );
INVx2_ASAP7_75t_L g171 ( .A(n_160), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_160), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_160), .A2(n_220), .B(n_221), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_160), .B(n_511), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_164), .Y(n_161) );
INVx1_ASAP7_75t_L g184 ( .A(n_164), .Y(n_184) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g435 ( .A(n_165), .Y(n_435) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx2_ASAP7_75t_L g241 ( .A(n_168), .Y(n_241) );
AND2x2_ASAP7_75t_L g246 ( .A(n_168), .B(n_247), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_171), .A2(n_186), .B(n_189), .C(n_190), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_171), .A2(n_198), .B(n_199), .Y(n_197) );
INVx2_ASAP7_75t_L g178 ( .A(n_173), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_173), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_174), .B(n_229), .Y(n_392) );
INVx1_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
OR2x2_ASAP7_75t_L g362 ( .A(n_175), .B(n_203), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_192), .Y(n_175) );
AND2x2_ASAP7_75t_L g238 ( .A(n_176), .B(n_229), .Y(n_238) );
INVx2_ASAP7_75t_L g250 ( .A(n_176), .Y(n_250) );
AND2x2_ASAP7_75t_L g284 ( .A(n_176), .B(n_232), .Y(n_284) );
AND2x2_ASAP7_75t_L g351 ( .A(n_176), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_177), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g231 ( .A(n_177), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g271 ( .A(n_177), .B(n_192), .Y(n_271) );
AND2x2_ASAP7_75t_L g288 ( .A(n_177), .B(n_289), .Y(n_288) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_191), .Y(n_177) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_178), .A2(n_218), .B(n_225), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_183), .C(n_184), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_182), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_182), .A2(n_489), .B(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_184), .A2(n_449), .B(n_450), .C(n_451), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_186), .A2(n_434), .B(n_436), .Y(n_433) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g214 ( .A(n_192), .B(n_215), .Y(n_214) );
INVx3_ASAP7_75t_L g232 ( .A(n_192), .Y(n_232) );
AND2x2_ASAP7_75t_L g237 ( .A(n_192), .B(n_217), .Y(n_237) );
AND2x2_ASAP7_75t_L g310 ( .A(n_192), .B(n_289), .Y(n_310) );
AND2x2_ASAP7_75t_L g375 ( .A(n_192), .B(n_365), .Y(n_375) );
OAI311xp33_ASAP7_75t_L g258 ( .A1(n_201), .A2(n_259), .A3(n_263), .B1(n_265), .C1(n_285), .Y(n_258) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g270 ( .A(n_202), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g329 ( .A(n_202), .B(n_237), .Y(n_329) );
AND2x2_ASAP7_75t_L g403 ( .A(n_202), .B(n_284), .Y(n_403) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_203), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g338 ( .A(n_203), .Y(n_338) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g229 ( .A(n_204), .Y(n_229) );
NOR2x1_ASAP7_75t_L g301 ( .A(n_204), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g358 ( .A(n_204), .B(n_232), .Y(n_358) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
INVx1_ASAP7_75t_L g255 ( .A(n_205), .Y(n_255) );
AO21x1_ASAP7_75t_L g254 ( .A1(n_207), .A2(n_210), .B(n_255), .Y(n_254) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_210), .A2(n_446), .B(n_455), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_210), .B(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_210), .B(n_468), .Y(n_467) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_210), .A2(n_484), .B(n_491), .Y(n_483) );
INVx3_ASAP7_75t_L g513 ( .A(n_210), .Y(n_513) );
AND2x2_ASAP7_75t_L g233 ( .A(n_213), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g286 ( .A(n_213), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g366 ( .A(n_213), .B(n_367), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g265 ( .A1(n_214), .A2(n_246), .B1(n_266), .B2(n_270), .C(n_272), .Y(n_265) );
INVx1_ASAP7_75t_L g390 ( .A(n_215), .Y(n_390) );
OR2x2_ASAP7_75t_L g356 ( .A(n_216), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g251 ( .A(n_217), .B(n_232), .Y(n_251) );
OR2x2_ASAP7_75t_L g253 ( .A(n_217), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g278 ( .A(n_217), .Y(n_278) );
INVx2_ASAP7_75t_L g289 ( .A(n_217), .Y(n_289) );
AND2x2_ASAP7_75t_L g316 ( .A(n_217), .B(n_254), .Y(n_316) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_217), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_233), .B1(n_236), .B2(n_239), .C(n_242), .Y(n_226) );
INVx1_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
AND2x2_ASAP7_75t_L g327 ( .A(n_229), .B(n_237), .Y(n_327) );
AND2x2_ASAP7_75t_L g377 ( .A(n_229), .B(n_231), .Y(n_377) );
INVx2_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g264 ( .A(n_231), .B(n_235), .Y(n_264) );
AND2x2_ASAP7_75t_L g343 ( .A(n_231), .B(n_316), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_232), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g302 ( .A(n_232), .Y(n_302) );
OAI21xp33_ASAP7_75t_L g312 ( .A1(n_233), .A2(n_313), .B(n_315), .Y(n_312) );
OR2x2_ASAP7_75t_L g256 ( .A(n_234), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g322 ( .A(n_234), .B(n_282), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_234), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g299 ( .A(n_235), .B(n_268), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_235), .B(n_382), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_236), .B(n_262), .Y(n_372) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
AND2x2_ASAP7_75t_L g295 ( .A(n_237), .B(n_250), .Y(n_295) );
INVx1_ASAP7_75t_L g311 ( .A(n_238), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_248), .B1(n_252), .B2(n_256), .Y(n_242) );
INVx2_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g274 ( .A(n_245), .Y(n_274) );
INVx1_ASAP7_75t_L g287 ( .A(n_245), .Y(n_287) );
INVx1_ASAP7_75t_L g257 ( .A(n_246), .Y(n_257) );
AND2x2_ASAP7_75t_L g328 ( .A(n_246), .B(n_274), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_246), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
OR2x2_ASAP7_75t_L g252 ( .A(n_249), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_249), .B(n_365), .Y(n_364) );
NOR2xp67_ASAP7_75t_L g396 ( .A(n_249), .B(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g399 ( .A(n_251), .B(n_351), .Y(n_399) );
INVx1_ASAP7_75t_SL g365 ( .A(n_253), .Y(n_365) );
AND2x2_ASAP7_75t_L g305 ( .A(n_254), .B(n_289), .Y(n_305) );
INVx1_ASAP7_75t_L g352 ( .A(n_254), .Y(n_352) );
OAI222xp33_ASAP7_75t_L g393 ( .A1(n_259), .A2(n_349), .B1(n_394), .B2(n_395), .C1(n_398), .C2(n_400), .Y(n_393) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g314 ( .A(n_261), .Y(n_314) );
AND2x2_ASAP7_75t_L g325 ( .A(n_262), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_262), .B(n_367), .Y(n_394) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_264), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g369 ( .A(n_266), .Y(n_369) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_SL g307 ( .A(n_269), .Y(n_307) );
AND2x2_ASAP7_75t_L g386 ( .A(n_269), .B(n_347), .Y(n_386) );
AND2x2_ASAP7_75t_L g409 ( .A(n_269), .B(n_293), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_271), .B(n_305), .Y(n_304) );
OAI32xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_275), .A3(n_277), .B1(n_279), .B2(n_283), .Y(n_272) );
BUFx2_ASAP7_75t_L g347 ( .A(n_274), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_275), .B(n_293), .Y(n_374) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g313 ( .A(n_276), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g381 ( .A(n_276), .B(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g370 ( .A(n_277), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AND2x2_ASAP7_75t_L g341 ( .A(n_280), .B(n_314), .Y(n_341) );
INVx2_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
OAI221xp5_ASAP7_75t_SL g303 ( .A1(n_282), .A2(n_304), .B1(n_306), .B2(n_308), .C(n_312), .Y(n_303) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g315 ( .A(n_284), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g321 ( .A(n_284), .B(n_305), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_288), .B1(n_290), .B2(n_295), .C(n_296), .Y(n_285) );
INVx1_ASAP7_75t_L g404 ( .A(n_286), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_287), .B(n_381), .Y(n_380) );
NAND2x1p5_ASAP7_75t_L g300 ( .A(n_288), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_293), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g359 ( .A(n_293), .Y(n_359) );
BUFx3_ASAP7_75t_L g382 ( .A(n_294), .Y(n_382) );
INVx1_ASAP7_75t_SL g323 ( .A(n_295), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_295), .B(n_337), .Y(n_336) );
AOI21xp33_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_298), .B(n_300), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_297), .A2(n_398), .B1(n_402), .B2(n_404), .C(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g344 ( .A(n_302), .B(n_305), .Y(n_344) );
INVx1_ASAP7_75t_L g408 ( .A(n_302), .Y(n_408) );
INVx2_ASAP7_75t_L g397 ( .A(n_305), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_305), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g350 ( .A(n_310), .B(n_351), .Y(n_350) );
OAI221xp5_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_320), .B1(n_322), .B2(n_323), .C(n_324), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B1(n_328), .B2(n_329), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_326), .A2(n_388), .B1(n_389), .B2(n_391), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g405 ( .A1(n_329), .A2(n_406), .B(n_409), .Y(n_405) );
NOR4xp25_ASAP7_75t_SL g330 ( .A(n_331), .B(n_339), .C(n_348), .D(n_368), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_336), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B1(n_345), .B2(n_346), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g384 ( .A(n_344), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_353), .B1(n_356), .B2(n_359), .C(n_360), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g371 ( .A(n_351), .Y(n_371) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI21xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_363), .B(n_366), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI211xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B(n_372), .C(n_373), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_376), .B2(n_377), .Y(n_373) );
CKINVDCx14_ASAP7_75t_R g383 ( .A(n_377), .Y(n_383) );
NOR3xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_393), .C(n_401), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B1(n_384), .B2(n_385), .C(n_387), .Y(n_379) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g721 ( .A(n_413), .Y(n_721) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g713 ( .A(n_415), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g719 ( .A(n_415), .Y(n_719) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g722 ( .A(n_419), .Y(n_722) );
AND3x1_ASAP7_75t_L g419 ( .A(n_420), .B(n_615), .C(n_672), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_560), .C(n_596), .Y(n_420) );
OAI211xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_469), .B(n_515), .C(n_547), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_442), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g518 ( .A(n_424), .B(n_519), .Y(n_518) );
INVx5_ASAP7_75t_L g546 ( .A(n_424), .Y(n_546) );
AND2x2_ASAP7_75t_L g619 ( .A(n_424), .B(n_535), .Y(n_619) );
AND2x2_ASAP7_75t_L g657 ( .A(n_424), .B(n_563), .Y(n_657) );
AND2x2_ASAP7_75t_L g677 ( .A(n_424), .B(n_520), .Y(n_677) );
OR2x6_ASAP7_75t_L g424 ( .A(n_425), .B(n_439), .Y(n_424) );
AOI21xp5_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_430), .B(n_438), .Y(n_425) );
BUFx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx5_ASAP7_75t_L g462 ( .A(n_431), .Y(n_462) );
INVx2_ASAP7_75t_L g437 ( .A(n_435), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_437), .A2(n_464), .B(n_465), .C(n_466), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_437), .A2(n_466), .B(n_499), .C(n_500), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_442), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_457), .Y(n_442) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_443), .Y(n_558) );
AND2x2_ASAP7_75t_L g572 ( .A(n_443), .B(n_519), .Y(n_572) );
INVx1_ASAP7_75t_L g595 ( .A(n_443), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_443), .B(n_546), .Y(n_634) );
OR2x2_ASAP7_75t_L g671 ( .A(n_443), .B(n_517), .Y(n_671) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_444), .Y(n_607) );
AND2x2_ASAP7_75t_L g614 ( .A(n_444), .B(n_520), .Y(n_614) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g535 ( .A(n_445), .B(n_520), .Y(n_535) );
BUFx2_ASAP7_75t_L g563 ( .A(n_445), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_454), .Y(n_446) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_453), .A2(n_462), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_453), .A2(n_462), .B(n_523), .C(n_524), .Y(n_522) );
INVx5_ASAP7_75t_L g517 ( .A(n_457), .Y(n_517) );
BUFx2_ASAP7_75t_L g539 ( .A(n_457), .Y(n_539) );
AND2x2_ASAP7_75t_L g696 ( .A(n_457), .B(n_550), .Y(n_696) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_467), .Y(n_457) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_502), .Y(n_470) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_471), .A2(n_597), .B1(n_604), .B2(n_605), .C(n_608), .Y(n_596) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
AND2x2_ASAP7_75t_L g503 ( .A(n_472), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_472), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g531 ( .A(n_473), .B(n_482), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_473), .B(n_483), .Y(n_541) );
OR2x2_ASAP7_75t_L g552 ( .A(n_473), .B(n_504), .Y(n_552) );
AND2x2_ASAP7_75t_L g555 ( .A(n_473), .B(n_543), .Y(n_555) );
AND2x2_ASAP7_75t_L g571 ( .A(n_473), .B(n_493), .Y(n_571) );
OR2x2_ASAP7_75t_L g587 ( .A(n_473), .B(n_483), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_473), .B(n_504), .Y(n_649) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_474), .B(n_493), .Y(n_641) );
AND2x2_ASAP7_75t_L g644 ( .A(n_474), .B(n_483), .Y(n_644) );
OR2x2_ASAP7_75t_L g565 ( .A(n_481), .B(n_552), .Y(n_565) );
INVx2_ASAP7_75t_L g591 ( .A(n_481), .Y(n_591) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_493), .Y(n_481) );
AND2x2_ASAP7_75t_L g514 ( .A(n_482), .B(n_494), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_482), .B(n_504), .Y(n_570) );
OR2x2_ASAP7_75t_L g581 ( .A(n_482), .B(n_494), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_482), .B(n_543), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_482), .A2(n_674), .B1(n_676), .B2(n_678), .C(n_681), .Y(n_673) );
INVx5_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_483), .B(n_504), .Y(n_612) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_487), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_493), .B(n_543), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_493), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g559 ( .A(n_493), .B(n_531), .Y(n_559) );
OR2x2_ASAP7_75t_L g603 ( .A(n_493), .B(n_504), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_493), .B(n_555), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_493), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g668 ( .A(n_493), .B(n_669), .Y(n_668) );
INVx5_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_SL g532 ( .A(n_494), .B(n_503), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_SL g536 ( .A1(n_494), .A2(n_537), .B(n_540), .C(n_544), .Y(n_536) );
OR2x2_ASAP7_75t_L g574 ( .A(n_494), .B(n_570), .Y(n_574) );
OR2x2_ASAP7_75t_L g610 ( .A(n_494), .B(n_552), .Y(n_610) );
OAI311xp33_ASAP7_75t_L g616 ( .A1(n_494), .A2(n_555), .A3(n_617), .B1(n_620), .C1(n_627), .Y(n_616) );
AND2x2_ASAP7_75t_L g667 ( .A(n_494), .B(n_504), .Y(n_667) );
AND2x2_ASAP7_75t_L g675 ( .A(n_494), .B(n_530), .Y(n_675) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_494), .Y(n_693) );
AND2x2_ASAP7_75t_L g710 ( .A(n_494), .B(n_531), .Y(n_710) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_501), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_514), .Y(n_502) );
AND2x2_ASAP7_75t_L g538 ( .A(n_503), .B(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g694 ( .A(n_503), .Y(n_694) );
AND2x2_ASAP7_75t_L g530 ( .A(n_504), .B(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g543 ( .A(n_504), .Y(n_543) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_504), .Y(n_586) );
INVxp67_ASAP7_75t_L g625 ( .A(n_504), .Y(n_625) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B(n_512), .Y(n_504) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_513), .A2(n_521), .B(n_529), .Y(n_520) );
AND2x2_ASAP7_75t_L g703 ( .A(n_514), .B(n_551), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_530), .B1(n_532), .B2(n_533), .C(n_536), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_517), .B(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g556 ( .A(n_517), .B(n_546), .Y(n_556) );
AND2x2_ASAP7_75t_L g564 ( .A(n_517), .B(n_519), .Y(n_564) );
OR2x2_ASAP7_75t_L g576 ( .A(n_517), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g594 ( .A(n_517), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g618 ( .A(n_517), .B(n_619), .Y(n_618) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_517), .Y(n_638) );
AND2x2_ASAP7_75t_L g690 ( .A(n_517), .B(n_614), .Y(n_690) );
OAI31xp33_ASAP7_75t_L g698 ( .A1(n_517), .A2(n_567), .A3(n_666), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_518), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_SL g662 ( .A(n_518), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_518), .B(n_671), .Y(n_670) );
AND2x4_ASAP7_75t_L g550 ( .A(n_519), .B(n_546), .Y(n_550) );
INVx1_ASAP7_75t_L g637 ( .A(n_519), .Y(n_637) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g687 ( .A(n_520), .B(n_546), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_SL g697 ( .A(n_530), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_531), .B(n_602), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_532), .A2(n_644), .B1(n_682), .B2(n_685), .Y(n_681) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g545 ( .A(n_535), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g604 ( .A(n_535), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_535), .B(n_556), .Y(n_709) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g679 ( .A(n_538), .B(n_680), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_539), .A2(n_598), .B(n_600), .Y(n_597) );
OR2x2_ASAP7_75t_L g605 ( .A(n_539), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g626 ( .A(n_539), .B(n_614), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_539), .B(n_637), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_539), .B(n_677), .Y(n_676) );
OAI221xp5_ASAP7_75t_SL g653 ( .A1(n_540), .A2(n_654), .B1(n_659), .B2(n_662), .C(n_663), .Y(n_653) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
OR2x2_ASAP7_75t_L g630 ( .A(n_541), .B(n_603), .Y(n_630) );
INVx1_ASAP7_75t_L g669 ( .A(n_541), .Y(n_669) );
INVx2_ASAP7_75t_L g645 ( .A(n_542), .Y(n_645) );
INVx1_ASAP7_75t_L g579 ( .A(n_543), .Y(n_579) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g584 ( .A(n_546), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_546), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g613 ( .A(n_546), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g701 ( .A(n_546), .B(n_671), .Y(n_701) );
AOI222xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_551), .B1(n_553), .B2(n_556), .C1(n_557), .C2(n_559), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g557 ( .A(n_550), .B(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_550), .A2(n_600), .B1(n_628), .B2(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_550), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
OAI21xp33_ASAP7_75t_SL g588 ( .A1(n_559), .A2(n_589), .B(n_592), .Y(n_588) );
OAI211xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_565), .B(n_566), .C(n_588), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
AOI221xp5_ASAP7_75t_L g566 ( .A1(n_564), .A2(n_567), .B1(n_572), .B2(n_573), .C(n_575), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_564), .B(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_L g658 ( .A(n_564), .Y(n_658) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
AND2x2_ASAP7_75t_L g660 ( .A(n_569), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g577 ( .A(n_572), .Y(n_577) );
AND2x2_ASAP7_75t_L g583 ( .A(n_572), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_578), .B1(n_582), .B2(n_585), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_579), .B(n_591), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_580), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g680 ( .A(n_584), .Y(n_680) );
AND2x2_ASAP7_75t_L g699 ( .A(n_584), .B(n_614), .Y(n_699) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_591), .B(n_648), .Y(n_707) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_594), .B(n_662), .Y(n_705) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g628 ( .A(n_606), .Y(n_628) );
BUFx2_ASAP7_75t_L g652 ( .A(n_607), .Y(n_652) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_611), .B(n_613), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR3xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_631), .C(n_653), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .B(n_626), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_635), .B(n_639), .C(n_642), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_632), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR2xp67_ASAP7_75t_SL g636 ( .A(n_637), .B(n_638), .Y(n_636) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_SL g661 ( .A(n_641), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B(n_650), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
AND2x2_ASAP7_75t_L g666 ( .A(n_644), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B1(n_668), .B2(n_670), .Y(n_663) );
INVx2_ASAP7_75t_SL g684 ( .A(n_671), .Y(n_684) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_688), .C(n_700), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_684), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B1(n_695), .B2(n_697), .C(n_698), .Y(n_688) );
A2O1A1Ixp33_ASAP7_75t_L g700 ( .A1(n_689), .A2(n_701), .B(n_702), .C(n_704), .Y(n_700) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_708), .B2(n_710), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g723 ( .A(n_712), .Y(n_723) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NOR2x2_ASAP7_75t_L g718 ( .A(n_714), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx3_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_729), .Y(n_724) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
BUFx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g733 ( .A(n_727), .Y(n_733) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_729), .A2(n_735), .B(n_738), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_732), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx5_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
CKINVDCx9p33_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_742), .Y(n_750) );
OR2x4_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .Y(n_742) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
endmodule