module fake_jpeg_16119_n_22 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_22);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_22;

wire n_13;
wire n_21;
wire n_10;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;

AOI22xp5_ASAP7_75t_L g8 ( 
.A1(n_4),
.A2(n_6),
.B1(n_5),
.B2(n_7),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_2),
.B(n_3),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_11),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_17),
.C(n_18),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_12),
.B1(n_8),
.B2(n_15),
.Y(n_19)
);

AOI321xp33_ASAP7_75t_L g21 ( 
.A1(n_20),
.A2(n_19),
.A3(n_10),
.B1(n_14),
.B2(n_13),
.C(n_17),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_21),
.A2(n_13),
.B(n_19),
.Y(n_22)
);


endmodule