module fake_jpeg_27772_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx6_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_24),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_23),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_14),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_1),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_10),
.B1(n_8),
.B2(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_13),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_30),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_21),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_11),
.Y(n_37)
);

OA21x2_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_8),
.B(n_17),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_40),
.B1(n_13),
.B2(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

OAI321xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_34),
.A3(n_35),
.B1(n_36),
.B2(n_33),
.C(n_3),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_43),
.B1(n_33),
.B2(n_41),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_47),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_5),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_50),
.A2(n_51),
.B(n_49),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_5),
.Y(n_54)
);


endmodule