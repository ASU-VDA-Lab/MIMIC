module fake_jpeg_1109_n_658 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_658);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_658;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_312;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_576;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g208 ( 
.A(n_59),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_61),
.Y(n_163)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_64),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_23),
.B(n_0),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_65),
.A2(n_109),
.B(n_118),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_66),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_67),
.Y(n_175)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_68),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_69),
.Y(n_178)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_72),
.Y(n_212)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_75),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_80),
.Y(n_188)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_82),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_83),
.B(n_111),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_84),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_85),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_88),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_90),
.Y(n_201)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_96),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_97),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_23),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_101),
.Y(n_143)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_20),
.B(n_1),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx11_ASAP7_75t_SL g104 ( 
.A(n_54),
.Y(n_104)
);

INVx5_ASAP7_75t_SL g182 ( 
.A(n_104),
.Y(n_182)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx11_ASAP7_75t_SL g106 ( 
.A(n_19),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_108),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_20),
.B(n_2),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_31),
.Y(n_112)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_25),
.Y(n_114)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_51),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_116),
.B(n_120),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_30),
.B(n_2),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_30),
.B(n_18),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_25),
.Y(n_122)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_26),
.Y(n_123)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_44),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_44),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_44),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g161 ( 
.A(n_126),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_46),
.Y(n_127)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_46),
.Y(n_128)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_26),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_129),
.B(n_57),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_61),
.A2(n_21),
.B1(n_52),
.B2(n_50),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_134),
.A2(n_21),
.B1(n_50),
.B2(n_52),
.Y(n_226)
);

BUFx12f_ASAP7_75t_SL g136 ( 
.A(n_104),
.Y(n_136)
);

INVx6_ASAP7_75t_SL g244 ( 
.A(n_136),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_109),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_150),
.B(n_165),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_65),
.B(n_55),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_156),
.B(n_36),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_128),
.B(n_55),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_173),
.B(n_52),
.Y(n_269)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_76),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_179),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_115),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_180),
.B(n_196),
.Y(n_279)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_66),
.Y(n_185)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_67),
.Y(n_189)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_59),
.Y(n_193)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_193),
.Y(n_259)
);

HAxp5_ASAP7_75t_SL g196 ( 
.A(n_108),
.B(n_57),
.CON(n_196),
.SN(n_196)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_198),
.Y(n_300)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_69),
.Y(n_204)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_75),
.Y(n_207)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_59),
.Y(n_209)
);

BUFx2_ASAP7_75t_SL g254 ( 
.A(n_209),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_40),
.Y(n_245)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_88),
.Y(n_214)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_214),
.Y(n_290)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_77),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_80),
.Y(n_216)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_216),
.Y(n_267)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_88),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_82),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_84),
.Y(n_221)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_221),
.Y(n_273)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_85),
.Y(n_222)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_222),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_173),
.A2(n_21),
.B(n_58),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_223),
.A2(n_155),
.B(n_168),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_150),
.A2(n_36),
.B1(n_34),
.B2(n_33),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_225),
.A2(n_287),
.B1(n_240),
.B2(n_298),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_226),
.A2(n_274),
.B1(n_278),
.B2(n_238),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_228),
.B(n_233),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_46),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_229),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_165),
.A2(n_40),
.B1(n_53),
.B2(n_58),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_231),
.A2(n_288),
.B1(n_292),
.B2(n_297),
.Y(n_313)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_232),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_161),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_58),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_238),
.Y(n_338)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_130),
.Y(n_239)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_239),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

BUFx16f_ASAP7_75t_L g243 ( 
.A(n_137),
.Y(n_243)
);

BUFx24_ASAP7_75t_L g322 ( 
.A(n_243),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_245),
.B(n_246),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_143),
.B(n_53),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_195),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_247),
.B(n_249),
.Y(n_321)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_248),
.Y(n_332)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_195),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_176),
.B(n_119),
.C(n_126),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_250),
.B(n_261),
.C(n_283),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_200),
.A2(n_86),
.B1(n_110),
.B2(n_103),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_253),
.A2(n_168),
.B1(n_178),
.B2(n_175),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_171),
.B(n_50),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_255),
.B(n_275),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_180),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_256),
.B(n_258),
.Y(n_336)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_169),
.Y(n_257)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_177),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_210),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_260),
.B(n_264),
.Y(n_342)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_157),
.B(n_96),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_171),
.B(n_200),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_135),
.B(n_47),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_174),
.B(n_56),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_197),
.B(n_47),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_265),
.Y(n_346)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_137),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_163),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_268),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_269),
.B(n_271),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_194),
.B(n_90),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_270),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_182),
.B(n_56),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_134),
.A2(n_89),
.B1(n_87),
.B2(n_42),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_131),
.B(n_42),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_158),
.B(n_34),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_276),
.B(n_281),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_152),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_277),
.B(n_208),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_140),
.A2(n_33),
.B1(n_32),
.B2(n_119),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_141),
.Y(n_280)
);

BUFx2_ASAP7_75t_SL g347 ( 
.A(n_280),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_146),
.B(n_32),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g283 ( 
.A(n_160),
.B(n_2),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_147),
.Y(n_284)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_172),
.Y(n_286)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_286),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_139),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_154),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_138),
.Y(n_289)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_289),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_151),
.B(n_3),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_291),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_154),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_141),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_293),
.Y(n_333)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_166),
.Y(n_294)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_294),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_170),
.B(n_6),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_295),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_142),
.B(n_9),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_296),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_212),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_172),
.Y(n_298)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_298),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_144),
.Y(n_299)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_188),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_301),
.Y(n_356)
);

OA22x2_ASAP7_75t_L g302 ( 
.A1(n_223),
.A2(n_133),
.B1(n_164),
.B2(n_183),
.Y(n_302)
);

OA22x2_ASAP7_75t_L g377 ( 
.A1(n_302),
.A2(n_323),
.B1(n_232),
.B2(n_239),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_303),
.B(n_307),
.Y(n_402)
);

AO22x1_ASAP7_75t_L g307 ( 
.A1(n_229),
.A2(n_196),
.B1(n_212),
.B2(n_206),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_308),
.B(n_324),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_255),
.A2(n_162),
.B1(n_184),
.B2(n_211),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_314),
.A2(n_317),
.B1(n_320),
.B2(n_337),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_242),
.A2(n_145),
.B(n_149),
.C(n_148),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_315),
.B(n_361),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_279),
.A2(n_132),
.B1(n_201),
.B2(n_205),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_279),
.A2(n_220),
.B1(n_203),
.B2(n_218),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_275),
.A2(n_159),
.B1(n_186),
.B2(n_152),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_178),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_350),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_244),
.A2(n_190),
.B1(n_167),
.B2(n_147),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_335),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_250),
.A2(n_218),
.B1(n_175),
.B2(n_153),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_238),
.A2(n_202),
.B1(n_208),
.B2(n_167),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_345),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_348),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_283),
.B(n_261),
.Y(n_350)
);

O2A1O1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_244),
.A2(n_202),
.B(n_14),
.C(n_15),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_351),
.A2(n_355),
.B(n_308),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_252),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_352),
.A2(n_254),
.B1(n_230),
.B2(n_266),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_261),
.A2(n_10),
.B1(n_16),
.B2(n_17),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_353),
.A2(n_354),
.B1(n_357),
.B2(n_358),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_270),
.A2(n_229),
.B1(n_301),
.B2(n_257),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_224),
.A2(n_10),
.B(n_16),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_270),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_252),
.A2(n_294),
.B1(n_235),
.B2(n_234),
.Y(n_358)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_347),
.Y(n_362)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_362),
.Y(n_423)
);

INVx13_ASAP7_75t_L g364 ( 
.A(n_322),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_364),
.Y(n_428)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_326),
.Y(n_367)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_367),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_329),
.A2(n_241),
.B1(n_300),
.B2(n_227),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_368),
.A2(n_379),
.B1(n_386),
.B2(n_388),
.Y(n_421)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_326),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_378),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_272),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_370),
.B(n_375),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_305),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_371),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_331),
.B(n_227),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_374),
.Y(n_409)
);

AND2x2_ASAP7_75t_SL g373 ( 
.A(n_350),
.B(n_273),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_373),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_282),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_290),
.C(n_273),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_267),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_376),
.B(n_393),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g413 ( 
.A1(n_377),
.A2(n_307),
.B(n_302),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_358),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_267),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_401),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_303),
.A2(n_241),
.B1(n_236),
.B2(n_237),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_382),
.A2(n_391),
.B1(n_394),
.B2(n_399),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_383),
.Y(n_446)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_384),
.B(n_387),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_317),
.A2(n_248),
.B1(n_300),
.B2(n_289),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_314),
.A2(n_236),
.B1(n_237),
.B2(n_251),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_309),
.A2(n_299),
.B1(n_284),
.B2(n_290),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_390),
.A2(n_397),
.B(n_345),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_323),
.A2(n_282),
.B1(n_251),
.B2(n_286),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_332),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_392),
.B(n_395),
.Y(n_432)
);

AND2x6_ASAP7_75t_L g393 ( 
.A(n_342),
.B(n_243),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_338),
.A2(n_268),
.B1(n_230),
.B2(n_259),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_327),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_346),
.B(n_285),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_396),
.B(n_403),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_320),
.A2(n_259),
.B1(n_266),
.B2(n_285),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_338),
.A2(n_243),
.B1(n_316),
.B2(n_344),
.Y(n_399)
);

AND2x6_ASAP7_75t_L g400 ( 
.A(n_342),
.B(n_360),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_400),
.B(n_404),
.Y(n_435)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_319),
.B(n_334),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_336),
.B(n_311),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_328),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_302),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_334),
.B(n_344),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_408),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_411),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_SL g467 ( 
.A1(n_413),
.A2(n_426),
.B(n_443),
.C(n_377),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_402),
.A2(n_324),
.B1(n_313),
.B2(n_316),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_416),
.A2(n_418),
.B1(n_425),
.B2(n_430),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_402),
.A2(n_360),
.B1(n_330),
.B2(n_302),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_381),
.A2(n_355),
.B(n_307),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_419),
.A2(n_420),
.B(n_424),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_381),
.A2(n_406),
.B(n_402),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_407),
.A2(n_390),
.B(n_398),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_366),
.A2(n_384),
.B1(n_378),
.B2(n_385),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_366),
.A2(n_330),
.B1(n_302),
.B2(n_359),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_374),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_433),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_380),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_385),
.A2(n_337),
.B1(n_321),
.B2(n_356),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_434),
.A2(n_438),
.B1(n_441),
.B2(n_372),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_363),
.A2(n_359),
.B1(n_336),
.B2(n_321),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_437),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_383),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_370),
.A2(n_356),
.B1(n_311),
.B2(n_357),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_382),
.A2(n_353),
.B1(n_315),
.B2(n_340),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_373),
.A2(n_340),
.B1(n_310),
.B2(n_343),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_364),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_348),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_407),
.A2(n_351),
.B(n_341),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_447),
.A2(n_389),
.B(n_398),
.Y(n_450)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_410),
.Y(n_448)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_448),
.Y(n_485)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_410),
.Y(n_449)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_449),
.Y(n_501)
);

A2O1A1Ixp33_ASAP7_75t_L g502 ( 
.A1(n_450),
.A2(n_475),
.B(n_416),
.C(n_447),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_420),
.A2(n_399),
.B(n_393),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_451),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_428),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_453),
.B(n_461),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_420),
.B(n_377),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_454),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_412),
.B(n_404),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_455),
.B(n_460),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_432),
.Y(n_456)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_456),
.Y(n_510)
);

CKINVDCx12_ASAP7_75t_R g458 ( 
.A(n_412),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_458),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_432),
.Y(n_459)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_459),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_417),
.B(n_304),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_445),
.Y(n_461)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_417),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_463),
.B(n_473),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_439),
.B(n_376),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_464),
.B(n_479),
.C(n_439),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_469),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_436),
.B(n_304),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_468),
.B(n_483),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_435),
.B(n_400),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_470),
.B(n_471),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_414),
.Y(n_471)
);

BUFx12_ASAP7_75t_L g472 ( 
.A(n_428),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_472),
.Y(n_490)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_445),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_426),
.A2(n_377),
.B(n_375),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_414),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_477),
.Y(n_491)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_409),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_478),
.A2(n_481),
.B1(n_440),
.B2(n_413),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_439),
.B(n_365),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_409),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_480),
.B(n_482),
.Y(n_512)
);

BUFx4f_ASAP7_75t_L g481 ( 
.A(n_428),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_431),
.B(n_373),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_435),
.B(n_362),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_448),
.B(n_438),
.Y(n_489)
);

CKINVDCx14_ASAP7_75t_R g523 ( 
.A(n_489),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_466),
.A2(n_415),
.B1(n_426),
.B2(n_433),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_492),
.A2(n_495),
.B1(n_503),
.B2(n_516),
.Y(n_527)
);

AO22x1_ASAP7_75t_L g494 ( 
.A1(n_449),
.A2(n_418),
.B1(n_430),
.B2(n_425),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_494),
.B(n_467),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_466),
.A2(n_475),
.B1(n_462),
.B2(n_480),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_496),
.B(n_497),
.C(n_498),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_464),
.B(n_415),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_365),
.C(n_442),
.Y(n_498)
);

OAI32xp33_ASAP7_75t_L g499 ( 
.A1(n_462),
.A2(n_429),
.A3(n_419),
.B1(n_413),
.B2(n_441),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_499),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_465),
.B(n_444),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_500),
.B(n_459),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_502),
.B(n_506),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_477),
.A2(n_429),
.B1(n_440),
.B2(n_441),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_451),
.B(n_434),
.C(n_387),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_505),
.B(n_507),
.C(n_518),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_478),
.B(n_416),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_465),
.A2(n_471),
.B1(n_476),
.B2(n_450),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_509),
.A2(n_511),
.B1(n_482),
.B2(n_467),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_454),
.A2(n_413),
.B1(n_440),
.B2(n_447),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_456),
.B(n_423),
.Y(n_514)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_514),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_454),
.A2(n_421),
.B1(n_413),
.B2(n_437),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_457),
.B(n_424),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_519),
.Y(n_563)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_520),
.Y(n_565)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_484),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_521),
.B(n_524),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_423),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_522),
.B(n_537),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_484),
.Y(n_524)
);

AOI22x1_ASAP7_75t_L g551 ( 
.A1(n_525),
.A2(n_526),
.B1(n_516),
.B2(n_487),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_515),
.A2(n_474),
.B1(n_452),
.B2(n_421),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_528),
.A2(n_542),
.B1(n_545),
.B2(n_546),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_490),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_532),
.B(n_535),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_509),
.A2(n_467),
.B1(n_452),
.B2(n_457),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_533),
.A2(n_540),
.B1(n_547),
.B2(n_502),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_496),
.B(n_473),
.C(n_461),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_534),
.B(n_513),
.Y(n_553)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_485),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_517),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_536),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_515),
.B(n_395),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_511),
.A2(n_467),
.B1(n_470),
.B2(n_469),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_490),
.Y(n_541)
);

INVxp33_ASAP7_75t_L g564 ( 
.A(n_541),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_503),
.A2(n_453),
.B1(n_443),
.B2(n_481),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_512),
.B(n_443),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_543),
.Y(n_555)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_485),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_544),
.Y(n_561)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_501),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_504),
.A2(n_481),
.B1(n_427),
.B2(n_428),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_504),
.A2(n_487),
.B1(n_493),
.B2(n_508),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_493),
.A2(n_411),
.B(n_422),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g560 ( 
.A1(n_548),
.A2(n_518),
.B(n_499),
.Y(n_560)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_501),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_549),
.A2(n_508),
.B1(n_513),
.B2(n_510),
.Y(n_550)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_550),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_551),
.A2(n_556),
.B1(n_572),
.B2(n_542),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_534),
.B(n_505),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_552),
.B(n_558),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_553),
.B(n_554),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_SL g554 ( 
.A(n_530),
.B(n_492),
.C(n_510),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_539),
.B(n_486),
.Y(n_557)
);

CKINVDCx14_ASAP7_75t_R g579 ( 
.A(n_557),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_529),
.B(n_530),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_560),
.A2(n_574),
.B(n_569),
.Y(n_593)
);

FAx1_ASAP7_75t_SL g566 ( 
.A(n_547),
.B(n_498),
.CI(n_495),
.CON(n_566),
.SN(n_566)
);

FAx1_ASAP7_75t_SL g589 ( 
.A(n_566),
.B(n_535),
.CI(n_394),
.CON(n_589),
.SN(n_589)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_529),
.B(n_497),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_568),
.B(n_569),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_540),
.B(n_507),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_533),
.B(n_494),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_570),
.B(n_574),
.C(n_549),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_538),
.A2(n_494),
.B1(n_491),
.B2(n_391),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_527),
.B(n_341),
.Y(n_574)
);

BUFx12_ASAP7_75t_L g575 ( 
.A(n_564),
.Y(n_575)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_575),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_576),
.A2(n_552),
.B1(n_446),
.B2(n_472),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_556),
.A2(n_538),
.B1(n_527),
.B2(n_531),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_578),
.A2(n_584),
.B1(n_401),
.B2(n_405),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_573),
.B(n_536),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_581),
.B(n_583),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_571),
.A2(n_555),
.B1(n_531),
.B2(n_562),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_582),
.A2(n_586),
.B1(n_566),
.B2(n_565),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_567),
.B(n_519),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_572),
.A2(n_531),
.B1(n_525),
.B2(n_523),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_570),
.A2(n_521),
.B1(n_543),
.B2(n_548),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_587),
.B(n_590),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_560),
.A2(n_545),
.B(n_544),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_588),
.A2(n_591),
.B(n_584),
.Y(n_612)
);

XOR2x2_ASAP7_75t_L g598 ( 
.A(n_589),
.B(n_593),
.Y(n_598)
);

INVx13_ASAP7_75t_L g590 ( 
.A(n_564),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_551),
.A2(n_532),
.B(n_541),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_559),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_592),
.B(n_367),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_563),
.B(n_561),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_594),
.A2(n_472),
.B(n_369),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_596),
.B(n_599),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_580),
.B(n_558),
.C(n_568),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_597),
.B(n_601),
.Y(n_625)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_600),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_579),
.B(n_446),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_591),
.A2(n_371),
.B1(n_392),
.B2(n_472),
.Y(n_602)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_602),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_605),
.B(n_611),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_606),
.B(n_608),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_581),
.B(n_327),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_607),
.A2(n_609),
.B(n_594),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_585),
.B(n_593),
.Y(n_608)
);

NOR2xp67_ASAP7_75t_SL g609 ( 
.A(n_577),
.B(n_312),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_580),
.B(n_310),
.Y(n_611)
);

AOI21x1_ASAP7_75t_L g618 ( 
.A1(n_612),
.A2(n_588),
.B(n_595),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_615),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_618),
.A2(n_604),
.B(n_589),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_603),
.B(n_577),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_619),
.B(n_624),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_603),
.B(n_585),
.C(n_587),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_620),
.B(n_621),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_597),
.B(n_578),
.C(n_595),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_SL g622 ( 
.A(n_596),
.B(n_582),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_622),
.B(n_598),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_604),
.B(n_583),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_608),
.B(n_576),
.C(n_586),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_626),
.B(n_610),
.C(n_612),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_627),
.B(n_629),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_623),
.A2(n_602),
.B1(n_598),
.B2(n_589),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_621),
.B(n_611),
.C(n_599),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_630),
.B(n_632),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_631),
.A2(n_617),
.B(n_614),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_614),
.A2(n_592),
.B1(n_590),
.B2(n_575),
.Y(n_632)
);

CKINVDCx14_ASAP7_75t_R g634 ( 
.A(n_625),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_634),
.B(n_636),
.Y(n_644)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_635),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_616),
.A2(n_590),
.B1(n_575),
.B2(n_305),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g638 ( 
.A(n_633),
.B(n_620),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_638),
.B(n_641),
.Y(n_650)
);

AOI221xp5_ASAP7_75t_L g639 ( 
.A1(n_637),
.A2(n_613),
.B1(n_626),
.B2(n_622),
.C(n_617),
.Y(n_639)
);

O2A1O1Ixp33_ASAP7_75t_SL g646 ( 
.A1(n_639),
.A2(n_631),
.B(n_628),
.C(n_629),
.Y(n_646)
);

CKINVDCx16_ASAP7_75t_R g641 ( 
.A(n_627),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_642),
.A2(n_630),
.B(n_575),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_646),
.A2(n_647),
.B(n_648),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_SL g648 ( 
.A1(n_645),
.A2(n_312),
.B(n_328),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_643),
.A2(n_318),
.B(n_306),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_649),
.B(n_348),
.Y(n_653)
);

AOI322xp5_ASAP7_75t_L g651 ( 
.A1(n_650),
.A2(n_644),
.A3(n_640),
.B1(n_641),
.B2(n_305),
.C1(n_343),
.C2(n_306),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_651),
.A2(n_653),
.B(n_325),
.Y(n_654)
);

NOR3xp33_ASAP7_75t_SL g655 ( 
.A(n_654),
.B(n_652),
.C(n_322),
.Y(n_655)
);

BUFx24_ASAP7_75t_SL g656 ( 
.A(n_655),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_656),
.B(n_325),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_657),
.A2(n_322),
.B(n_522),
.Y(n_658)
);


endmodule