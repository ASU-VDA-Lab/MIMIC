module fake_jpeg_26991_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_44),
.Y(n_60)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_36),
.Y(n_62)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_57),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_36),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_45),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_30),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_30),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_17),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_81),
.Y(n_103)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_39),
.B1(n_37),
.B2(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_96),
.B1(n_52),
.B2(n_42),
.Y(n_108)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_39),
.B1(n_47),
.B2(n_38),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_76),
.A2(n_38),
.B1(n_47),
.B2(n_37),
.Y(n_127)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_79),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_22),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_82),
.Y(n_129)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_87),
.Y(n_105)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx6f_ASAP7_75t_SL g123 ( 
.A(n_85),
.Y(n_123)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_91),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_98),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_19),
.B1(n_39),
.B2(n_34),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_22),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_33),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_19),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_58),
.B(n_44),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_75),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_128),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_112),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_21),
.B(n_23),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_119),
.B(n_121),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_127),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_45),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_73),
.A2(n_58),
.B(n_76),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_73),
.A2(n_19),
.B1(n_34),
.B2(n_21),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_101),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_23),
.Y(n_128)
);

MAJx3_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_73),
.C(n_42),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_137),
.B(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_122),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_0),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_120),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_140),
.Y(n_180)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_145),
.B1(n_155),
.B2(n_158),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_149),
.Y(n_167)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_33),
.Y(n_146)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_126),
.B1(n_93),
.B2(n_85),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_156),
.B1(n_129),
.B2(n_64),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_28),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_28),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_157),
.Y(n_168)
);

CKINVDCx12_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_113),
.A2(n_79),
.B1(n_78),
.B2(n_65),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_30),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_108),
.B1(n_119),
.B2(n_115),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_178),
.B1(n_183),
.B2(n_156),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_121),
.C(n_103),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_179),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_134),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_174),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_103),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_77),
.B1(n_109),
.B2(n_102),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_128),
.B(n_111),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_130),
.A2(n_64),
.B1(n_102),
.B2(n_109),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_182),
.B1(n_74),
.B2(n_49),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_133),
.A2(n_129),
.B1(n_43),
.B2(n_37),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_49),
.C(n_104),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_189),
.Y(n_218)
);

NAND2x1_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_148),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_186),
.A2(n_190),
.B(n_118),
.Y(n_221)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_191),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_49),
.C(n_104),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_145),
.A2(n_43),
.B1(n_47),
.B2(n_38),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_122),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_194),
.B(n_195),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_199),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_197),
.Y(n_247)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_200),
.A2(n_204),
.B(n_211),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_171),
.B(n_135),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_174),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_219),
.Y(n_233)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_205),
.Y(n_237)
);

AND2x2_ASAP7_75t_SL g204 ( 
.A(n_177),
.B(n_67),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_215),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_141),
.B1(n_25),
.B2(n_31),
.Y(n_207)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_25),
.B1(n_36),
.B2(n_35),
.Y(n_208)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

AO21x2_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_142),
.B(n_74),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_216),
.B1(n_176),
.B2(n_67),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_172),
.B(n_24),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_210),
.B(n_212),
.Y(n_230)
);

NAND2xp33_ASAP7_75t_SL g211 ( 
.A(n_169),
.B(n_69),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_118),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_213),
.A2(n_221),
.B(n_187),
.Y(n_246)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_160),
.A2(n_94),
.B1(n_92),
.B2(n_95),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_160),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_184),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_35),
.B1(n_31),
.B2(n_24),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_82),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_24),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_162),
.C(n_163),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_214),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_225),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_229),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_218),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_217),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_238),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_170),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_246),
.B(n_197),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_161),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_176),
.Y(n_252)
);

AOI22x1_ASAP7_75t_SL g245 ( 
.A1(n_209),
.A2(n_161),
.B1(n_180),
.B2(n_159),
.Y(n_245)
);

OAI22x1_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_248),
.B1(n_204),
.B2(n_216),
.Y(n_257)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_198),
.B(n_1),
.C(n_2),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_249),
.B(n_1),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_250),
.Y(n_286)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_239),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_266),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_193),
.C(n_211),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_256),
.B(n_270),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_257),
.A2(n_260),
.B1(n_264),
.B2(n_235),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_237),
.A2(n_219),
.B1(n_218),
.B2(n_202),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_263),
.C(n_268),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_193),
.C(n_223),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_69),
.B1(n_67),
.B2(n_50),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_224),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_234),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_269),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_26),
.C(n_20),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_231),
.B1(n_226),
.B2(n_240),
.Y(n_271)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_271),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_260),
.C(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_278),
.B(n_282),
.Y(n_294)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_287),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_246),
.C(n_228),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_284),
.C(n_285),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_228),
.C(n_241),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_241),
.C(n_232),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_244),
.C(n_248),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_254),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_259),
.B1(n_269),
.B2(n_236),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_289),
.A2(n_300),
.B1(n_4),
.B2(n_5),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_247),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_291),
.A2(n_299),
.B(n_1),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_301),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_247),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_298),
.Y(n_307)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_248),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_227),
.B(n_248),
.C(n_229),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_283),
.A2(n_35),
.B1(n_31),
.B2(n_3),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_26),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_26),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_279),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_272),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_4),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_297),
.B(n_284),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_309),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_275),
.C(n_286),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_314),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_10),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_290),
.C(n_295),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_292),
.C(n_299),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_294),
.A2(n_2),
.B(n_3),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_289),
.B(n_7),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_316),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_304),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_318),
.B(n_321),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_319),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_306),
.B(n_10),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_324),
.B(n_325),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_312),
.B(n_10),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_308),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_329),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_317),
.A2(n_318),
.B(n_325),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_309),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_332),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_318),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_307),
.C(n_20),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_334),
.A2(n_332),
.B1(n_327),
.B2(n_328),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_333),
.B(n_335),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_11),
.B(n_12),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_11),
.Y(n_339)
);

OAI21x1_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_12),
.B(n_13),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_14),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_14),
.B(n_26),
.Y(n_342)
);


endmodule