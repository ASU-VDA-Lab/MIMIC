module fake_ibex_1564_n_4545 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_840, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_232, n_380, n_749, n_281, n_559, n_425, n_4545);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_840;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4545;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4449;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2607;
wire n_1382;
wire n_3548;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_845;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_4514;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_3605;
wire n_930;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4343;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4353;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4421;
wire n_4179;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_963;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3904;
wire n_3135;
wire n_3440;
wire n_4378;
wire n_850;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_4477;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_4418;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_875;
wire n_1307;
wire n_4431;
wire n_1327;
wire n_2644;
wire n_4445;
wire n_876;
wire n_3211;
wire n_3479;
wire n_1840;
wire n_2837;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_4470;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3896;
wire n_3753;
wire n_2192;
wire n_4423;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_3353;
wire n_2918;
wire n_3976;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_4450;
wire n_3969;
wire n_4467;
wire n_1081;
wire n_4437;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_4447;
wire n_4491;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3949;
wire n_3507;
wire n_3884;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_4389;
wire n_4510;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_4312;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_4430;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_4433;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_4428;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_3809;
wire n_979;
wire n_4503;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4517;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_4511;
wire n_1007;
wire n_2253;
wire n_4479;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_4422;
wire n_1219;
wire n_4513;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_4481;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_1326;
wire n_971;
wire n_4444;
wire n_1350;
wire n_3627;
wire n_906;
wire n_4499;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_4533;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4455;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4518;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_4480;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_4535;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_4290;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_4252;
wire n_1332;
wire n_2660;
wire n_3971;
wire n_4505;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4522;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_4476;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4126;
wire n_3583;
wire n_2019;
wire n_4103;
wire n_1407;
wire n_3282;
wire n_4435;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_4411;
wire n_4523;
wire n_4408;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_4489;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_4419;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_2599;
wire n_974;
wire n_1036;
wire n_3626;
wire n_1831;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_4494;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_4542;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_4374;
wire n_1140;
wire n_1985;
wire n_4375;
wire n_4501;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_4403;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_4230;
wire n_859;
wire n_3849;
wire n_965;
wire n_1109;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4469;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_4460;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4504;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_4527;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_4485;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_3364;
wire n_1236;
wire n_4384;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_4537;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4407;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_4462;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_4540;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_4490;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_3503;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_4362;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2910;
wire n_2552;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_4414;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_4525;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_4443;
wire n_1682;
wire n_4151;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_847;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_4424;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_4415;
wire n_1345;
wire n_4215;
wire n_4456;
wire n_4315;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_3578;
wire n_954;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_4492;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_4500;
wire n_998;
wire n_1395;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_4427;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_3829;
wire n_1864;
wire n_943;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_2398;
wire n_1836;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_3646;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_863;
wire n_2185;
wire n_4141;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_4496;
wire n_2507;
wire n_2759;
wire n_3682;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3434;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1185;
wire n_1683;
wire n_4256;
wire n_3575;
wire n_4454;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_4278;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_4458;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_3158;
wire n_2045;
wire n_2427;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_4276;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1941;
wire n_1707;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_4185;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_920;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_4441;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_2997;
wire n_3314;
wire n_961;
wire n_991;
wire n_1331;
wire n_1223;
wire n_1349;
wire n_2127;
wire n_3891;
wire n_3747;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_4536;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_4497;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_4512;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_4483;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4488;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1601;
wire n_1294;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4142;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1458;
wire n_1694;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3696;
wire n_3113;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_4286;
wire n_4429;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1962;
wire n_1225;
wire n_2346;
wire n_982;
wire n_4438;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3912;
wire n_3778;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_2959;
wire n_1625;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_4498;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1348;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_3356;
wire n_1191;
wire n_2004;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_3899;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_4149;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_4319;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_3773;
wire n_2528;
wire n_4383;
wire n_3216;
wire n_2548;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_4543;
wire n_4466;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1946;
wire n_1726;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_3506;
wire n_2845;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_3162;
wire n_2732;
wire n_2984;
wire n_4436;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_4538;
wire n_3333;
wire n_3096;
wire n_4509;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_4434;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_4367;
wire n_950;
wire n_3139;
wire n_2700;
wire n_1222;
wire n_4282;
wire n_1630;
wire n_3408;
wire n_4475;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_4410;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_4440;
wire n_1885;
wire n_1989;
wire n_1740;
wire n_3604;
wire n_1838;
wire n_3540;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_4529;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2576;
wire n_2348;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_4200;
wire n_4162;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_4439;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_4487;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4519;
wire n_4148;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_4541;
wire n_4515;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_4530;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_2816;
wire n_2433;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_2658;
wire n_3576;
wire n_3236;
wire n_3109;
wire n_1961;
wire n_3491;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_4265;
wire n_3062;
wire n_4524;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2864;
wire n_2406;
wire n_1632;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4017;
wire n_1542;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1547;
wire n_3497;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_956;
wire n_3561;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_2574;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_2911;
wire n_1623;
wire n_861;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_4453;
wire n_1098;
wire n_4474;
wire n_1518;
wire n_1366;
wire n_4350;
wire n_4380;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_3102;
wire n_2872;
wire n_3173;
wire n_4345;
wire n_4281;
wire n_4478;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_4473;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_4464;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_854;
wire n_4432;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_3543;
wire n_1734;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4461;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_4516;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_4528;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_4502;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_914;
wire n_4147;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_4471;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_4386;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_3296;
wire n_1911;
wire n_2293;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_4482;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_4493;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_1488;
wire n_849;
wire n_980;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3557;
wire n_1074;
wire n_3225;
wire n_3380;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_1022;
wire n_4412;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3286;
wire n_999;
wire n_2634;
wire n_3124;
wire n_2982;
wire n_1092;
wire n_4038;
wire n_4472;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_4521;
wire n_1230;
wire n_4459;
wire n_1027;
wire n_1516;
wire n_3893;
wire n_4484;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2303;
wire n_949;
wire n_2104;
wire n_2653;
wire n_2357;
wire n_2618;
wire n_2855;
wire n_3938;
wire n_4354;
wire n_924;
wire n_4448;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4401;
wire n_4532;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_3056;
wire n_2453;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_3052;
wire n_2443;
wire n_3189;
wire n_4544;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_2066;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_4275;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_4468;
wire n_1736;
wire n_4442;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2749;
wire n_888;
wire n_2378;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_4539;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_3275;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_2670;
wire n_4486;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2726;
wire n_2917;
wire n_2619;
wire n_3873;
wire n_3738;
wire n_4506;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_4327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_4465;
wire n_1355;
wire n_3691;
wire n_4452;
wire n_2544;
wire n_856;
wire n_3193;
wire n_4534;
wire n_3635;
wire n_3501;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_4183;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_4508;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_4425;
wire n_3980;
wire n_2673;
wire n_2430;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_3180;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_795),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_96),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_164),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_678),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_655),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_216),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_750),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_495),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_542),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_141),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_164),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_266),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_183),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_836),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_530),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_123),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_761),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_762),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_364),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_691),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_84),
.Y(n_862)
);

BUFx8_ASAP7_75t_SL g863 ( 
.A(n_482),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_784),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_287),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_805),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_626),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_522),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_723),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_540),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_782),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_125),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_48),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_793),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_570),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_47),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_63),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_692),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_554),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_343),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_354),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_395),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_302),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_673),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_552),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_92),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_89),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_599),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_665),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_433),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_71),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_361),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_315),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_317),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_786),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_242),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_210),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_293),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_267),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_266),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_216),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_124),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_776),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_79),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_405),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_709),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_212),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_222),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_690),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_394),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_837),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_328),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_504),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_691),
.Y(n_914)
);

BUFx10_ASAP7_75t_L g915 ( 
.A(n_430),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_417),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_788),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_739),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_753),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_692),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_171),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_401),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_464),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_434),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_357),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_138),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_126),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_794),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_562),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_722),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_427),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_320),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_569),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_242),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_787),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_751),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_234),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_443),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_588),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_358),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_489),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_81),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_720),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_451),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_498),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_610),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_774),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_624),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_260),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_363),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_182),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_828),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_751),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_832),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_807),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_481),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_407),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_641),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_227),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_655),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_572),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_137),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_49),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_672),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_391),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_745),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_340),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_754),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_396),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_58),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_15),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_150),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_209),
.Y(n_973)
);

BUFx2_ASAP7_75t_R g974 ( 
.A(n_570),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_149),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_799),
.Y(n_976)
);

BUFx10_ASAP7_75t_L g977 ( 
.A(n_457),
.Y(n_977)
);

CKINVDCx16_ASAP7_75t_R g978 ( 
.A(n_73),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_287),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_277),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_177),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_64),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_227),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_391),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_532),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_770),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_262),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_749),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_85),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_210),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_17),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_673),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_693),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_693),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_550),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_779),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_746),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_624),
.Y(n_998)
);

BUFx10_ASAP7_75t_L g999 ( 
.A(n_39),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_82),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_594),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_370),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_783),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_595),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_498),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_122),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_409),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_798),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_533),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_234),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_333),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_594),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_528),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_703),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_797),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_807),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_470),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_244),
.Y(n_1018)
);

BUFx10_ASAP7_75t_L g1019 ( 
.A(n_404),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_395),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_204),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_176),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_764),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_712),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_697),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_778),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_764),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_3),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_269),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_438),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_626),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_756),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_201),
.Y(n_1033)
);

CKINVDCx16_ASAP7_75t_R g1034 ( 
.A(n_504),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_318),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_707),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_219),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_351),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_48),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_250),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_630),
.Y(n_1041)
);

CKINVDCx16_ASAP7_75t_R g1042 ( 
.A(n_194),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_789),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_172),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_33),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_615),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_729),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_747),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_838),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_17),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_501),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_687),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_43),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_432),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_763),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_439),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_380),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_15),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_748),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_268),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_796),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_100),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_326),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_638),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_638),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_679),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_258),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_620),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_147),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_271),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_722),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_606),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_646),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_428),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_736),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_777),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_307),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_471),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_200),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_798),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_96),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_381),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_635),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_468),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_772),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_458),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_88),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_679),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_384),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_85),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_84),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_610),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_125),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_604),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_273),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_450),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_603),
.Y(n_1097)
);

BUFx10_ASAP7_75t_L g1098 ( 
.A(n_388),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_702),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_706),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_398),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_567),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_810),
.Y(n_1103)
);

CKINVDCx14_ASAP7_75t_R g1104 ( 
.A(n_552),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_200),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_718),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_485),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_20),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_471),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_573),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_777),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_110),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_781),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_127),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_559),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_441),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_768),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_767),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_549),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_265),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_482),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_418),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_246),
.Y(n_1123)
);

BUFx10_ASAP7_75t_L g1124 ( 
.A(n_377),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_677),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_201),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_670),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_198),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_180),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_520),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_230),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_90),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_295),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_836),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_791),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_773),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_123),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_66),
.Y(n_1138)
);

BUFx2_ASAP7_75t_SL g1139 ( 
.A(n_483),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_689),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_105),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_328),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_158),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_473),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_790),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_631),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_675),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_780),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_113),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_209),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_10),
.Y(n_1151)
);

CKINVDCx14_ASAP7_75t_R g1152 ( 
.A(n_62),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_627),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_792),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_90),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_58),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_94),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_775),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_335),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_569),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_780),
.Y(n_1161)
);

CKINVDCx16_ASAP7_75t_R g1162 ( 
.A(n_664),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_547),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_513),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_453),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_384),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_145),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_701),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_253),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_406),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_132),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_405),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_735),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_618),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_657),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_232),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_60),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_215),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_136),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_346),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_392),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_94),
.Y(n_1182)
);

BUFx10_ASAP7_75t_L g1183 ( 
.A(n_483),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_787),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_666),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_416),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_540),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_71),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_704),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_745),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_343),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_680),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_658),
.Y(n_1193)
);

CKINVDCx16_ASAP7_75t_R g1194 ( 
.A(n_40),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_612),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_713),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_238),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_416),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_766),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_718),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_298),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_306),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_55),
.Y(n_1203)
);

BUFx5_ASAP7_75t_L g1204 ( 
.A(n_750),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_130),
.Y(n_1205)
);

INVxp33_ASAP7_75t_SL g1206 ( 
.A(n_833),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_643),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_477),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_803),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_689),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_485),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_276),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_765),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_233),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_467),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_805),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_758),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_20),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_327),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_43),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_579),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_785),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_35),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_759),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_717),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_301),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_526),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_269),
.Y(n_1228)
);

CKINVDCx16_ASAP7_75t_R g1229 ( 
.A(n_35),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_67),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_363),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_390),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_324),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_497),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_360),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_385),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_833),
.Y(n_1237)
);

BUFx10_ASAP7_75t_L g1238 ( 
.A(n_160),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_279),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_588),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_104),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_399),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_98),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_738),
.Y(n_1244)
);

BUFx8_ASAP7_75t_SL g1245 ( 
.A(n_648),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_428),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_812),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_480),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_822),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_98),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_374),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_606),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_712),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_401),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_759),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_105),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_808),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_771),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_118),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_427),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_809),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_284),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_766),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_839),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_258),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_506),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_527),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_436),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_61),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_755),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_184),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_340),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_121),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_505),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_366),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_177),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_93),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_248),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_549),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_313),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_282),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_207),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_826),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_146),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_59),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_189),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_148),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_472),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_651),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_653),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_708),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_145),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_103),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_479),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_120),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_352),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_183),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_179),
.Y(n_1298)
);

BUFx10_ASAP7_75t_L g1299 ( 
.A(n_114),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_757),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_649),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_198),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_546),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_318),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_509),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_645),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_320),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_814),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_319),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_675),
.Y(n_1310)
);

BUFx5_ASAP7_75t_L g1311 ( 
.A(n_63),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_92),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_180),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_772),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_24),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_559),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_816),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_659),
.Y(n_1318)
);

BUFx5_ASAP7_75t_L g1319 ( 
.A(n_211),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_421),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_211),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_562),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_434),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_429),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_80),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_40),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_508),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_752),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_213),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_760),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_544),
.Y(n_1331)
);

BUFx10_ASAP7_75t_L g1332 ( 
.A(n_567),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_367),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_356),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_762),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_389),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_346),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_744),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_31),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_414),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_589),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_537),
.Y(n_1342)
);

BUFx5_ASAP7_75t_L g1343 ( 
.A(n_621),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_295),
.Y(n_1344)
);

INVxp67_ASAP7_75t_SL g1345 ( 
.A(n_769),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_800),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_645),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_816),
.Y(n_1348)
);

BUFx5_ASAP7_75t_L g1349 ( 
.A(n_616),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_338),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_619),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1204),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_880),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_941),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_908),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_867),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_863),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_908),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_867),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_956),
.B(n_0),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1204),
.Y(n_1361)
);

INVx5_ASAP7_75t_L g1362 ( 
.A(n_1061),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_976),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1204),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_966),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1061),
.B(n_0),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_908),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1017),
.B(n_0),
.Y(n_1368)
);

BUFx12f_ASAP7_75t_L g1369 ( 
.A(n_915),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_908),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_981),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1131),
.B(n_1),
.Y(n_1372)
);

XNOR2xp5_ASAP7_75t_L g1373 ( 
.A(n_1028),
.B(n_1),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1154),
.B(n_1179),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_981),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1103),
.B(n_1),
.Y(n_1376)
);

INVx5_ASAP7_75t_L g1377 ( 
.A(n_1061),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1204),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_863),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_886),
.B(n_2),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_915),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1204),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_915),
.Y(n_1383)
);

INVx5_ASAP7_75t_L g1384 ( 
.A(n_981),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_977),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1223),
.B(n_886),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1204),
.Y(n_1387)
);

INVx5_ASAP7_75t_L g1388 ( 
.A(n_981),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1205),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_895),
.B(n_2),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_895),
.B(n_2),
.Y(n_1391)
);

INVxp67_ASAP7_75t_L g1392 ( 
.A(n_942),
.Y(n_1392)
);

AND2x6_ASAP7_75t_L g1393 ( 
.A(n_966),
.B(n_3),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_978),
.B(n_3),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1205),
.Y(n_1395)
);

INVx5_ASAP7_75t_L g1396 ( 
.A(n_1205),
.Y(n_1396)
);

BUFx12f_ASAP7_75t_L g1397 ( 
.A(n_977),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_986),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1204),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_942),
.B(n_4),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_996),
.B(n_4),
.Y(n_1401)
);

INVx5_ASAP7_75t_L g1402 ( 
.A(n_1205),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1243),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1243),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_996),
.B(n_6),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1243),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1034),
.B(n_5),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1243),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1000),
.B(n_6),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_977),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1104),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_999),
.Y(n_1412)
);

INVx5_ASAP7_75t_L g1413 ( 
.A(n_1244),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_999),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1244),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1000),
.B(n_7),
.Y(n_1416)
);

INVx5_ASAP7_75t_L g1417 ( 
.A(n_1244),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1042),
.B(n_5),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1244),
.Y(n_1419)
);

CKINVDCx14_ASAP7_75t_R g1420 ( 
.A(n_1152),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1311),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1162),
.B(n_7),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1006),
.B(n_9),
.Y(n_1423)
);

INVx5_ASAP7_75t_L g1424 ( 
.A(n_1264),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1194),
.B(n_8),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1006),
.B(n_8),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1206),
.B(n_9),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1206),
.B(n_10),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1311),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1302),
.B(n_11),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1302),
.B(n_12),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_878),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_878),
.Y(n_1433)
);

INVx5_ASAP7_75t_L g1434 ( 
.A(n_1264),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_999),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1351),
.B(n_11),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_1028),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_986),
.B(n_12),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_993),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1264),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_993),
.B(n_1059),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1264),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_843),
.B(n_13),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1059),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1313),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1062),
.Y(n_1446)
);

INVx5_ASAP7_75t_L g1447 ( 
.A(n_1313),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1062),
.B(n_13),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1229),
.B(n_16),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1311),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1019),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1072),
.Y(n_1452)
);

BUFx12f_ASAP7_75t_L g1453 ( 
.A(n_1019),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1311),
.Y(n_1454)
);

INVx5_ASAP7_75t_L g1455 ( 
.A(n_1313),
.Y(n_1455)
);

INVx5_ASAP7_75t_L g1456 ( 
.A(n_1313),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1072),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_859),
.B(n_16),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1311),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1311),
.B(n_14),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_948),
.B(n_14),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1145),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1151),
.B(n_19),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1311),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_SL g1465 ( 
.A(n_1319),
.B(n_18),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1145),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1236),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1236),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1019),
.B(n_18),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1319),
.Y(n_1470)
);

BUFx8_ASAP7_75t_L g1471 ( 
.A(n_1319),
.Y(n_1471)
);

INVx5_ASAP7_75t_L g1472 ( 
.A(n_1098),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1258),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1319),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1258),
.B(n_1261),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_845),
.B(n_19),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1319),
.B(n_21),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1098),
.B(n_21),
.Y(n_1478)
);

NAND2x1p5_ASAP7_75t_L g1479 ( 
.A(n_1261),
.B(n_22),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1353),
.A2(n_882),
.B1(n_883),
.B2(n_881),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1374),
.B(n_1098),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1432),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1354),
.B(n_1363),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1449),
.A2(n_881),
.B1(n_883),
.B2(n_882),
.Y(n_1484)
);

AO22x2_ASAP7_75t_L g1485 ( 
.A1(n_1394),
.A2(n_974),
.B1(n_1139),
.B2(n_1345),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1433),
.A2(n_887),
.B1(n_889),
.B2(n_884),
.Y(n_1486)
);

AO22x2_ASAP7_75t_L g1487 ( 
.A1(n_1407),
.A2(n_874),
.B1(n_888),
.B2(n_869),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1366),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1357),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1360),
.A2(n_887),
.B1(n_889),
.B2(n_884),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1376),
.A2(n_892),
.B1(n_894),
.B2(n_891),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1462),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1366),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1379),
.A2(n_892),
.B1(n_894),
.B2(n_891),
.Y(n_1494)
);

AO22x2_ASAP7_75t_L g1495 ( 
.A1(n_1418),
.A2(n_997),
.B1(n_1030),
.B2(n_905),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_SL g1496 ( 
.A(n_1380),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1411),
.B(n_1124),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1369),
.B(n_1245),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1400),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1420),
.B(n_1124),
.Y(n_1500)
);

AO22x2_ASAP7_75t_L g1501 ( 
.A1(n_1422),
.A2(n_1425),
.B1(n_1400),
.B2(n_1401),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1479),
.A2(n_898),
.B1(n_1340),
.B2(n_896),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1386),
.B(n_1348),
.Y(n_1503)
);

OAI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1436),
.A2(n_898),
.B1(n_1340),
.B2(n_896),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1472),
.B(n_1124),
.Y(n_1505)
);

AO22x2_ASAP7_75t_L g1506 ( 
.A1(n_1401),
.A2(n_1080),
.B1(n_1114),
.B2(n_1058),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1426),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1368),
.A2(n_1344),
.B1(n_1347),
.B2(n_1342),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1462),
.Y(n_1509)
);

NOR2x1p5_ASAP7_75t_L g1510 ( 
.A(n_1397),
.B(n_1342),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1372),
.A2(n_1347),
.B1(n_1348),
.B2(n_1344),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1392),
.B(n_842),
.Y(n_1512)
);

OAI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1465),
.A2(n_1350),
.B1(n_1463),
.B2(n_1458),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1380),
.A2(n_1350),
.B1(n_847),
.B2(n_849),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1426),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1462),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1393),
.A2(n_850),
.B1(n_852),
.B2(n_844),
.Y(n_1517)
);

BUFx10_ASAP7_75t_L g1518 ( 
.A(n_1430),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1452),
.B(n_855),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1472),
.B(n_1183),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1430),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1437),
.A2(n_890),
.B1(n_909),
.B2(n_853),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1393),
.A2(n_858),
.B1(n_861),
.B2(n_860),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1393),
.A2(n_865),
.B1(n_870),
.B2(n_868),
.Y(n_1524)
);

AND2x2_ASAP7_75t_SL g1525 ( 
.A(n_1478),
.B(n_851),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1472),
.B(n_1183),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1436),
.A2(n_1341),
.B1(n_1335),
.B2(n_890),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1393),
.A2(n_871),
.B1(n_875),
.B2(n_873),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1465),
.A2(n_877),
.B1(n_899),
.B2(n_876),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1373),
.A2(n_909),
.B1(n_962),
.B2(n_853),
.Y(n_1530)
);

NAND3x1_ASAP7_75t_L g1531 ( 
.A(n_1427),
.B(n_1245),
.C(n_982),
.Y(n_1531)
);

OAI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1443),
.A2(n_982),
.B1(n_989),
.B2(n_962),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1466),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1457),
.B(n_1183),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1438),
.Y(n_1535)
);

AO22x2_ASAP7_75t_L g1536 ( 
.A1(n_1438),
.A2(n_1167),
.B1(n_1170),
.B2(n_1122),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1467),
.B(n_1238),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1466),
.Y(n_1538)
);

NAND3x1_ASAP7_75t_L g1539 ( 
.A(n_1428),
.B(n_991),
.C(n_989),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1448),
.A2(n_901),
.B1(n_903),
.B2(n_900),
.Y(n_1540)
);

OAI22xp33_ASAP7_75t_SL g1541 ( 
.A1(n_1390),
.A2(n_906),
.B1(n_912),
.B2(n_904),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1383),
.B(n_1238),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1448),
.A2(n_917),
.B1(n_918),
.B2(n_914),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1410),
.A2(n_921),
.B1(n_922),
.B2(n_920),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1414),
.A2(n_931),
.B1(n_932),
.B2(n_930),
.Y(n_1545)
);

OR2x6_ASAP7_75t_L g1546 ( 
.A(n_1435),
.B(n_933),
.Y(n_1546)
);

OAI22xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1391),
.A2(n_936),
.B1(n_938),
.B2(n_934),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1383),
.B(n_1238),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1385),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_SL g1550 ( 
.A1(n_1453),
.A2(n_1071),
.B1(n_1091),
.B2(n_991),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1381),
.A2(n_944),
.B1(n_945),
.B2(n_943),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1466),
.Y(n_1552)
);

OAI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1443),
.A2(n_1091),
.B1(n_1093),
.B2(n_1071),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1441),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1356),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1441),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1359),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1475),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1385),
.B(n_1412),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1451),
.A2(n_949),
.B1(n_950),
.B2(n_947),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1365),
.Y(n_1561)
);

OA22x2_ASAP7_75t_L g1562 ( 
.A1(n_1412),
.A2(n_1476),
.B1(n_1475),
.B2(n_1409),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1476),
.A2(n_954),
.B1(n_955),
.B2(n_953),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1362),
.B(n_1299),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1398),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1405),
.A2(n_1341),
.B1(n_1335),
.B2(n_1097),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1439),
.Y(n_1567)
);

AO22x2_ASAP7_75t_L g1568 ( 
.A1(n_1416),
.A2(n_1177),
.B1(n_1187),
.B2(n_1172),
.Y(n_1568)
);

OAI22xp33_ASAP7_75t_SL g1569 ( 
.A1(n_1423),
.A2(n_958),
.B1(n_960),
.B2(n_957),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_R g1570 ( 
.A1(n_1469),
.A2(n_1227),
.B1(n_848),
.B2(n_854),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1444),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1362),
.B(n_1299),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1471),
.B(n_1343),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1431),
.B(n_1031),
.Y(n_1574)
);

OA22x2_ASAP7_75t_L g1575 ( 
.A1(n_1460),
.A2(n_963),
.B1(n_1002),
.B2(n_972),
.Y(n_1575)
);

OAI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1477),
.A2(n_964),
.B1(n_969),
.B2(n_961),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1446),
.Y(n_1577)
);

OR2x6_ASAP7_75t_L g1578 ( 
.A(n_1461),
.B(n_1027),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1468),
.Y(n_1579)
);

AO22x2_ASAP7_75t_L g1580 ( 
.A1(n_1473),
.A2(n_1338),
.B1(n_1339),
.B2(n_1333),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1471),
.A2(n_971),
.B1(n_973),
.B2(n_970),
.Y(n_1581)
);

OR2x6_ASAP7_75t_L g1582 ( 
.A(n_1382),
.B(n_851),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1362),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1382),
.B(n_925),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1377),
.B(n_1299),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1377),
.B(n_1324),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1377),
.A2(n_984),
.B1(n_992),
.B2(n_979),
.Y(n_1587)
);

OAI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1387),
.A2(n_1097),
.B1(n_1105),
.B2(n_1093),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1384),
.B(n_1337),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1387),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1421),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1384),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1474),
.A2(n_1001),
.B1(n_1003),
.B2(n_998),
.Y(n_1593)
);

AO22x2_ASAP7_75t_L g1594 ( 
.A1(n_1421),
.A2(n_1346),
.B1(n_1331),
.B2(n_856),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1429),
.B(n_1324),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1384),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1388),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1429),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1450),
.A2(n_1007),
.B1(n_1009),
.B2(n_1005),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1450),
.A2(n_1012),
.B1(n_1014),
.B2(n_1010),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1388),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1474),
.A2(n_1016),
.B1(n_1018),
.B2(n_1015),
.Y(n_1602)
);

BUFx10_ASAP7_75t_L g1603 ( 
.A(n_1355),
.Y(n_1603)
);

AO22x2_ASAP7_75t_L g1604 ( 
.A1(n_1352),
.A2(n_1326),
.B1(n_1325),
.B2(n_857),
.Y(n_1604)
);

OAI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1361),
.A2(n_1142),
.B1(n_1147),
.B2(n_1105),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1364),
.B(n_1324),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1388),
.B(n_1337),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1396),
.Y(n_1608)
);

NOR2x1p5_ASAP7_75t_L g1609 ( 
.A(n_1378),
.B(n_872),
.Y(n_1609)
);

AO22x2_ASAP7_75t_L g1610 ( 
.A1(n_1399),
.A2(n_862),
.B1(n_864),
.B2(n_846),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1454),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1459),
.B(n_866),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1464),
.Y(n_1613)
);

AO22x2_ASAP7_75t_L g1614 ( 
.A1(n_1470),
.A2(n_885),
.B1(n_893),
.B2(n_879),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1396),
.A2(n_1320),
.B1(n_1147),
.B2(n_1155),
.Y(n_1615)
);

OAI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1396),
.A2(n_1320),
.B1(n_1155),
.B2(n_1161),
.Y(n_1616)
);

AO22x2_ASAP7_75t_L g1617 ( 
.A1(n_1402),
.A2(n_902),
.B1(n_907),
.B2(n_897),
.Y(n_1617)
);

AO22x2_ASAP7_75t_L g1618 ( 
.A1(n_1402),
.A2(n_911),
.B1(n_913),
.B2(n_910),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1402),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1413),
.Y(n_1620)
);

NAND3x1_ASAP7_75t_L g1621 ( 
.A(n_1413),
.B(n_1161),
.C(n_1142),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1413),
.A2(n_1021),
.B1(n_1024),
.B2(n_1020),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1456),
.B(n_1332),
.Y(n_1623)
);

AO22x2_ASAP7_75t_L g1624 ( 
.A1(n_1417),
.A2(n_919),
.B1(n_923),
.B2(n_916),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1417),
.A2(n_1029),
.B1(n_1032),
.B2(n_1025),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1417),
.A2(n_1038),
.B1(n_1039),
.B2(n_1033),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1424),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1424),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1424),
.B(n_1332),
.Y(n_1629)
);

OR2x6_ASAP7_75t_L g1630 ( 
.A(n_1355),
.B(n_951),
.Y(n_1630)
);

OAI22xp33_ASAP7_75t_SL g1631 ( 
.A1(n_1434),
.A2(n_1041),
.B1(n_1045),
.B2(n_1040),
.Y(n_1631)
);

NAND3x1_ASAP7_75t_L g1632 ( 
.A(n_1434),
.B(n_1180),
.C(n_1169),
.Y(n_1632)
);

OA22x2_ASAP7_75t_L g1633 ( 
.A1(n_1434),
.A2(n_1069),
.B1(n_1079),
.B2(n_1049),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1447),
.B(n_1332),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1447),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1447),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1455),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1455),
.A2(n_1055),
.B1(n_1060),
.B2(n_1053),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1455),
.Y(n_1639)
);

OAI22xp33_ASAP7_75t_SL g1640 ( 
.A1(n_1456),
.A2(n_1064),
.B1(n_1065),
.B2(n_1063),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1456),
.B(n_1319),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1355),
.B(n_925),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1358),
.Y(n_1643)
);

OR2x6_ASAP7_75t_L g1644 ( 
.A(n_1358),
.B(n_985),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1358),
.B(n_1319),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1367),
.B(n_1343),
.Y(n_1646)
);

AO22x2_ASAP7_75t_L g1647 ( 
.A1(n_1367),
.A2(n_926),
.B1(n_927),
.B2(n_924),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_SL g1648 ( 
.A1(n_1367),
.A2(n_1180),
.B1(n_1182),
.B2(n_1169),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1370),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1370),
.A2(n_1067),
.B1(n_1068),
.B2(n_1066),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1370),
.B(n_1070),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1371),
.Y(n_1652)
);

OAI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1371),
.A2(n_1184),
.B1(n_1235),
.B2(n_1182),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1371),
.Y(n_1654)
);

XOR2xp5_ASAP7_75t_L g1655 ( 
.A(n_1375),
.B(n_1184),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1375),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1375),
.Y(n_1657)
);

NAND3x1_ASAP7_75t_L g1658 ( 
.A(n_1389),
.B(n_1255),
.C(n_1235),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1389),
.A2(n_1074),
.B1(n_1076),
.B2(n_1073),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1389),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1395),
.Y(n_1661)
);

OAI22xp33_ASAP7_75t_SL g1662 ( 
.A1(n_1395),
.A2(n_1082),
.B1(n_1084),
.B2(n_1077),
.Y(n_1662)
);

NAND2xp33_ASAP7_75t_SL g1663 ( 
.A(n_1395),
.B(n_1255),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1403),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1403),
.Y(n_1665)
);

AO22x2_ASAP7_75t_L g1666 ( 
.A1(n_1403),
.A2(n_929),
.B1(n_935),
.B2(n_928),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1404),
.B(n_1085),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1404),
.B(n_1343),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1404),
.B(n_1087),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1406),
.B(n_1343),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1406),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1406),
.Y(n_1672)
);

OAI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1408),
.A2(n_1284),
.B1(n_1310),
.B2(n_1276),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1408),
.A2(n_1284),
.B1(n_1310),
.B2(n_1276),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1408),
.B(n_1343),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1415),
.B(n_1343),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1415),
.B(n_1321),
.Y(n_1677)
);

OAI22xp33_ASAP7_75t_SL g1678 ( 
.A1(n_1415),
.A2(n_1089),
.B1(n_1090),
.B2(n_1088),
.Y(n_1678)
);

OAI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1419),
.A2(n_937),
.B1(n_940),
.B2(n_939),
.Y(n_1679)
);

OAI22xp33_ASAP7_75t_SL g1680 ( 
.A1(n_1419),
.A2(n_1094),
.B1(n_1095),
.B2(n_1092),
.Y(n_1680)
);

AO22x2_ASAP7_75t_L g1681 ( 
.A1(n_1419),
.A2(n_946),
.B1(n_959),
.B2(n_952),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1440),
.A2(n_1099),
.B1(n_1100),
.B2(n_1096),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1440),
.A2(n_1110),
.B1(n_1111),
.B2(n_1101),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1440),
.A2(n_1115),
.B1(n_1117),
.B2(n_1112),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1442),
.Y(n_1685)
);

OAI22xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1442),
.A2(n_1119),
.B1(n_1121),
.B2(n_1118),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1442),
.A2(n_1129),
.B1(n_1133),
.B2(n_1127),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1445),
.A2(n_1136),
.B1(n_1138),
.B2(n_1135),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1445),
.B(n_965),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1445),
.B(n_1343),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1374),
.B(n_1349),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1353),
.A2(n_1141),
.B1(n_1143),
.B2(n_1140),
.Y(n_1692)
);

OAI22xp33_ASAP7_75t_SL g1693 ( 
.A1(n_1479),
.A2(n_1146),
.B1(n_1148),
.B2(n_1144),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1462),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1353),
.A2(n_1150),
.B1(n_1163),
.B2(n_1149),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1353),
.A2(n_1174),
.B1(n_1175),
.B2(n_1173),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1353),
.A2(n_1186),
.B1(n_1188),
.B2(n_1185),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1483),
.B(n_1189),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1554),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1503),
.B(n_1315),
.Y(n_1700)
);

CKINVDCx20_ASAP7_75t_R g1701 ( 
.A(n_1522),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1481),
.B(n_1190),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1556),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1558),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1604),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1604),
.Y(n_1706)
);

XOR2xp5_ASAP7_75t_L g1707 ( 
.A(n_1530),
.B(n_1322),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1610),
.Y(n_1708)
);

NAND2xp33_ASAP7_75t_R g1709 ( 
.A(n_1489),
.B(n_1192),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1610),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1614),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1689),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1614),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1482),
.B(n_1193),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1559),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1488),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1493),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1538),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1499),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_1656),
.Y(n_1720)
);

XNOR2xp5_ASAP7_75t_L g1721 ( 
.A(n_1539),
.B(n_1195),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1647),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1507),
.Y(n_1723)
);

NOR2xp67_ASAP7_75t_L g1724 ( 
.A(n_1517),
.B(n_933),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1647),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1549),
.B(n_1542),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1515),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1521),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1548),
.B(n_1197),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1518),
.Y(n_1730)
);

CKINVDCx14_ASAP7_75t_R g1731 ( 
.A(n_1498),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1594),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1534),
.B(n_1198),
.Y(n_1733)
);

INVxp67_ASAP7_75t_SL g1734 ( 
.A(n_1666),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1594),
.Y(n_1735)
);

CKINVDCx20_ASAP7_75t_R g1736 ( 
.A(n_1550),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1497),
.B(n_1199),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1666),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1681),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1519),
.B(n_1200),
.Y(n_1740)
);

XOR2xp5_ASAP7_75t_L g1741 ( 
.A(n_1485),
.B(n_1336),
.Y(n_1741)
);

BUFx8_ASAP7_75t_L g1742 ( 
.A(n_1496),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_SL g1743 ( 
.A(n_1498),
.Y(n_1743)
);

INVxp33_ASAP7_75t_L g1744 ( 
.A(n_1655),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1681),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1567),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1606),
.B(n_1201),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1595),
.B(n_1349),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1535),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1505),
.B(n_1202),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1546),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1651),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1537),
.B(n_1203),
.Y(n_1753)
);

XOR2xp5_ASAP7_75t_L g1754 ( 
.A(n_1485),
.B(n_1308),
.Y(n_1754)
);

OR2x6_ASAP7_75t_L g1755 ( 
.A(n_1546),
.B(n_951),
.Y(n_1755)
);

XOR2xp5_ASAP7_75t_L g1756 ( 
.A(n_1648),
.B(n_1312),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1677),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1598),
.B(n_1349),
.Y(n_1758)
);

BUFx3_ASAP7_75t_L g1759 ( 
.A(n_1577),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1612),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1580),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1480),
.B(n_1314),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1580),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1691),
.B(n_1582),
.Y(n_1764)
);

INVxp33_ASAP7_75t_SL g1765 ( 
.A(n_1490),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1520),
.B(n_1207),
.Y(n_1766)
);

INVx4_ASAP7_75t_SL g1767 ( 
.A(n_1682),
.Y(n_1767)
);

XOR2xp5_ASAP7_75t_L g1768 ( 
.A(n_1674),
.B(n_1615),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1526),
.B(n_967),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1641),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1525),
.B(n_1208),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1562),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1609),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1583),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1523),
.B(n_985),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1574),
.Y(n_1776)
);

XOR2xp5_ASAP7_75t_L g1777 ( 
.A(n_1616),
.B(n_1327),
.Y(n_1777)
);

CKINVDCx20_ASAP7_75t_R g1778 ( 
.A(n_1486),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1500),
.B(n_1212),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1642),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1589),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1607),
.Y(n_1782)
);

XNOR2x2_ASAP7_75t_L g1783 ( 
.A(n_1487),
.B(n_968),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1501),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1512),
.B(n_1214),
.Y(n_1785)
);

INVx5_ASAP7_75t_L g1786 ( 
.A(n_1630),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1501),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1555),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1557),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1561),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1579),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1565),
.Y(n_1792)
);

CKINVDCx20_ASAP7_75t_R g1793 ( 
.A(n_1508),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1571),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1564),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1572),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1538),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1590),
.A2(n_980),
.B(n_975),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1585),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1524),
.B(n_1026),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1586),
.Y(n_1801)
);

CKINVDCx20_ASAP7_75t_R g1802 ( 
.A(n_1511),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1645),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1668),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1582),
.Y(n_1805)
);

XNOR2x2_ASAP7_75t_L g1806 ( 
.A(n_1487),
.B(n_983),
.Y(n_1806)
);

INVxp67_ASAP7_75t_SL g1807 ( 
.A(n_1591),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1692),
.B(n_1217),
.Y(n_1808)
);

XNOR2x2_ASAP7_75t_L g1809 ( 
.A(n_1495),
.B(n_987),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1584),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1670),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1695),
.B(n_1218),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1584),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1675),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1540),
.B(n_1219),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1543),
.B(n_1220),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1514),
.B(n_1221),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1563),
.B(n_1222),
.Y(n_1818)
);

AOI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1646),
.A2(n_1318),
.B(n_1317),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1504),
.B(n_1349),
.Y(n_1820)
);

AND2x2_ASAP7_75t_SL g1821 ( 
.A(n_1528),
.B(n_1696),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1587),
.B(n_1224),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1623),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1676),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1629),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1634),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1690),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1630),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1544),
.Y(n_1829)
);

XOR2xp5_ASAP7_75t_L g1830 ( 
.A(n_1588),
.B(n_1328),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1644),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1574),
.B(n_988),
.Y(n_1832)
);

INVx2_ASAP7_75t_SL g1833 ( 
.A(n_1578),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1644),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1492),
.Y(n_1835)
);

INVxp33_ASAP7_75t_L g1836 ( 
.A(n_1697),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1617),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1509),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1491),
.B(n_1349),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1551),
.B(n_1226),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1617),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1618),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1516),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1560),
.B(n_1228),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1618),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1624),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1533),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1624),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1667),
.Y(n_1849)
);

CKINVDCx20_ASAP7_75t_R g1850 ( 
.A(n_1663),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1669),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1633),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1679),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1575),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1578),
.B(n_990),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1552),
.Y(n_1856)
);

OAI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1611),
.A2(n_995),
.B(n_994),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1619),
.Y(n_1858)
);

NAND2xp33_ASAP7_75t_R g1859 ( 
.A(n_1531),
.B(n_1621),
.Y(n_1859)
);

CKINVDCx16_ASAP7_75t_R g1860 ( 
.A(n_1581),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1620),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1627),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1628),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1506),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1625),
.B(n_1004),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1506),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1626),
.B(n_1230),
.Y(n_1867)
);

INVxp67_ASAP7_75t_L g1868 ( 
.A(n_1536),
.Y(n_1868)
);

OAI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1573),
.A2(n_1613),
.B(n_1599),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1545),
.Y(n_1870)
);

XNOR2xp5_ASAP7_75t_L g1871 ( 
.A(n_1632),
.B(n_1233),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1593),
.B(n_1234),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1662),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1678),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1680),
.Y(n_1875)
);

BUFx3_ASAP7_75t_L g1876 ( 
.A(n_1592),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1694),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1600),
.B(n_1237),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1686),
.Y(n_1879)
);

CKINVDCx20_ASAP7_75t_R g1880 ( 
.A(n_1602),
.Y(n_1880)
);

CKINVDCx20_ASAP7_75t_R g1881 ( 
.A(n_1638),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1650),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1484),
.B(n_1239),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1659),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1683),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1510),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1513),
.B(n_1349),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1684),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1596),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1687),
.Y(n_1890)
);

NOR2xp67_ASAP7_75t_L g1891 ( 
.A(n_1597),
.B(n_1026),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1688),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1495),
.B(n_1241),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1601),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1502),
.B(n_1349),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1536),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1622),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1608),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1635),
.Y(n_1899)
);

OR2x2_ASAP7_75t_SL g1900 ( 
.A(n_1527),
.B(n_1008),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1636),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1637),
.B(n_1011),
.Y(n_1902)
);

XOR2xp5_ASAP7_75t_L g1903 ( 
.A(n_1532),
.B(n_1329),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1639),
.Y(n_1904)
);

INVxp33_ASAP7_75t_SL g1905 ( 
.A(n_1568),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1568),
.B(n_1249),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1603),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1576),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1529),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1541),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1494),
.B(n_1250),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1547),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1631),
.Y(n_1913)
);

INVxp67_ASAP7_75t_SL g1914 ( 
.A(n_1605),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1640),
.Y(n_1915)
);

NAND2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1660),
.B(n_1013),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1693),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1569),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1570),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1658),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1643),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1654),
.Y(n_1922)
);

CKINVDCx20_ASAP7_75t_R g1923 ( 
.A(n_1653),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1665),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1657),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1661),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1672),
.Y(n_1927)
);

NOR2xp67_ASAP7_75t_L g1928 ( 
.A(n_1649),
.B(n_1027),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1685),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1553),
.B(n_1298),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1652),
.Y(n_1931)
);

BUFx6f_ASAP7_75t_SL g1932 ( 
.A(n_1673),
.Y(n_1932)
);

INVxp67_ASAP7_75t_L g1933 ( 
.A(n_1566),
.Y(n_1933)
);

NAND2xp33_ASAP7_75t_SL g1934 ( 
.A(n_1664),
.B(n_1300),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1671),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1489),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1595),
.B(n_1031),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1554),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1595),
.B(n_1056),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1554),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1689),
.Y(n_1941)
);

INVxp67_ASAP7_75t_SL g1942 ( 
.A(n_1647),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1554),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1503),
.B(n_1303),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1554),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1554),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1554),
.Y(n_1947)
);

CKINVDCx20_ASAP7_75t_R g1948 ( 
.A(n_1522),
.Y(n_1948)
);

INVxp67_ASAP7_75t_SL g1949 ( 
.A(n_1647),
.Y(n_1949)
);

AND2x2_ASAP7_75t_SL g1950 ( 
.A(n_1483),
.B(n_1056),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1483),
.B(n_1251),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1554),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1554),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1549),
.B(n_1252),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1554),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1554),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1483),
.B(n_1257),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1689),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1554),
.Y(n_1959)
);

BUFx6f_ASAP7_75t_L g1960 ( 
.A(n_1538),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1554),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1483),
.B(n_1260),
.Y(n_1962)
);

INVxp33_ASAP7_75t_L g1963 ( 
.A(n_1655),
.Y(n_1963)
);

XOR2x2_ASAP7_75t_L g1964 ( 
.A(n_1530),
.B(n_22),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1689),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1595),
.B(n_1022),
.Y(n_1966)
);

XNOR2xp5_ASAP7_75t_L g1967 ( 
.A(n_1530),
.B(n_1262),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1483),
.B(n_1263),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_SL g1969 ( 
.A(n_1496),
.B(n_1266),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1595),
.B(n_1120),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1595),
.B(n_1023),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1483),
.B(n_1267),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1554),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1554),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1554),
.Y(n_1975)
);

XNOR2xp5_ASAP7_75t_L g1976 ( 
.A(n_1530),
.B(n_1268),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1554),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1549),
.B(n_1270),
.Y(n_1978)
);

INVx2_ASAP7_75t_SL g1979 ( 
.A(n_1518),
.Y(n_1979)
);

INVx2_ASAP7_75t_SL g1980 ( 
.A(n_1518),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1554),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1595),
.B(n_1120),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1554),
.Y(n_1983)
);

INVxp33_ASAP7_75t_L g1984 ( 
.A(n_1655),
.Y(n_1984)
);

XNOR2x2_ASAP7_75t_L g1985 ( 
.A(n_1485),
.B(n_1035),
.Y(n_1985)
);

OR2x6_ASAP7_75t_L g1986 ( 
.A(n_1498),
.B(n_1164),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1554),
.Y(n_1987)
);

XNOR2xp5_ASAP7_75t_L g1988 ( 
.A(n_1530),
.B(n_1271),
.Y(n_1988)
);

BUFx8_ASAP7_75t_L g1989 ( 
.A(n_1496),
.Y(n_1989)
);

CKINVDCx16_ASAP7_75t_R g1990 ( 
.A(n_1498),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1554),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1554),
.Y(n_1992)
);

INVx3_ASAP7_75t_L g1993 ( 
.A(n_1786),
.Y(n_1993)
);

INVx2_ASAP7_75t_SL g1994 ( 
.A(n_1979),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1731),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1950),
.B(n_1272),
.Y(n_1996)
);

OAI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1887),
.A2(n_1037),
.B(n_1036),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1770),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1930),
.B(n_1919),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1807),
.B(n_1273),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1805),
.B(n_1043),
.Y(n_2001)
);

OAI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1887),
.A2(n_1046),
.B(n_1044),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1714),
.B(n_1275),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1743),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1715),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1698),
.B(n_1277),
.Y(n_2006)
);

BUFx3_ASAP7_75t_L g2007 ( 
.A(n_1742),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1836),
.B(n_1279),
.Y(n_2008)
);

BUFx6f_ASAP7_75t_L g2009 ( 
.A(n_1786),
.Y(n_2009)
);

AND2x4_ASAP7_75t_SL g2010 ( 
.A(n_1755),
.B(n_1164),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1719),
.B(n_1280),
.Y(n_2011)
);

INVx2_ASAP7_75t_SL g2012 ( 
.A(n_1980),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1723),
.B(n_1282),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1951),
.B(n_1283),
.Y(n_2014)
);

INVx3_ASAP7_75t_L g2015 ( 
.A(n_1786),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1902),
.Y(n_2016)
);

BUFx6f_ASAP7_75t_L g2017 ( 
.A(n_1718),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1876),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1727),
.B(n_1285),
.Y(n_2019)
);

OAI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1820),
.A2(n_1048),
.B(n_1047),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1902),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1774),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1712),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1861),
.Y(n_2024)
);

INVxp67_ASAP7_75t_L g2025 ( 
.A(n_1734),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_1810),
.B(n_1050),
.Y(n_2026)
);

INVx1_ASAP7_75t_SL g2027 ( 
.A(n_1722),
.Y(n_2027)
);

AND2x4_ASAP7_75t_SL g2028 ( 
.A(n_1755),
.B(n_1171),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1742),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1941),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1862),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1958),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1965),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_L g2034 ( 
.A(n_1718),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1722),
.B(n_1286),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1728),
.B(n_1287),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1863),
.Y(n_2037)
);

HB1xp67_ASAP7_75t_L g2038 ( 
.A(n_1720),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1716),
.B(n_1288),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1725),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1813),
.B(n_1051),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1717),
.Y(n_2042)
);

INVxp33_ASAP7_75t_L g2043 ( 
.A(n_1830),
.Y(n_2043)
);

OAI21x1_ASAP7_75t_L g2044 ( 
.A1(n_1819),
.A2(n_1215),
.B(n_1171),
.Y(n_2044)
);

INVx2_ASAP7_75t_SL g2045 ( 
.A(n_1755),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1966),
.B(n_1289),
.Y(n_2046)
);

INVxp67_ASAP7_75t_L g2047 ( 
.A(n_1942),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1699),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_1966),
.B(n_1052),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1957),
.B(n_1290),
.Y(n_2050)
);

BUFx4f_ASAP7_75t_L g2051 ( 
.A(n_1986),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1971),
.B(n_1291),
.Y(n_2052)
);

INVxp67_ASAP7_75t_SL g2053 ( 
.A(n_1949),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_1725),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1971),
.B(n_1749),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1889),
.Y(n_2056)
);

AND2x2_ASAP7_75t_SL g2057 ( 
.A(n_1990),
.B(n_1215),
.Y(n_2057)
);

BUFx6f_ASAP7_75t_L g2058 ( 
.A(n_1718),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1962),
.B(n_1292),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1703),
.Y(n_2060)
);

INVx4_ASAP7_75t_L g2061 ( 
.A(n_1986),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1760),
.B(n_1294),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1704),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1938),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1968),
.B(n_1295),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1940),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1960),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1853),
.B(n_1296),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1784),
.B(n_1054),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1798),
.B(n_1304),
.Y(n_2070)
);

HB1xp67_ASAP7_75t_L g2071 ( 
.A(n_1739),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1894),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1898),
.Y(n_2073)
);

AND2x2_ASAP7_75t_SL g2074 ( 
.A(n_1969),
.B(n_1265),
.Y(n_2074)
);

INVx2_ASAP7_75t_SL g2075 ( 
.A(n_1730),
.Y(n_2075)
);

HB1xp67_ASAP7_75t_L g2076 ( 
.A(n_1739),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1972),
.B(n_1305),
.Y(n_2077)
);

INVx3_ASAP7_75t_L g2078 ( 
.A(n_1803),
.Y(n_2078)
);

BUFx6f_ASAP7_75t_L g2079 ( 
.A(n_1960),
.Y(n_2079)
);

INVx1_ASAP7_75t_SL g2080 ( 
.A(n_1738),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1933),
.B(n_1306),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1943),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1960),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1945),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_L g2085 ( 
.A(n_1700),
.B(n_1307),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1798),
.B(n_1772),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1771),
.B(n_1309),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1804),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1946),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1702),
.B(n_1893),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1947),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1787),
.B(n_1057),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1944),
.B(n_1323),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1733),
.B(n_1330),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1811),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1753),
.B(n_1334),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1808),
.B(n_1075),
.Y(n_2097)
);

OAI21xp5_ASAP7_75t_L g2098 ( 
.A1(n_1820),
.A2(n_1081),
.B(n_1078),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1952),
.Y(n_2099)
);

INVx1_ASAP7_75t_SL g2100 ( 
.A(n_1745),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1732),
.B(n_1083),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_L g2102 ( 
.A(n_1776),
.B(n_1256),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1735),
.B(n_1086),
.Y(n_2103)
);

NAND2x1p5_ASAP7_75t_L g2104 ( 
.A(n_1705),
.B(n_1265),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1812),
.B(n_1102),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1953),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_1795),
.B(n_1106),
.Y(n_2107)
);

INVxp67_ASAP7_75t_SL g2108 ( 
.A(n_1916),
.Y(n_2108)
);

INVx2_ASAP7_75t_SL g2109 ( 
.A(n_1989),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1955),
.Y(n_2110)
);

BUFx2_ASAP7_75t_L g2111 ( 
.A(n_1989),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1882),
.B(n_1107),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1956),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1959),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_1796),
.B(n_1108),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1814),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1884),
.B(n_1109),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1906),
.B(n_1113),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_1911),
.B(n_1116),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1914),
.B(n_1123),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1961),
.Y(n_2121)
);

OAI21xp5_ASAP7_75t_L g2122 ( 
.A1(n_1839),
.A2(n_1126),
.B(n_1125),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1916),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1885),
.B(n_1128),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1888),
.B(n_1130),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1973),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1974),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1890),
.B(n_1132),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1824),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1827),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_1903),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1899),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_1969),
.B(n_1134),
.Y(n_2133)
);

INVxp67_ASAP7_75t_L g2134 ( 
.A(n_1832),
.Y(n_2134)
);

NAND2x1p5_ASAP7_75t_L g2135 ( 
.A(n_1706),
.B(n_1137),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_1832),
.B(n_1153),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1901),
.Y(n_2137)
);

BUFx6f_ASAP7_75t_L g2138 ( 
.A(n_1708),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1872),
.B(n_1156),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_1878),
.B(n_1157),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1710),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1975),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1892),
.B(n_1158),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_1743),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1762),
.B(n_1159),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_SL g2146 ( 
.A(n_1837),
.B(n_1841),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1977),
.Y(n_2147)
);

INVx3_ASAP7_75t_L g2148 ( 
.A(n_1907),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1748),
.B(n_1160),
.Y(n_2149)
);

OR2x6_ASAP7_75t_L g2150 ( 
.A(n_1986),
.B(n_1165),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1748),
.B(n_1166),
.Y(n_2151)
);

OAI21xp5_ASAP7_75t_L g2152 ( 
.A1(n_1839),
.A2(n_1176),
.B(n_1168),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1777),
.B(n_1178),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1981),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1937),
.B(n_1982),
.Y(n_2155)
);

AND2x4_ASAP7_75t_L g2156 ( 
.A(n_1799),
.B(n_1181),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_1897),
.B(n_1247),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_L g2158 ( 
.A(n_1833),
.B(n_1248),
.Y(n_2158)
);

INVx3_ASAP7_75t_L g2159 ( 
.A(n_1788),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1937),
.B(n_1191),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1939),
.B(n_1196),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1939),
.B(n_1209),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1983),
.Y(n_2163)
);

BUFx6f_ASAP7_75t_L g2164 ( 
.A(n_1711),
.Y(n_2164)
);

BUFx6f_ASAP7_75t_L g2165 ( 
.A(n_1713),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1970),
.B(n_1210),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1904),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1789),
.Y(n_2168)
);

HB1xp67_ASAP7_75t_L g2169 ( 
.A(n_1756),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_1855),
.B(n_1737),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1970),
.B(n_1211),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_1855),
.B(n_1747),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1987),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1982),
.B(n_1213),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_1817),
.B(n_1216),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1857),
.B(n_1225),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1991),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1769),
.B(n_1231),
.Y(n_2178)
);

OAI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_1895),
.A2(n_1240),
.B(n_1232),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1857),
.B(n_1242),
.Y(n_2180)
);

BUFx4f_ASAP7_75t_L g2181 ( 
.A(n_1920),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1992),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1769),
.B(n_1246),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1790),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1791),
.Y(n_2185)
);

BUFx3_ASAP7_75t_L g2186 ( 
.A(n_1746),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1752),
.B(n_1757),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_1865),
.B(n_1253),
.Y(n_2188)
);

AOI22xp5_ASAP7_75t_L g2189 ( 
.A1(n_1821),
.A2(n_1259),
.B1(n_1269),
.B2(n_1254),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1801),
.Y(n_2190)
);

OAI21xp5_ASAP7_75t_L g2191 ( 
.A1(n_1895),
.A2(n_1278),
.B(n_1274),
.Y(n_2191)
);

BUFx2_ASAP7_75t_L g2192 ( 
.A(n_1936),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1792),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_1900),
.B(n_1910),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1794),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_1852),
.B(n_1281),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1823),
.Y(n_2197)
);

INVx3_ASAP7_75t_L g2198 ( 
.A(n_1759),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1780),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1825),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_1865),
.B(n_1293),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_1779),
.B(n_1297),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1764),
.B(n_1301),
.Y(n_2203)
);

AND2x4_ASAP7_75t_L g2204 ( 
.A(n_1826),
.B(n_1316),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_1854),
.B(n_23),
.Y(n_2205)
);

INVx3_ASAP7_75t_L g2206 ( 
.A(n_1828),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_L g2207 ( 
.A(n_1765),
.B(n_23),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1764),
.B(n_840),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_1709),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1891),
.Y(n_2210)
);

AND2x4_ASAP7_75t_L g2211 ( 
.A(n_1908),
.B(n_24),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1835),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1724),
.B(n_1909),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_1729),
.B(n_841),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1724),
.B(n_841),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1912),
.B(n_25),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1869),
.B(n_25),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1868),
.B(n_824),
.Y(n_2218)
);

HB1xp67_ASAP7_75t_L g2219 ( 
.A(n_1768),
.Y(n_2219)
);

BUFx3_ASAP7_75t_L g2220 ( 
.A(n_1751),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1891),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1838),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1869),
.B(n_824),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_1868),
.B(n_825),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_L g2225 ( 
.A(n_1815),
.B(n_1816),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_1831),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1918),
.B(n_1726),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_1834),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1913),
.B(n_825),
.Y(n_2229)
);

OR2x2_ASAP7_75t_SL g2230 ( 
.A(n_1860),
.B(n_26),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1915),
.B(n_826),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1843),
.Y(n_2232)
);

BUFx6f_ASAP7_75t_L g2233 ( 
.A(n_1842),
.Y(n_2233)
);

OAI21xp5_ASAP7_75t_L g2234 ( 
.A1(n_1758),
.A2(n_1800),
.B(n_1775),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_L g2235 ( 
.A(n_1845),
.Y(n_2235)
);

HB1xp67_ASAP7_75t_L g2236 ( 
.A(n_1964),
.Y(n_2236)
);

INVx2_ASAP7_75t_SL g2237 ( 
.A(n_1858),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_1707),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_1740),
.B(n_827),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1849),
.B(n_827),
.Y(n_2240)
);

BUFx3_ASAP7_75t_L g2241 ( 
.A(n_1781),
.Y(n_2241)
);

OR2x2_ASAP7_75t_L g2242 ( 
.A(n_1744),
.B(n_828),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1761),
.Y(n_2243)
);

BUFx4f_ASAP7_75t_L g2244 ( 
.A(n_1886),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1851),
.B(n_829),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1847),
.Y(n_2246)
);

BUFx6f_ASAP7_75t_L g2247 ( 
.A(n_1846),
.Y(n_2247)
);

OAI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_1758),
.A2(n_26),
.B(n_27),
.Y(n_2248)
);

HB1xp67_ASAP7_75t_L g2249 ( 
.A(n_1967),
.Y(n_2249)
);

INVx4_ASAP7_75t_L g2250 ( 
.A(n_1932),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1763),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_1840),
.B(n_1844),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_1883),
.B(n_830),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1848),
.B(n_830),
.Y(n_2254)
);

INVx4_ASAP7_75t_L g2255 ( 
.A(n_1932),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1773),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_1924),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_1818),
.B(n_831),
.Y(n_2258)
);

INVx1_ASAP7_75t_SL g2259 ( 
.A(n_1923),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_1976),
.B(n_831),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_1988),
.B(n_832),
.Y(n_2261)
);

BUFx6f_ASAP7_75t_L g2262 ( 
.A(n_1797),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_1917),
.B(n_1721),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1782),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_1822),
.B(n_834),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_1867),
.B(n_27),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_1954),
.B(n_835),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_1978),
.B(n_835),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_1785),
.B(n_28),
.Y(n_2269)
);

INVx3_ASAP7_75t_L g2270 ( 
.A(n_1873),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1874),
.B(n_837),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1856),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_1875),
.B(n_838),
.Y(n_2273)
);

INVx4_ASAP7_75t_L g2274 ( 
.A(n_1767),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_1750),
.B(n_28),
.Y(n_2275)
);

HB1xp67_ASAP7_75t_L g2276 ( 
.A(n_1783),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1879),
.B(n_840),
.Y(n_2277)
);

INVx2_ASAP7_75t_SL g2278 ( 
.A(n_1871),
.Y(n_2278)
);

BUFx3_ASAP7_75t_L g2279 ( 
.A(n_1850),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1864),
.Y(n_2280)
);

HB1xp67_ASAP7_75t_L g2281 ( 
.A(n_1806),
.Y(n_2281)
);

HB1xp67_ASAP7_75t_L g2282 ( 
.A(n_1809),
.Y(n_2282)
);

INVx3_ASAP7_75t_L g2283 ( 
.A(n_1877),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_1793),
.B(n_29),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1921),
.Y(n_2285)
);

INVx4_ASAP7_75t_L g2286 ( 
.A(n_1767),
.Y(n_2286)
);

OAI21xp5_ASAP7_75t_L g2287 ( 
.A1(n_1766),
.A2(n_29),
.B(n_30),
.Y(n_2287)
);

INVx3_ASAP7_75t_L g2288 ( 
.A(n_1866),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_1802),
.B(n_811),
.Y(n_2289)
);

AND2x6_ASAP7_75t_L g2290 ( 
.A(n_1896),
.B(n_30),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_1922),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1925),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_L g2293 ( 
.A(n_1880),
.B(n_31),
.Y(n_2293)
);

INVxp67_ASAP7_75t_L g2294 ( 
.A(n_1934),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_1778),
.B(n_1829),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1928),
.Y(n_2296)
);

BUFx4f_ASAP7_75t_L g2297 ( 
.A(n_1859),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1928),
.Y(n_2298)
);

INVx2_ASAP7_75t_SL g2299 ( 
.A(n_1985),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_1926),
.B(n_813),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1927),
.Y(n_2301)
);

BUFx6f_ASAP7_75t_L g2302 ( 
.A(n_1929),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1870),
.B(n_813),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1905),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_1741),
.B(n_814),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1931),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_1754),
.B(n_815),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1935),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_1881),
.Y(n_2309)
);

INVx2_ASAP7_75t_SL g2310 ( 
.A(n_1701),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_1948),
.Y(n_2311)
);

OAI21xp5_ASAP7_75t_L g2312 ( 
.A1(n_1963),
.A2(n_32),
.B(n_33),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_1736),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1984),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1770),
.Y(n_2315)
);

INVx3_ASAP7_75t_L g2316 ( 
.A(n_1786),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_1807),
.B(n_817),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_1950),
.B(n_817),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_1807),
.B(n_818),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1715),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_1950),
.B(n_818),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1807),
.B(n_819),
.Y(n_2322)
);

BUFx6f_ASAP7_75t_L g2323 ( 
.A(n_1786),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_1836),
.B(n_32),
.Y(n_2324)
);

INVx3_ASAP7_75t_L g2325 ( 
.A(n_1786),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_1807),
.B(n_820),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_1770),
.Y(n_2327)
);

AND2x2_ASAP7_75t_SL g2328 ( 
.A(n_1990),
.B(n_34),
.Y(n_2328)
);

HB1xp67_ASAP7_75t_L g2329 ( 
.A(n_1720),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_1836),
.B(n_34),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1715),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1715),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_1770),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_L g2334 ( 
.A(n_2225),
.B(n_821),
.Y(n_2334)
);

INVxp67_ASAP7_75t_L g2335 ( 
.A(n_2187),
.Y(n_2335)
);

INVxp67_ASAP7_75t_L g2336 ( 
.A(n_2187),
.Y(n_2336)
);

INVx5_ASAP7_75t_L g2337 ( 
.A(n_2009),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_SL g2338 ( 
.A(n_2051),
.B(n_36),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2155),
.B(n_2023),
.Y(n_2339)
);

INVx4_ASAP7_75t_L g2340 ( 
.A(n_2009),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_L g2341 ( 
.A(n_2134),
.B(n_821),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2193),
.Y(n_2342)
);

BUFx6f_ASAP7_75t_L g2343 ( 
.A(n_2017),
.Y(n_2343)
);

AND2x4_ASAP7_75t_L g2344 ( 
.A(n_2108),
.B(n_36),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2155),
.B(n_37),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_2045),
.B(n_37),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2030),
.B(n_38),
.Y(n_2347)
);

AND2x4_ASAP7_75t_L g2348 ( 
.A(n_2061),
.B(n_38),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_2061),
.B(n_39),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2145),
.B(n_2093),
.Y(n_2350)
);

INVx4_ASAP7_75t_L g2351 ( 
.A(n_2009),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2032),
.B(n_2033),
.Y(n_2352)
);

OR2x6_ASAP7_75t_L g2353 ( 
.A(n_2007),
.B(n_41),
.Y(n_2353)
);

BUFx3_ASAP7_75t_L g2354 ( 
.A(n_2029),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2194),
.B(n_41),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2195),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2042),
.Y(n_2357)
);

BUFx6f_ASAP7_75t_L g2358 ( 
.A(n_2017),
.Y(n_2358)
);

BUFx6f_ASAP7_75t_L g2359 ( 
.A(n_2017),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2189),
.B(n_42),
.Y(n_2360)
);

NAND2x1p5_ASAP7_75t_L g2361 ( 
.A(n_2051),
.B(n_44),
.Y(n_2361)
);

NAND2x1p5_ASAP7_75t_L g2362 ( 
.A(n_2111),
.B(n_44),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2138),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_2134),
.B(n_42),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2048),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2055),
.B(n_45),
.Y(n_2366)
);

BUFx12f_ASAP7_75t_L g2367 ( 
.A(n_2109),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2138),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2060),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2055),
.B(n_45),
.Y(n_2370)
);

AO21x2_ASAP7_75t_L g2371 ( 
.A1(n_2217),
.A2(n_46),
.B(n_47),
.Y(n_2371)
);

CKINVDCx11_ASAP7_75t_R g2372 ( 
.A(n_2192),
.Y(n_2372)
);

BUFx8_ASAP7_75t_L g2373 ( 
.A(n_2220),
.Y(n_2373)
);

AND2x2_ASAP7_75t_SL g2374 ( 
.A(n_2074),
.B(n_46),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2003),
.B(n_49),
.Y(n_2375)
);

NAND2x1p5_ASAP7_75t_L g2376 ( 
.A(n_2323),
.B(n_51),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2120),
.B(n_50),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2252),
.B(n_811),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2081),
.B(n_50),
.Y(n_2379)
);

BUFx2_ASAP7_75t_SL g2380 ( 
.A(n_2123),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2227),
.B(n_51),
.Y(n_2381)
);

BUFx4f_ASAP7_75t_L g2382 ( 
.A(n_2150),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2170),
.B(n_52),
.Y(n_2383)
);

CKINVDCx6p67_ASAP7_75t_R g2384 ( 
.A(n_2150),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2227),
.B(n_52),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2119),
.B(n_53),
.Y(n_2386)
);

INVx6_ASAP7_75t_L g2387 ( 
.A(n_2323),
.Y(n_2387)
);

AND2x4_ASAP7_75t_L g2388 ( 
.A(n_2274),
.B(n_53),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2063),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2068),
.B(n_54),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_SL g2391 ( 
.A(n_1995),
.B(n_54),
.Y(n_2391)
);

NAND2xp33_ASAP7_75t_L g2392 ( 
.A(n_2034),
.B(n_55),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2064),
.Y(n_2393)
);

BUFx6f_ASAP7_75t_L g2394 ( 
.A(n_2034),
.Y(n_2394)
);

BUFx3_ASAP7_75t_L g2395 ( 
.A(n_2186),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2066),
.Y(n_2396)
);

BUFx2_ASAP7_75t_L g2397 ( 
.A(n_2150),
.Y(n_2397)
);

AND2x6_ASAP7_75t_L g2398 ( 
.A(n_2123),
.B(n_56),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2082),
.Y(n_2399)
);

BUFx8_ASAP7_75t_SL g2400 ( 
.A(n_2004),
.Y(n_2400)
);

BUFx4f_ASAP7_75t_L g2401 ( 
.A(n_2328),
.Y(n_2401)
);

AND2x2_ASAP7_75t_SL g2402 ( 
.A(n_2057),
.B(n_56),
.Y(n_2402)
);

NAND2x1p5_ASAP7_75t_L g2403 ( 
.A(n_2323),
.B(n_59),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2172),
.B(n_57),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2138),
.Y(n_2405)
);

AND2x4_ASAP7_75t_L g2406 ( 
.A(n_2274),
.B(n_57),
.Y(n_2406)
);

BUFx4f_ASAP7_75t_L g2407 ( 
.A(n_2290),
.Y(n_2407)
);

CKINVDCx8_ASAP7_75t_R g2408 ( 
.A(n_2144),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2068),
.B(n_60),
.Y(n_2409)
);

AND2x4_ASAP7_75t_L g2410 ( 
.A(n_2286),
.B(n_2075),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_2034),
.Y(n_2411)
);

OR2x2_ASAP7_75t_L g2412 ( 
.A(n_2259),
.B(n_1999),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2084),
.B(n_61),
.Y(n_2413)
);

BUFx6f_ASAP7_75t_L g2414 ( 
.A(n_2058),
.Y(n_2414)
);

AND2x4_ASAP7_75t_L g2415 ( 
.A(n_2286),
.B(n_62),
.Y(n_2415)
);

BUFx3_ASAP7_75t_L g2416 ( 
.A(n_2038),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_2089),
.B(n_64),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2091),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2153),
.B(n_65),
.Y(n_2419)
);

INVxp67_ASAP7_75t_L g2420 ( 
.A(n_2211),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_2123),
.B(n_65),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_SL g2422 ( 
.A(n_2297),
.B(n_66),
.Y(n_2422)
);

INVx4_ASAP7_75t_L g2423 ( 
.A(n_2058),
.Y(n_2423)
);

INVx5_ASAP7_75t_L g2424 ( 
.A(n_2058),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2099),
.B(n_67),
.Y(n_2425)
);

BUFx4f_ASAP7_75t_L g2426 ( 
.A(n_2290),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2141),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_2106),
.B(n_68),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2087),
.B(n_2090),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2008),
.B(n_812),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2284),
.B(n_2289),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2110),
.B(n_68),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2113),
.Y(n_2433)
);

AND2x4_ASAP7_75t_L g2434 ( 
.A(n_2114),
.B(n_69),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2121),
.B(n_69),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_SL g2436 ( 
.A(n_2297),
.B(n_2250),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2126),
.B(n_70),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2141),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2127),
.B(n_70),
.Y(n_2439)
);

BUFx4f_ASAP7_75t_L g2440 ( 
.A(n_2290),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2006),
.B(n_72),
.Y(n_2441)
);

INVx3_ASAP7_75t_L g2442 ( 
.A(n_1993),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2309),
.B(n_822),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2142),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2147),
.Y(n_2445)
);

BUFx6f_ASAP7_75t_L g2446 ( 
.A(n_2067),
.Y(n_2446)
);

OR2x6_ASAP7_75t_L g2447 ( 
.A(n_2250),
.B(n_72),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2014),
.B(n_73),
.Y(n_2448)
);

BUFx6f_ASAP7_75t_L g2449 ( 
.A(n_2067),
.Y(n_2449)
);

AND2x4_ASAP7_75t_L g2450 ( 
.A(n_2154),
.B(n_74),
.Y(n_2450)
);

INVx1_ASAP7_75t_SL g2451 ( 
.A(n_2010),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2163),
.Y(n_2452)
);

NOR2xp33_ASAP7_75t_L g2453 ( 
.A(n_2304),
.B(n_834),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2173),
.B(n_74),
.Y(n_2454)
);

AND2x4_ASAP7_75t_L g2455 ( 
.A(n_2177),
.B(n_75),
.Y(n_2455)
);

CKINVDCx6p67_ASAP7_75t_R g2456 ( 
.A(n_2279),
.Y(n_2456)
);

BUFx6f_ASAP7_75t_L g2457 ( 
.A(n_2067),
.Y(n_2457)
);

AND2x6_ASAP7_75t_L g2458 ( 
.A(n_2211),
.B(n_75),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2182),
.B(n_76),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2086),
.B(n_76),
.Y(n_2460)
);

BUFx2_ASAP7_75t_SL g2461 ( 
.A(n_2079),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2016),
.Y(n_2462)
);

AND2x2_ASAP7_75t_SL g2463 ( 
.A(n_2205),
.B(n_77),
.Y(n_2463)
);

OR2x2_ASAP7_75t_L g2464 ( 
.A(n_2259),
.B(n_77),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2141),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2164),
.Y(n_2466)
);

OR2x2_ASAP7_75t_L g2467 ( 
.A(n_2131),
.B(n_78),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2050),
.B(n_78),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2086),
.B(n_2157),
.Y(n_2469)
);

HB1xp67_ASAP7_75t_L g2470 ( 
.A(n_2329),
.Y(n_2470)
);

OR2x2_ASAP7_75t_L g2471 ( 
.A(n_2219),
.B(n_79),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2097),
.B(n_80),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2105),
.B(n_81),
.Y(n_2473)
);

BUFx2_ASAP7_75t_L g2474 ( 
.A(n_2040),
.Y(n_2474)
);

NOR2xp67_ASAP7_75t_L g2475 ( 
.A(n_2255),
.B(n_82),
.Y(n_2475)
);

INVx5_ASAP7_75t_L g2476 ( 
.A(n_2079),
.Y(n_2476)
);

BUFx3_ASAP7_75t_L g2477 ( 
.A(n_2198),
.Y(n_2477)
);

AND2x6_ASAP7_75t_L g2478 ( 
.A(n_2205),
.B(n_83),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2118),
.B(n_83),
.Y(n_2479)
);

INVxp67_ASAP7_75t_L g2480 ( 
.A(n_2094),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2021),
.Y(n_2481)
);

NOR2xp67_ASAP7_75t_L g2482 ( 
.A(n_2255),
.B(n_86),
.Y(n_2482)
);

AND2x4_ASAP7_75t_L g2483 ( 
.A(n_2005),
.B(n_86),
.Y(n_2483)
);

AND2x4_ASAP7_75t_L g2484 ( 
.A(n_2320),
.B(n_87),
.Y(n_2484)
);

AND2x4_ASAP7_75t_L g2485 ( 
.A(n_2331),
.B(n_87),
.Y(n_2485)
);

INVx4_ASAP7_75t_L g2486 ( 
.A(n_2079),
.Y(n_2486)
);

NAND2x1p5_ASAP7_75t_L g2487 ( 
.A(n_1993),
.B(n_2015),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2139),
.B(n_88),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2059),
.B(n_89),
.Y(n_2489)
);

NAND2x1p5_ASAP7_75t_L g2490 ( 
.A(n_2015),
.B(n_93),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2140),
.B(n_91),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_SL g2492 ( 
.A(n_2027),
.B(n_91),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2070),
.B(n_95),
.Y(n_2493)
);

CKINVDCx8_ASAP7_75t_R g2494 ( 
.A(n_2290),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2164),
.Y(n_2495)
);

INVxp67_ASAP7_75t_L g2496 ( 
.A(n_2096),
.Y(n_2496)
);

BUFx3_ASAP7_75t_L g2497 ( 
.A(n_2198),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2190),
.Y(n_2498)
);

OR2x6_ASAP7_75t_L g2499 ( 
.A(n_1994),
.B(n_2012),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2070),
.B(n_95),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2332),
.Y(n_2501)
);

CKINVDCx11_ASAP7_75t_R g2502 ( 
.A(n_2314),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2164),
.Y(n_2503)
);

INVxp67_ASAP7_75t_L g2504 ( 
.A(n_2065),
.Y(n_2504)
);

NOR2xp33_ASAP7_75t_L g2505 ( 
.A(n_1996),
.B(n_2077),
.Y(n_2505)
);

OR2x2_ASAP7_75t_L g2506 ( 
.A(n_2295),
.B(n_97),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2318),
.B(n_97),
.Y(n_2507)
);

AND2x4_ASAP7_75t_L g2508 ( 
.A(n_2270),
.B(n_99),
.Y(n_2508)
);

BUFx4f_ASAP7_75t_L g2509 ( 
.A(n_2028),
.Y(n_2509)
);

INVx2_ASAP7_75t_SL g2510 ( 
.A(n_2244),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2197),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2270),
.B(n_99),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2175),
.B(n_100),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2069),
.B(n_101),
.Y(n_2514)
);

INVx2_ASAP7_75t_SL g2515 ( 
.A(n_2244),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2243),
.Y(n_2516)
);

BUFx6f_ASAP7_75t_L g2517 ( 
.A(n_2083),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2069),
.B(n_101),
.Y(n_2518)
);

AND2x4_ASAP7_75t_L g2519 ( 
.A(n_2200),
.B(n_102),
.Y(n_2519)
);

BUFx12f_ASAP7_75t_L g2520 ( 
.A(n_2230),
.Y(n_2520)
);

OR2x2_ASAP7_75t_L g2521 ( 
.A(n_2062),
.B(n_102),
.Y(n_2521)
);

BUFx2_ASAP7_75t_L g2522 ( 
.A(n_2054),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2165),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2092),
.B(n_103),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2251),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2083),
.Y(n_2526)
);

BUFx6f_ASAP7_75t_L g2527 ( 
.A(n_2083),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2165),
.Y(n_2528)
);

AND2x4_ASAP7_75t_L g2529 ( 
.A(n_2316),
.B(n_104),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2165),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2024),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2233),
.Y(n_2532)
);

NOR2xp33_ASAP7_75t_SL g2533 ( 
.A(n_2027),
.B(n_106),
.Y(n_2533)
);

AND2x4_ASAP7_75t_L g2534 ( 
.A(n_2316),
.B(n_106),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2233),
.Y(n_2535)
);

AND2x2_ASAP7_75t_SL g2536 ( 
.A(n_2321),
.B(n_107),
.Y(n_2536)
);

BUFx3_ASAP7_75t_L g2537 ( 
.A(n_2148),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2188),
.B(n_107),
.Y(n_2538)
);

NAND2x1p5_ASAP7_75t_L g2539 ( 
.A(n_2325),
.B(n_109),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2031),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2201),
.B(n_2207),
.Y(n_2541)
);

AND2x4_ASAP7_75t_L g2542 ( 
.A(n_2325),
.B(n_108),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2092),
.B(n_108),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2202),
.B(n_2000),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2037),
.Y(n_2545)
);

BUFx3_ASAP7_75t_L g2546 ( 
.A(n_2148),
.Y(n_2546)
);

AND2x4_ASAP7_75t_L g2547 ( 
.A(n_2237),
.B(n_109),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2000),
.B(n_110),
.Y(n_2548)
);

OR2x6_ASAP7_75t_L g2549 ( 
.A(n_2310),
.B(n_111),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2049),
.B(n_111),
.Y(n_2550)
);

BUFx6f_ASAP7_75t_L g2551 ( 
.A(n_2257),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2233),
.Y(n_2552)
);

INVx1_ASAP7_75t_SL g2553 ( 
.A(n_2242),
.Y(n_2553)
);

BUFx2_ASAP7_75t_SL g2554 ( 
.A(n_2071),
.Y(n_2554)
);

AND2x4_ASAP7_75t_L g2555 ( 
.A(n_2206),
.B(n_112),
.Y(n_2555)
);

OR2x6_ASAP7_75t_L g2556 ( 
.A(n_2209),
.B(n_112),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2049),
.B(n_113),
.Y(n_2557)
);

AND2x6_ASAP7_75t_L g2558 ( 
.A(n_2235),
.B(n_114),
.Y(n_2558)
);

BUFx3_ASAP7_75t_L g2559 ( 
.A(n_2241),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2168),
.Y(n_2560)
);

NAND2x1p5_ASAP7_75t_L g2561 ( 
.A(n_2018),
.B(n_116),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2062),
.B(n_115),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2235),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2136),
.B(n_115),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2203),
.B(n_116),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2203),
.B(n_117),
.Y(n_2566)
);

INVx5_ASAP7_75t_L g2567 ( 
.A(n_2018),
.Y(n_2567)
);

AND2x4_ASAP7_75t_L g2568 ( 
.A(n_2206),
.B(n_117),
.Y(n_2568)
);

NAND2x1p5_ASAP7_75t_L g2569 ( 
.A(n_2133),
.B(n_119),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2112),
.B(n_2117),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2112),
.B(n_118),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2235),
.Y(n_2572)
);

NAND2x1_ASAP7_75t_L g2573 ( 
.A(n_2247),
.B(n_2283),
.Y(n_2573)
);

BUFx6f_ASAP7_75t_L g2574 ( 
.A(n_2257),
.Y(n_2574)
);

BUFx6f_ASAP7_75t_L g2575 ( 
.A(n_2257),
.Y(n_2575)
);

BUFx10_ASAP7_75t_L g2576 ( 
.A(n_2196),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2088),
.Y(n_2577)
);

INVx5_ASAP7_75t_L g2578 ( 
.A(n_2302),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2085),
.B(n_119),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2095),
.Y(n_2580)
);

AND2x4_ASAP7_75t_L g2581 ( 
.A(n_2226),
.B(n_120),
.Y(n_2581)
);

AND2x4_ASAP7_75t_L g2582 ( 
.A(n_2226),
.B(n_121),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2116),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2117),
.B(n_122),
.Y(n_2584)
);

NOR2x1p5_ASAP7_75t_L g2585 ( 
.A(n_2313),
.B(n_124),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2247),
.Y(n_2586)
);

OR2x2_ASAP7_75t_L g2587 ( 
.A(n_2046),
.B(n_2052),
.Y(n_2587)
);

AND2x4_ASAP7_75t_L g2588 ( 
.A(n_2228),
.B(n_126),
.Y(n_2588)
);

BUFx3_ASAP7_75t_L g2589 ( 
.A(n_2078),
.Y(n_2589)
);

BUFx12f_ASAP7_75t_L g2590 ( 
.A(n_2278),
.Y(n_2590)
);

NOR2xp33_ASAP7_75t_SL g2591 ( 
.A(n_2311),
.B(n_127),
.Y(n_2591)
);

AND2x4_ASAP7_75t_L g2592 ( 
.A(n_2228),
.B(n_128),
.Y(n_2592)
);

BUFx2_ASAP7_75t_L g2593 ( 
.A(n_2076),
.Y(n_2593)
);

OR2x6_ASAP7_75t_L g2594 ( 
.A(n_2312),
.B(n_128),
.Y(n_2594)
);

OR2x2_ASAP7_75t_L g2595 ( 
.A(n_2046),
.B(n_129),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2263),
.B(n_129),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2238),
.Y(n_2597)
);

HB1xp67_ASAP7_75t_L g2598 ( 
.A(n_2025),
.Y(n_2598)
);

HB1xp67_ASAP7_75t_L g2599 ( 
.A(n_2025),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2129),
.Y(n_2600)
);

BUFx2_ASAP7_75t_L g2601 ( 
.A(n_2053),
.Y(n_2601)
);

NAND2x1p5_ASAP7_75t_L g2602 ( 
.A(n_2159),
.B(n_131),
.Y(n_2602)
);

NOR2xp33_ASAP7_75t_L g2603 ( 
.A(n_2052),
.B(n_823),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2124),
.B(n_130),
.Y(n_2604)
);

BUFx3_ASAP7_75t_L g2605 ( 
.A(n_2078),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2178),
.B(n_131),
.Y(n_2606)
);

BUFx8_ASAP7_75t_SL g2607 ( 
.A(n_2181),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2130),
.Y(n_2608)
);

AND2x6_ASAP7_75t_L g2609 ( 
.A(n_2247),
.B(n_132),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_SL g2610 ( 
.A(n_2047),
.B(n_133),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2124),
.B(n_133),
.Y(n_2611)
);

AND2x6_ASAP7_75t_L g2612 ( 
.A(n_2080),
.B(n_134),
.Y(n_2612)
);

INVx3_ASAP7_75t_L g2613 ( 
.A(n_2159),
.Y(n_2613)
);

BUFx8_ASAP7_75t_L g2614 ( 
.A(n_2305),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2125),
.B(n_134),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2184),
.Y(n_2616)
);

CKINVDCx16_ASAP7_75t_R g2617 ( 
.A(n_2249),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_1998),
.Y(n_2618)
);

AO21x2_ASAP7_75t_L g2619 ( 
.A1(n_2217),
.A2(n_135),
.B(n_136),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2315),
.Y(n_2620)
);

BUFx4f_ASAP7_75t_L g2621 ( 
.A(n_2135),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2213),
.B(n_802),
.Y(n_2622)
);

NOR2xp33_ASAP7_75t_SL g2623 ( 
.A(n_2169),
.B(n_135),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2125),
.B(n_137),
.Y(n_2624)
);

BUFx6f_ASAP7_75t_L g2625 ( 
.A(n_2302),
.Y(n_2625)
);

NAND2x1p5_ASAP7_75t_L g2626 ( 
.A(n_2327),
.B(n_139),
.Y(n_2626)
);

OR2x6_ASAP7_75t_L g2627 ( 
.A(n_2312),
.B(n_138),
.Y(n_2627)
);

OR2x2_ASAP7_75t_L g2628 ( 
.A(n_2303),
.B(n_139),
.Y(n_2628)
);

INVx4_ASAP7_75t_L g2629 ( 
.A(n_2302),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2185),
.Y(n_2630)
);

BUFx3_ASAP7_75t_L g2631 ( 
.A(n_2181),
.Y(n_2631)
);

INVx1_ASAP7_75t_SL g2632 ( 
.A(n_2218),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2285),
.Y(n_2633)
);

BUFx4f_ASAP7_75t_L g2634 ( 
.A(n_2135),
.Y(n_2634)
);

INVx6_ASAP7_75t_L g2635 ( 
.A(n_2196),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2333),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2128),
.B(n_2143),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2291),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2292),
.Y(n_2639)
);

BUFx3_ASAP7_75t_L g2640 ( 
.A(n_2107),
.Y(n_2640)
);

INVx3_ASAP7_75t_L g2641 ( 
.A(n_2104),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2301),
.Y(n_2642)
);

HB1xp67_ASAP7_75t_L g2643 ( 
.A(n_2047),
.Y(n_2643)
);

INVx4_ASAP7_75t_L g2644 ( 
.A(n_2104),
.Y(n_2644)
);

AND2x4_ASAP7_75t_L g2645 ( 
.A(n_2280),
.B(n_140),
.Y(n_2645)
);

NAND2x1_ASAP7_75t_SL g2646 ( 
.A(n_2276),
.B(n_140),
.Y(n_2646)
);

NOR2x1_ASAP7_75t_L g2647 ( 
.A(n_2287),
.B(n_141),
.Y(n_2647)
);

INVxp67_ASAP7_75t_L g2648 ( 
.A(n_2208),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2288),
.Y(n_2649)
);

CKINVDCx20_ASAP7_75t_R g2650 ( 
.A(n_2236),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2128),
.B(n_142),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2132),
.Y(n_2652)
);

BUFx12f_ASAP7_75t_L g2653 ( 
.A(n_2001),
.Y(n_2653)
);

NOR2xp33_ASAP7_75t_SL g2654 ( 
.A(n_2293),
.B(n_142),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2143),
.B(n_143),
.Y(n_2655)
);

NAND2x1p5_ASAP7_75t_L g2656 ( 
.A(n_2035),
.B(n_2137),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2213),
.B(n_143),
.Y(n_2657)
);

CKINVDCx20_ASAP7_75t_R g2658 ( 
.A(n_2260),
.Y(n_2658)
);

OR2x2_ASAP7_75t_L g2659 ( 
.A(n_2303),
.B(n_144),
.Y(n_2659)
);

BUFx6f_ASAP7_75t_SL g2660 ( 
.A(n_2001),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2167),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2306),
.Y(n_2662)
);

NAND2x1p5_ASAP7_75t_L g2663 ( 
.A(n_2224),
.B(n_2026),
.Y(n_2663)
);

INVx1_ASAP7_75t_SL g2664 ( 
.A(n_2183),
.Y(n_2664)
);

NOR2xp33_ASAP7_75t_L g2665 ( 
.A(n_2011),
.B(n_819),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2011),
.B(n_144),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2022),
.Y(n_2667)
);

INVx1_ASAP7_75t_SL g2668 ( 
.A(n_2317),
.Y(n_2668)
);

INVxp67_ASAP7_75t_L g2669 ( 
.A(n_2208),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2288),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2261),
.B(n_146),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2264),
.Y(n_2672)
);

NOR2xp33_ASAP7_75t_SL g2673 ( 
.A(n_2299),
.B(n_147),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2317),
.Y(n_2674)
);

INVxp67_ASAP7_75t_L g2675 ( 
.A(n_2319),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2013),
.B(n_148),
.Y(n_2676)
);

AND2x4_ASAP7_75t_L g2677 ( 
.A(n_2026),
.B(n_149),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2319),
.Y(n_2678)
);

OR2x2_ASAP7_75t_L g2679 ( 
.A(n_2043),
.B(n_150),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2013),
.B(n_151),
.Y(n_2680)
);

OR2x2_ASAP7_75t_L g2681 ( 
.A(n_2160),
.B(n_151),
.Y(n_2681)
);

NAND2x1_ASAP7_75t_SL g2682 ( 
.A(n_2281),
.B(n_152),
.Y(n_2682)
);

INVx3_ASAP7_75t_L g2683 ( 
.A(n_2056),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2072),
.Y(n_2684)
);

AND2x4_ASAP7_75t_L g2685 ( 
.A(n_2041),
.B(n_2199),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2322),
.Y(n_2686)
);

INVx2_ASAP7_75t_SL g2687 ( 
.A(n_2107),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2019),
.B(n_152),
.Y(n_2688)
);

CKINVDCx20_ASAP7_75t_R g2689 ( 
.A(n_2307),
.Y(n_2689)
);

CKINVDCx20_ASAP7_75t_R g2690 ( 
.A(n_2282),
.Y(n_2690)
);

INVxp67_ASAP7_75t_SL g2691 ( 
.A(n_2322),
.Y(n_2691)
);

BUFx6f_ASAP7_75t_L g2692 ( 
.A(n_2262),
.Y(n_2692)
);

OR2x6_ASAP7_75t_L g2693 ( 
.A(n_2287),
.B(n_153),
.Y(n_2693)
);

BUFx6f_ASAP7_75t_L g2694 ( 
.A(n_2262),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2073),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2019),
.B(n_153),
.Y(n_2696)
);

BUFx3_ASAP7_75t_L g2697 ( 
.A(n_2115),
.Y(n_2697)
);

BUFx4f_ASAP7_75t_L g2698 ( 
.A(n_2041),
.Y(n_2698)
);

BUFx2_ASAP7_75t_L g2699 ( 
.A(n_2326),
.Y(n_2699)
);

BUFx4f_ASAP7_75t_L g2700 ( 
.A(n_2115),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2326),
.Y(n_2701)
);

AND2x4_ASAP7_75t_L g2702 ( 
.A(n_2156),
.B(n_154),
.Y(n_2702)
);

INVx3_ASAP7_75t_L g2703 ( 
.A(n_2283),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_2324),
.Y(n_2704)
);

INVx1_ASAP7_75t_SL g2705 ( 
.A(n_2156),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_SL g2706 ( 
.A(n_2330),
.B(n_154),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2036),
.B(n_2039),
.Y(n_2707)
);

NAND2x1p5_ASAP7_75t_L g2708 ( 
.A(n_2204),
.B(n_156),
.Y(n_2708)
);

NAND2x1p5_ASAP7_75t_L g2709 ( 
.A(n_2204),
.B(n_156),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2308),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2240),
.Y(n_2711)
);

AND2x6_ASAP7_75t_L g2712 ( 
.A(n_2080),
.B(n_155),
.Y(n_2712)
);

OR2x6_ASAP7_75t_L g2713 ( 
.A(n_2248),
.B(n_155),
.Y(n_2713)
);

INVx6_ASAP7_75t_L g2714 ( 
.A(n_2265),
.Y(n_2714)
);

NOR2x1_ASAP7_75t_L g2715 ( 
.A(n_2223),
.B(n_157),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2036),
.B(n_157),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2039),
.B(n_158),
.Y(n_2717)
);

CKINVDCx6p67_ASAP7_75t_R g2718 ( 
.A(n_2216),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2240),
.Y(n_2719)
);

BUFx3_ASAP7_75t_L g2720 ( 
.A(n_2256),
.Y(n_2720)
);

BUFx3_ASAP7_75t_L g2721 ( 
.A(n_2210),
.Y(n_2721)
);

INVx6_ASAP7_75t_L g2722 ( 
.A(n_2258),
.Y(n_2722)
);

BUFx4f_ASAP7_75t_L g2723 ( 
.A(n_2214),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2212),
.Y(n_2724)
);

OR2x2_ASAP7_75t_L g2725 ( 
.A(n_2160),
.B(n_159),
.Y(n_2725)
);

INVx4_ASAP7_75t_L g2726 ( 
.A(n_2262),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2245),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2158),
.B(n_810),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2222),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2161),
.B(n_159),
.Y(n_2730)
);

OR2x2_ASAP7_75t_L g2731 ( 
.A(n_2161),
.B(n_160),
.Y(n_2731)
);

OR2x2_ASAP7_75t_L g2732 ( 
.A(n_2162),
.B(n_161),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2253),
.B(n_161),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2245),
.Y(n_2734)
);

BUFx3_ASAP7_75t_L g2735 ( 
.A(n_2221),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2300),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2162),
.B(n_162),
.Y(n_2737)
);

BUFx2_ASAP7_75t_L g2738 ( 
.A(n_2248),
.Y(n_2738)
);

AND2x4_ASAP7_75t_L g2739 ( 
.A(n_2294),
.B(n_162),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2300),
.Y(n_2740)
);

INVx3_ASAP7_75t_L g2741 ( 
.A(n_2232),
.Y(n_2741)
);

NAND2x1p5_ASAP7_75t_L g2742 ( 
.A(n_2239),
.B(n_165),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2166),
.B(n_163),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2246),
.Y(n_2744)
);

NAND2x1p5_ASAP7_75t_L g2745 ( 
.A(n_2267),
.B(n_2268),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2166),
.B(n_163),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2100),
.Y(n_2747)
);

OR2x6_ASAP7_75t_L g2748 ( 
.A(n_2216),
.B(n_2229),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2100),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2171),
.B(n_165),
.Y(n_2750)
);

INVx4_ASAP7_75t_L g2751 ( 
.A(n_2272),
.Y(n_2751)
);

BUFx12f_ASAP7_75t_L g2752 ( 
.A(n_2294),
.Y(n_2752)
);

OR2x2_ASAP7_75t_L g2753 ( 
.A(n_2171),
.B(n_166),
.Y(n_2753)
);

BUFx6f_ASAP7_75t_L g2754 ( 
.A(n_2044),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2146),
.Y(n_2755)
);

BUFx2_ASAP7_75t_L g2756 ( 
.A(n_2254),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2174),
.B(n_2176),
.Y(n_2757)
);

BUFx6f_ASAP7_75t_L g2758 ( 
.A(n_2254),
.Y(n_2758)
);

BUFx6f_ASAP7_75t_L g2759 ( 
.A(n_2215),
.Y(n_2759)
);

BUFx2_ASAP7_75t_L g2760 ( 
.A(n_2174),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2176),
.B(n_166),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2180),
.B(n_2266),
.Y(n_2762)
);

CKINVDCx5p33_ASAP7_75t_R g2763 ( 
.A(n_2215),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2296),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2298),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_2269),
.B(n_167),
.Y(n_2766)
);

INVx3_ASAP7_75t_L g2767 ( 
.A(n_2229),
.Y(n_2767)
);

BUFx6f_ASAP7_75t_L g2768 ( 
.A(n_2231),
.Y(n_2768)
);

AND2x4_ASAP7_75t_L g2769 ( 
.A(n_2101),
.B(n_167),
.Y(n_2769)
);

OR2x6_ASAP7_75t_L g2770 ( 
.A(n_2231),
.B(n_168),
.Y(n_2770)
);

AND2x4_ASAP7_75t_L g2771 ( 
.A(n_2101),
.B(n_2103),
.Y(n_2771)
);

INVx2_ASAP7_75t_SL g2772 ( 
.A(n_2271),
.Y(n_2772)
);

INVx3_ASAP7_75t_L g2773 ( 
.A(n_2223),
.Y(n_2773)
);

NAND2x1_ASAP7_75t_L g2774 ( 
.A(n_2234),
.B(n_2103),
.Y(n_2774)
);

AND2x4_ASAP7_75t_L g2775 ( 
.A(n_1997),
.B(n_168),
.Y(n_2775)
);

BUFx8_ASAP7_75t_L g2776 ( 
.A(n_2102),
.Y(n_2776)
);

AND2x4_ASAP7_75t_L g2777 ( 
.A(n_1997),
.B(n_169),
.Y(n_2777)
);

INVx3_ASAP7_75t_L g2778 ( 
.A(n_2271),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2180),
.B(n_169),
.Y(n_2779)
);

AND2x4_ASAP7_75t_L g2780 ( 
.A(n_2002),
.B(n_170),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2149),
.Y(n_2781)
);

AND2x4_ASAP7_75t_L g2782 ( 
.A(n_2002),
.B(n_170),
.Y(n_2782)
);

BUFx12f_ASAP7_75t_L g2783 ( 
.A(n_2273),
.Y(n_2783)
);

OR2x2_ASAP7_75t_SL g2784 ( 
.A(n_2273),
.B(n_171),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2179),
.B(n_172),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2179),
.B(n_173),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_SL g2787 ( 
.A(n_2275),
.B(n_173),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2191),
.B(n_174),
.Y(n_2788)
);

NOR2x1_ASAP7_75t_SL g2789 ( 
.A(n_2149),
.B(n_174),
.Y(n_2789)
);

AND2x6_ASAP7_75t_L g2790 ( 
.A(n_2277),
.B(n_175),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2277),
.Y(n_2791)
);

AND2x4_ASAP7_75t_L g2792 ( 
.A(n_2234),
.B(n_175),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2191),
.B(n_176),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2151),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2151),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2020),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2122),
.B(n_178),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2122),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2152),
.Y(n_2799)
);

NOR2xp33_ASAP7_75t_L g2800 ( 
.A(n_2152),
.B(n_820),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2020),
.Y(n_2801)
);

CKINVDCx5p33_ASAP7_75t_R g2802 ( 
.A(n_2098),
.Y(n_2802)
);

AND2x4_ASAP7_75t_L g2803 ( 
.A(n_2098),
.B(n_178),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2187),
.Y(n_2804)
);

AND2x4_ASAP7_75t_L g2805 ( 
.A(n_2187),
.B(n_179),
.Y(n_2805)
);

OR2x2_ASAP7_75t_L g2806 ( 
.A(n_2259),
.B(n_181),
.Y(n_2806)
);

INVx1_ASAP7_75t_SL g2807 ( 
.A(n_2010),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2187),
.B(n_181),
.Y(n_2808)
);

NOR2xp33_ASAP7_75t_SL g2809 ( 
.A(n_2051),
.B(n_182),
.Y(n_2809)
);

INVx8_ASAP7_75t_L g2810 ( 
.A(n_2150),
.Y(n_2810)
);

AND2x4_ASAP7_75t_L g2811 ( 
.A(n_2187),
.B(n_184),
.Y(n_2811)
);

BUFx6f_ASAP7_75t_L g2812 ( 
.A(n_2017),
.Y(n_2812)
);

NOR2xp33_ASAP7_75t_SL g2813 ( 
.A(n_2051),
.B(n_185),
.Y(n_2813)
);

AND2x2_ASAP7_75t_SL g2814 ( 
.A(n_2074),
.B(n_185),
.Y(n_2814)
);

BUFx8_ASAP7_75t_SL g2815 ( 
.A(n_2111),
.Y(n_2815)
);

BUFx12f_ASAP7_75t_L g2816 ( 
.A(n_2111),
.Y(n_2816)
);

CKINVDCx20_ASAP7_75t_R g2817 ( 
.A(n_2007),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2187),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2225),
.B(n_801),
.Y(n_2819)
);

AO21x2_ASAP7_75t_L g2820 ( 
.A1(n_2217),
.A2(n_186),
.B(n_187),
.Y(n_2820)
);

NOR2x1p5_ASAP7_75t_SL g2821 ( 
.A(n_2296),
.B(n_186),
.Y(n_2821)
);

AND2x4_ASAP7_75t_L g2822 ( 
.A(n_2187),
.B(n_187),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_L g2823 ( 
.A(n_2017),
.Y(n_2823)
);

OR2x2_ASAP7_75t_L g2824 ( 
.A(n_2259),
.B(n_188),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2187),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2193),
.Y(n_2826)
);

AO21x2_ASAP7_75t_L g2827 ( 
.A1(n_2217),
.A2(n_188),
.B(n_189),
.Y(n_2827)
);

OR2x2_ASAP7_75t_L g2828 ( 
.A(n_2259),
.B(n_190),
.Y(n_2828)
);

AND2x4_ASAP7_75t_L g2829 ( 
.A(n_2187),
.B(n_190),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2145),
.B(n_191),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2145),
.B(n_191),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2187),
.B(n_192),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_SL g2833 ( 
.A(n_2123),
.B(n_192),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2187),
.Y(n_2834)
);

BUFx2_ASAP7_75t_L g2835 ( 
.A(n_2108),
.Y(n_2835)
);

NOR2xp33_ASAP7_75t_L g2836 ( 
.A(n_2225),
.B(n_808),
.Y(n_2836)
);

CKINVDCx8_ASAP7_75t_R g2837 ( 
.A(n_2111),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2804),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2818),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2825),
.Y(n_2840)
);

CKINVDCx5p33_ASAP7_75t_R g2841 ( 
.A(n_2400),
.Y(n_2841)
);

INVxp67_ASAP7_75t_SL g2842 ( 
.A(n_2335),
.Y(n_2842)
);

BUFx8_ASAP7_75t_SL g2843 ( 
.A(n_2815),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2336),
.B(n_193),
.Y(n_2844)
);

INVx5_ASAP7_75t_SL g2845 ( 
.A(n_2384),
.Y(n_2845)
);

BUFx3_ASAP7_75t_L g2846 ( 
.A(n_2817),
.Y(n_2846)
);

INVx3_ASAP7_75t_L g2847 ( 
.A(n_2621),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2834),
.B(n_193),
.Y(n_2848)
);

INVx3_ASAP7_75t_L g2849 ( 
.A(n_2621),
.Y(n_2849)
);

BUFx2_ASAP7_75t_L g2850 ( 
.A(n_2634),
.Y(n_2850)
);

BUFx12f_ASAP7_75t_L g2851 ( 
.A(n_2373),
.Y(n_2851)
);

INVxp67_ASAP7_75t_SL g2852 ( 
.A(n_2382),
.Y(n_2852)
);

OR2x2_ASAP7_75t_L g2853 ( 
.A(n_2412),
.B(n_2664),
.Y(n_2853)
);

INVx3_ASAP7_75t_L g2854 ( 
.A(n_2634),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2760),
.B(n_194),
.Y(n_2855)
);

BUFx4f_ASAP7_75t_L g2856 ( 
.A(n_2810),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2339),
.B(n_2570),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2352),
.Y(n_2858)
);

BUFx6f_ASAP7_75t_L g2859 ( 
.A(n_2343),
.Y(n_2859)
);

INVx1_ASAP7_75t_SL g2860 ( 
.A(n_2372),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2637),
.B(n_2350),
.Y(n_2861)
);

BUFx3_ASAP7_75t_L g2862 ( 
.A(n_2354),
.Y(n_2862)
);

INVx4_ASAP7_75t_L g2863 ( 
.A(n_2810),
.Y(n_2863)
);

BUFx2_ASAP7_75t_SL g2864 ( 
.A(n_2494),
.Y(n_2864)
);

INVx5_ASAP7_75t_L g2865 ( 
.A(n_2398),
.Y(n_2865)
);

INVx1_ASAP7_75t_SL g2866 ( 
.A(n_2835),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2710),
.Y(n_2867)
);

BUFx3_ASAP7_75t_L g2868 ( 
.A(n_2373),
.Y(n_2868)
);

CKINVDCx5p33_ASAP7_75t_R g2869 ( 
.A(n_2816),
.Y(n_2869)
);

BUFx3_ASAP7_75t_L g2870 ( 
.A(n_2367),
.Y(n_2870)
);

INVx3_ASAP7_75t_L g2871 ( 
.A(n_2644),
.Y(n_2871)
);

BUFx6f_ASAP7_75t_L g2872 ( 
.A(n_2343),
.Y(n_2872)
);

CKINVDCx11_ASAP7_75t_R g2873 ( 
.A(n_2837),
.Y(n_2873)
);

OR2x6_ASAP7_75t_L g2874 ( 
.A(n_2353),
.B(n_195),
.Y(n_2874)
);

INVx1_ASAP7_75t_SL g2875 ( 
.A(n_2416),
.Y(n_2875)
);

INVx3_ASAP7_75t_SL g2876 ( 
.A(n_2456),
.Y(n_2876)
);

BUFx2_ASAP7_75t_L g2877 ( 
.A(n_2382),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2516),
.Y(n_2878)
);

OR2x2_ASAP7_75t_L g2879 ( 
.A(n_2705),
.B(n_195),
.Y(n_2879)
);

BUFx6f_ASAP7_75t_L g2880 ( 
.A(n_2343),
.Y(n_2880)
);

AOI22xp33_ASAP7_75t_L g2881 ( 
.A1(n_2401),
.A2(n_199),
.B1(n_196),
.B2(n_197),
.Y(n_2881)
);

INVx3_ASAP7_75t_L g2882 ( 
.A(n_2644),
.Y(n_2882)
);

NAND2x1p5_ASAP7_75t_L g2883 ( 
.A(n_2509),
.B(n_196),
.Y(n_2883)
);

BUFx2_ASAP7_75t_L g2884 ( 
.A(n_2653),
.Y(n_2884)
);

INVx4_ASAP7_75t_L g2885 ( 
.A(n_2337),
.Y(n_2885)
);

BUFx12f_ASAP7_75t_L g2886 ( 
.A(n_2353),
.Y(n_2886)
);

BUFx2_ASAP7_75t_L g2887 ( 
.A(n_2397),
.Y(n_2887)
);

INVx5_ASAP7_75t_L g2888 ( 
.A(n_2398),
.Y(n_2888)
);

AND2x2_ASAP7_75t_SL g2889 ( 
.A(n_2407),
.B(n_197),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2516),
.Y(n_2890)
);

BUFx3_ASAP7_75t_L g2891 ( 
.A(n_2395),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2536),
.B(n_199),
.Y(n_2892)
);

AOI22xp33_ASAP7_75t_L g2893 ( 
.A1(n_2401),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_2893)
);

AND2x4_ASAP7_75t_L g2894 ( 
.A(n_2794),
.B(n_202),
.Y(n_2894)
);

BUFx2_ASAP7_75t_L g2895 ( 
.A(n_2700),
.Y(n_2895)
);

BUFx2_ASAP7_75t_L g2896 ( 
.A(n_2700),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2578),
.Y(n_2897)
);

BUFx3_ASAP7_75t_L g2898 ( 
.A(n_2559),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2525),
.Y(n_2899)
);

BUFx6f_ASAP7_75t_SL g2900 ( 
.A(n_2447),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2342),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2544),
.B(n_203),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2525),
.Y(n_2903)
);

INVx3_ASAP7_75t_SL g2904 ( 
.A(n_2499),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2356),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2771),
.B(n_205),
.Y(n_2906)
);

INVx1_ASAP7_75t_SL g2907 ( 
.A(n_2451),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2531),
.Y(n_2908)
);

INVx3_ASAP7_75t_L g2909 ( 
.A(n_2578),
.Y(n_2909)
);

BUFx12f_ASAP7_75t_L g2910 ( 
.A(n_2502),
.Y(n_2910)
);

BUFx2_ASAP7_75t_L g2911 ( 
.A(n_2698),
.Y(n_2911)
);

CKINVDCx20_ASAP7_75t_R g2912 ( 
.A(n_2408),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2357),
.Y(n_2913)
);

BUFx3_ASAP7_75t_L g2914 ( 
.A(n_2509),
.Y(n_2914)
);

AOI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_2802),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_2915)
);

INVx3_ASAP7_75t_L g2916 ( 
.A(n_2578),
.Y(n_2916)
);

BUFx12f_ASAP7_75t_L g2917 ( 
.A(n_2447),
.Y(n_2917)
);

BUFx6f_ASAP7_75t_L g2918 ( 
.A(n_2358),
.Y(n_2918)
);

BUFx6f_ASAP7_75t_L g2919 ( 
.A(n_2358),
.Y(n_2919)
);

INVx2_ASAP7_75t_SL g2920 ( 
.A(n_2337),
.Y(n_2920)
);

INVx1_ASAP7_75t_SL g2921 ( 
.A(n_2807),
.Y(n_2921)
);

INVx1_ASAP7_75t_SL g2922 ( 
.A(n_2344),
.Y(n_2922)
);

BUFx6f_ASAP7_75t_L g2923 ( 
.A(n_2358),
.Y(n_2923)
);

BUFx6f_ASAP7_75t_L g2924 ( 
.A(n_2359),
.Y(n_2924)
);

INVx3_ASAP7_75t_L g2925 ( 
.A(n_2337),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2357),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2771),
.B(n_206),
.Y(n_2927)
);

AOI22xp33_ASAP7_75t_SL g2928 ( 
.A1(n_2463),
.A2(n_2402),
.B1(n_2814),
.B2(n_2374),
.Y(n_2928)
);

NAND2x1p5_ASAP7_75t_L g2929 ( 
.A(n_2698),
.B(n_208),
.Y(n_2929)
);

CKINVDCx5p33_ASAP7_75t_R g2930 ( 
.A(n_2520),
.Y(n_2930)
);

CKINVDCx5p33_ASAP7_75t_R g2931 ( 
.A(n_2607),
.Y(n_2931)
);

INVx3_ASAP7_75t_L g2932 ( 
.A(n_2340),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2429),
.B(n_2795),
.Y(n_2933)
);

CKINVDCx5p33_ASAP7_75t_R g2934 ( 
.A(n_2590),
.Y(n_2934)
);

BUFx6f_ASAP7_75t_L g2935 ( 
.A(n_2359),
.Y(n_2935)
);

BUFx2_ASAP7_75t_SL g2936 ( 
.A(n_2424),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2365),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2365),
.Y(n_2938)
);

AOI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2505),
.A2(n_213),
.B1(n_208),
.B2(n_212),
.Y(n_2939)
);

INVxp67_ASAP7_75t_SL g2940 ( 
.A(n_2805),
.Y(n_2940)
);

INVx2_ASAP7_75t_SL g2941 ( 
.A(n_2576),
.Y(n_2941)
);

CKINVDCx11_ASAP7_75t_R g2942 ( 
.A(n_2650),
.Y(n_2942)
);

INVx5_ASAP7_75t_L g2943 ( 
.A(n_2398),
.Y(n_2943)
);

BUFx2_ASAP7_75t_SL g2944 ( 
.A(n_2424),
.Y(n_2944)
);

OR2x6_ASAP7_75t_L g2945 ( 
.A(n_2361),
.B(n_214),
.Y(n_2945)
);

CKINVDCx20_ASAP7_75t_R g2946 ( 
.A(n_2617),
.Y(n_2946)
);

CKINVDCx6p67_ASAP7_75t_R g2947 ( 
.A(n_2660),
.Y(n_2947)
);

INVx1_ASAP7_75t_SL g2948 ( 
.A(n_2344),
.Y(n_2948)
);

INVx8_ASAP7_75t_L g2949 ( 
.A(n_2499),
.Y(n_2949)
);

INVx1_ASAP7_75t_SL g2950 ( 
.A(n_2554),
.Y(n_2950)
);

BUFx2_ASAP7_75t_SL g2951 ( 
.A(n_2424),
.Y(n_2951)
);

INVx2_ASAP7_75t_SL g2952 ( 
.A(n_2576),
.Y(n_2952)
);

BUFx6f_ASAP7_75t_L g2953 ( 
.A(n_2359),
.Y(n_2953)
);

INVx2_ASAP7_75t_SL g2954 ( 
.A(n_2387),
.Y(n_2954)
);

BUFx12f_ASAP7_75t_L g2955 ( 
.A(n_2362),
.Y(n_2955)
);

AOI22xp33_ASAP7_75t_L g2956 ( 
.A1(n_2458),
.A2(n_217),
.B1(n_214),
.B2(n_215),
.Y(n_2956)
);

BUFx6f_ASAP7_75t_L g2957 ( 
.A(n_2394),
.Y(n_2957)
);

BUFx3_ASAP7_75t_L g2958 ( 
.A(n_2387),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2369),
.Y(n_2959)
);

INVx3_ASAP7_75t_L g2960 ( 
.A(n_2340),
.Y(n_2960)
);

INVx2_ASAP7_75t_SL g2961 ( 
.A(n_2635),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2369),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2444),
.Y(n_2963)
);

INVx4_ASAP7_75t_L g2964 ( 
.A(n_2398),
.Y(n_2964)
);

CKINVDCx14_ASAP7_75t_R g2965 ( 
.A(n_2597),
.Y(n_2965)
);

BUFx4_ASAP7_75t_SL g2966 ( 
.A(n_2549),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2444),
.Y(n_2967)
);

BUFx2_ASAP7_75t_L g2968 ( 
.A(n_2601),
.Y(n_2968)
);

BUFx2_ASAP7_75t_SL g2969 ( 
.A(n_2476),
.Y(n_2969)
);

AOI22xp33_ASAP7_75t_L g2970 ( 
.A1(n_2458),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_2970)
);

AOI22xp33_ASAP7_75t_SL g2971 ( 
.A1(n_2458),
.A2(n_221),
.B1(n_218),
.B2(n_220),
.Y(n_2971)
);

NAND2x1p5_ASAP7_75t_L g2972 ( 
.A(n_2407),
.B(n_220),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2445),
.Y(n_2973)
);

BUFx2_ASAP7_75t_SL g2974 ( 
.A(n_2476),
.Y(n_2974)
);

CKINVDCx20_ASAP7_75t_R g2975 ( 
.A(n_2776),
.Y(n_2975)
);

BUFx4_ASAP7_75t_SL g2976 ( 
.A(n_2549),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2445),
.Y(n_2977)
);

BUFx6f_ASAP7_75t_L g2978 ( 
.A(n_2394),
.Y(n_2978)
);

BUFx6f_ASAP7_75t_L g2979 ( 
.A(n_2394),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2452),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2452),
.Y(n_2981)
);

BUFx6f_ASAP7_75t_L g2982 ( 
.A(n_2411),
.Y(n_2982)
);

INVx3_ASAP7_75t_L g2983 ( 
.A(n_2351),
.Y(n_2983)
);

BUFx2_ASAP7_75t_R g2984 ( 
.A(n_2704),
.Y(n_2984)
);

INVx1_ASAP7_75t_SL g2985 ( 
.A(n_2554),
.Y(n_2985)
);

AND2x2_ASAP7_75t_L g2986 ( 
.A(n_2541),
.B(n_221),
.Y(n_2986)
);

INVx1_ASAP7_75t_SL g2987 ( 
.A(n_2470),
.Y(n_2987)
);

BUFx3_ASAP7_75t_L g2988 ( 
.A(n_2477),
.Y(n_2988)
);

BUFx2_ASAP7_75t_SL g2989 ( 
.A(n_2476),
.Y(n_2989)
);

BUFx4_ASAP7_75t_SL g2990 ( 
.A(n_2556),
.Y(n_2990)
);

BUFx8_ASAP7_75t_L g2991 ( 
.A(n_2660),
.Y(n_2991)
);

BUFx12f_ASAP7_75t_L g2992 ( 
.A(n_2510),
.Y(n_2992)
);

BUFx12f_ASAP7_75t_L g2993 ( 
.A(n_2515),
.Y(n_2993)
);

INVx3_ASAP7_75t_L g2994 ( 
.A(n_2351),
.Y(n_2994)
);

BUFx3_ASAP7_75t_L g2995 ( 
.A(n_2497),
.Y(n_2995)
);

BUFx3_ASAP7_75t_L g2996 ( 
.A(n_2537),
.Y(n_2996)
);

INVx3_ASAP7_75t_SL g2997 ( 
.A(n_2388),
.Y(n_2997)
);

BUFx10_ASAP7_75t_L g2998 ( 
.A(n_2348),
.Y(n_2998)
);

INVx5_ASAP7_75t_L g2999 ( 
.A(n_2558),
.Y(n_2999)
);

INVx5_ASAP7_75t_L g3000 ( 
.A(n_2558),
.Y(n_3000)
);

BUFx4f_ASAP7_75t_L g3001 ( 
.A(n_2478),
.Y(n_3001)
);

CKINVDCx5p33_ASAP7_75t_R g3002 ( 
.A(n_2752),
.Y(n_3002)
);

NAND2x1p5_ASAP7_75t_L g3003 ( 
.A(n_2426),
.B(n_222),
.Y(n_3003)
);

CKINVDCx5p33_ASAP7_75t_R g3004 ( 
.A(n_2776),
.Y(n_3004)
);

INVx1_ASAP7_75t_SL g3005 ( 
.A(n_2474),
.Y(n_3005)
);

AND2x4_ASAP7_75t_L g3006 ( 
.A(n_2641),
.B(n_223),
.Y(n_3006)
);

NAND2x1p5_ASAP7_75t_L g3007 ( 
.A(n_2426),
.B(n_223),
.Y(n_3007)
);

BUFx2_ASAP7_75t_L g3008 ( 
.A(n_2478),
.Y(n_3008)
);

BUFx2_ASAP7_75t_L g3009 ( 
.A(n_2478),
.Y(n_3009)
);

INVx5_ASAP7_75t_L g3010 ( 
.A(n_2558),
.Y(n_3010)
);

INVx3_ASAP7_75t_SL g3011 ( 
.A(n_2388),
.Y(n_3011)
);

INVx4_ASAP7_75t_L g3012 ( 
.A(n_2440),
.Y(n_3012)
);

INVx6_ASAP7_75t_SL g3013 ( 
.A(n_2556),
.Y(n_3013)
);

INVx5_ASAP7_75t_L g3014 ( 
.A(n_2558),
.Y(n_3014)
);

INVxp67_ASAP7_75t_SL g3015 ( 
.A(n_2805),
.Y(n_3015)
);

NAND2x1p5_ASAP7_75t_L g3016 ( 
.A(n_2440),
.B(n_224),
.Y(n_3016)
);

INVxp67_ASAP7_75t_L g3017 ( 
.A(n_2458),
.Y(n_3017)
);

BUFx6f_ASAP7_75t_L g3018 ( 
.A(n_2411),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2781),
.B(n_224),
.Y(n_3019)
);

INVx4_ASAP7_75t_L g3020 ( 
.A(n_2478),
.Y(n_3020)
);

INVxp67_ASAP7_75t_SL g3021 ( 
.A(n_2811),
.Y(n_3021)
);

INVx1_ASAP7_75t_SL g3022 ( 
.A(n_2522),
.Y(n_3022)
);

BUFx6f_ASAP7_75t_SL g3023 ( 
.A(n_2406),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2389),
.Y(n_3024)
);

BUFx6f_ASAP7_75t_L g3025 ( 
.A(n_2411),
.Y(n_3025)
);

BUFx10_ASAP7_75t_L g3026 ( 
.A(n_2348),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2393),
.Y(n_3027)
);

INVx1_ASAP7_75t_SL g3028 ( 
.A(n_2593),
.Y(n_3028)
);

NAND2x1p5_ASAP7_75t_L g3029 ( 
.A(n_2349),
.B(n_225),
.Y(n_3029)
);

INVx8_ASAP7_75t_L g3030 ( 
.A(n_2349),
.Y(n_3030)
);

BUFx12f_ASAP7_75t_L g3031 ( 
.A(n_2406),
.Y(n_3031)
);

CKINVDCx5p33_ASAP7_75t_R g3032 ( 
.A(n_2614),
.Y(n_3032)
);

HB1xp67_ASAP7_75t_L g3033 ( 
.A(n_2811),
.Y(n_3033)
);

BUFx2_ASAP7_75t_SL g3034 ( 
.A(n_2609),
.Y(n_3034)
);

BUFx3_ASAP7_75t_L g3035 ( 
.A(n_2546),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2545),
.Y(n_3036)
);

INVx6_ASAP7_75t_L g3037 ( 
.A(n_2614),
.Y(n_3037)
);

AND2x2_ASAP7_75t_L g3038 ( 
.A(n_2431),
.B(n_225),
.Y(n_3038)
);

BUFx6f_ASAP7_75t_L g3039 ( 
.A(n_2414),
.Y(n_3039)
);

AND2x4_ASAP7_75t_L g3040 ( 
.A(n_2641),
.B(n_226),
.Y(n_3040)
);

BUFx12f_ASAP7_75t_L g3041 ( 
.A(n_2415),
.Y(n_3041)
);

INVx5_ASAP7_75t_L g3042 ( 
.A(n_2609),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2781),
.B(n_226),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2633),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2396),
.Y(n_3045)
);

BUFx2_ASAP7_75t_L g3046 ( 
.A(n_2822),
.Y(n_3046)
);

CKINVDCx6p67_ASAP7_75t_R g3047 ( 
.A(n_2631),
.Y(n_3047)
);

BUFx6f_ASAP7_75t_L g3048 ( 
.A(n_2414),
.Y(n_3048)
);

INVxp67_ASAP7_75t_SL g3049 ( 
.A(n_2822),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2638),
.Y(n_3050)
);

BUFx3_ASAP7_75t_L g3051 ( 
.A(n_2640),
.Y(n_3051)
);

INVx8_ASAP7_75t_L g3052 ( 
.A(n_2609),
.Y(n_3052)
);

BUFx3_ASAP7_75t_L g3053 ( 
.A(n_2697),
.Y(n_3053)
);

CKINVDCx20_ASAP7_75t_R g3054 ( 
.A(n_2689),
.Y(n_3054)
);

BUFx2_ASAP7_75t_SL g3055 ( 
.A(n_2609),
.Y(n_3055)
);

INVxp67_ASAP7_75t_SL g3056 ( 
.A(n_2829),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2399),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2418),
.Y(n_3058)
);

BUFx12f_ASAP7_75t_L g3059 ( 
.A(n_2415),
.Y(n_3059)
);

BUFx3_ASAP7_75t_L g3060 ( 
.A(n_2410),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2433),
.Y(n_3061)
);

INVx2_ASAP7_75t_SL g3062 ( 
.A(n_2635),
.Y(n_3062)
);

INVx6_ASAP7_75t_SL g3063 ( 
.A(n_2702),
.Y(n_3063)
);

BUFx6f_ASAP7_75t_SL g3064 ( 
.A(n_2739),
.Y(n_3064)
);

BUFx6f_ASAP7_75t_L g3065 ( 
.A(n_2414),
.Y(n_3065)
);

INVx2_ASAP7_75t_SL g3066 ( 
.A(n_2567),
.Y(n_3066)
);

BUFx4f_ASAP7_75t_L g3067 ( 
.A(n_2708),
.Y(n_3067)
);

BUFx4_ASAP7_75t_SL g3068 ( 
.A(n_2720),
.Y(n_3068)
);

CKINVDCx11_ASAP7_75t_R g3069 ( 
.A(n_2658),
.Y(n_3069)
);

BUFx12f_ASAP7_75t_L g3070 ( 
.A(n_2709),
.Y(n_3070)
);

BUFx6f_ASAP7_75t_L g3071 ( 
.A(n_2446),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2707),
.B(n_228),
.Y(n_3072)
);

AND2x4_ASAP7_75t_L g3073 ( 
.A(n_2829),
.B(n_228),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2639),
.Y(n_3074)
);

BUFx2_ASAP7_75t_L g3075 ( 
.A(n_2783),
.Y(n_3075)
);

INVx1_ASAP7_75t_SL g3076 ( 
.A(n_2702),
.Y(n_3076)
);

BUFx2_ASAP7_75t_SL g3077 ( 
.A(n_2446),
.Y(n_3077)
);

BUFx6f_ASAP7_75t_L g3078 ( 
.A(n_2446),
.Y(n_3078)
);

BUFx3_ASAP7_75t_L g3079 ( 
.A(n_2410),
.Y(n_3079)
);

INVx6_ASAP7_75t_SL g3080 ( 
.A(n_2677),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2642),
.Y(n_3081)
);

INVx3_ASAP7_75t_SL g3082 ( 
.A(n_2529),
.Y(n_3082)
);

INVx2_ASAP7_75t_SL g3083 ( 
.A(n_2567),
.Y(n_3083)
);

INVx5_ASAP7_75t_L g3084 ( 
.A(n_2625),
.Y(n_3084)
);

HB1xp67_ASAP7_75t_L g3085 ( 
.A(n_2598),
.Y(n_3085)
);

INVx3_ASAP7_75t_L g3086 ( 
.A(n_2629),
.Y(n_3086)
);

BUFx3_ASAP7_75t_L g3087 ( 
.A(n_2589),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2826),
.Y(n_3088)
);

INVx2_ASAP7_75t_SL g3089 ( 
.A(n_2567),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2560),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2587),
.B(n_229),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2540),
.Y(n_3092)
);

INVx2_ASAP7_75t_L g3093 ( 
.A(n_2616),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2667),
.Y(n_3094)
);

BUFx3_ASAP7_75t_L g3095 ( 
.A(n_2605),
.Y(n_3095)
);

BUFx2_ASAP7_75t_SL g3096 ( 
.A(n_2449),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2630),
.Y(n_3097)
);

BUFx5_ASAP7_75t_L g3098 ( 
.A(n_2528),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2684),
.Y(n_3099)
);

INVx3_ASAP7_75t_SL g3100 ( 
.A(n_2529),
.Y(n_3100)
);

BUFx3_ASAP7_75t_L g3101 ( 
.A(n_2534),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2695),
.Y(n_3102)
);

CKINVDCx20_ASAP7_75t_R g3103 ( 
.A(n_2690),
.Y(n_3103)
);

INVx4_ASAP7_75t_L g3104 ( 
.A(n_2629),
.Y(n_3104)
);

BUFx3_ASAP7_75t_L g3105 ( 
.A(n_2534),
.Y(n_3105)
);

INVx8_ASAP7_75t_L g3106 ( 
.A(n_2677),
.Y(n_3106)
);

INVx3_ASAP7_75t_L g3107 ( 
.A(n_2751),
.Y(n_3107)
);

BUFx5_ASAP7_75t_L g3108 ( 
.A(n_2528),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2757),
.B(n_229),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2724),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2652),
.Y(n_3111)
);

AND2x4_ASAP7_75t_L g3112 ( 
.A(n_2498),
.B(n_230),
.Y(n_3112)
);

BUFx3_ASAP7_75t_L g3113 ( 
.A(n_2542),
.Y(n_3113)
);

INVx4_ASAP7_75t_L g3114 ( 
.A(n_2417),
.Y(n_3114)
);

BUFx3_ASAP7_75t_L g3115 ( 
.A(n_2542),
.Y(n_3115)
);

CKINVDCx5p33_ASAP7_75t_R g3116 ( 
.A(n_2585),
.Y(n_3116)
);

BUFx3_ASAP7_75t_L g3117 ( 
.A(n_2487),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2729),
.Y(n_3118)
);

INVx3_ASAP7_75t_L g3119 ( 
.A(n_2751),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2661),
.Y(n_3120)
);

CKINVDCx5p33_ASAP7_75t_R g3121 ( 
.A(n_2679),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2744),
.Y(n_3122)
);

INVx8_ASAP7_75t_L g3123 ( 
.A(n_2417),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2501),
.B(n_231),
.Y(n_3124)
);

BUFx6f_ASAP7_75t_L g3125 ( 
.A(n_2449),
.Y(n_3125)
);

BUFx2_ASAP7_75t_L g3126 ( 
.A(n_2364),
.Y(n_3126)
);

INVxp67_ASAP7_75t_SL g3127 ( 
.A(n_2519),
.Y(n_3127)
);

HB1xp67_ASAP7_75t_L g3128 ( 
.A(n_2599),
.Y(n_3128)
);

AND2x2_ASAP7_75t_L g3129 ( 
.A(n_2419),
.B(n_231),
.Y(n_3129)
);

INVx1_ASAP7_75t_SL g3130 ( 
.A(n_2550),
.Y(n_3130)
);

INVx2_ASAP7_75t_SL g3131 ( 
.A(n_2555),
.Y(n_3131)
);

BUFx6f_ASAP7_75t_L g3132 ( 
.A(n_2449),
.Y(n_3132)
);

NAND2x1p5_ASAP7_75t_L g3133 ( 
.A(n_2364),
.B(n_232),
.Y(n_3133)
);

INVx2_ASAP7_75t_SL g3134 ( 
.A(n_2555),
.Y(n_3134)
);

AND2x4_ASAP7_75t_L g3135 ( 
.A(n_2511),
.B(n_233),
.Y(n_3135)
);

CKINVDCx5p33_ASAP7_75t_R g3136 ( 
.A(n_2467),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2662),
.Y(n_3137)
);

BUFx6f_ASAP7_75t_L g3138 ( 
.A(n_2457),
.Y(n_3138)
);

INVx4_ASAP7_75t_L g3139 ( 
.A(n_2428),
.Y(n_3139)
);

AND2x4_ASAP7_75t_L g3140 ( 
.A(n_2685),
.B(n_235),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2747),
.Y(n_3141)
);

BUFx6f_ASAP7_75t_L g3142 ( 
.A(n_2457),
.Y(n_3142)
);

CKINVDCx14_ASAP7_75t_R g3143 ( 
.A(n_2471),
.Y(n_3143)
);

AND2x4_ASAP7_75t_L g3144 ( 
.A(n_2685),
.B(n_235),
.Y(n_3144)
);

INVx3_ASAP7_75t_L g3145 ( 
.A(n_2625),
.Y(n_3145)
);

BUFx6f_ASAP7_75t_L g3146 ( 
.A(n_2457),
.Y(n_3146)
);

INVx3_ASAP7_75t_L g3147 ( 
.A(n_2625),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2747),
.Y(n_3148)
);

BUFx3_ASAP7_75t_L g3149 ( 
.A(n_2568),
.Y(n_3149)
);

INVx2_ASAP7_75t_SL g3150 ( 
.A(n_2568),
.Y(n_3150)
);

INVx1_ASAP7_75t_SL g3151 ( 
.A(n_2557),
.Y(n_3151)
);

BUFx2_ASAP7_75t_L g3152 ( 
.A(n_2581),
.Y(n_3152)
);

NOR2xp33_ASAP7_75t_L g3153 ( 
.A(n_2420),
.B(n_236),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2749),
.Y(n_3154)
);

BUFx6f_ASAP7_75t_L g3155 ( 
.A(n_2517),
.Y(n_3155)
);

BUFx6f_ASAP7_75t_L g3156 ( 
.A(n_2517),
.Y(n_3156)
);

INVx3_ASAP7_75t_L g3157 ( 
.A(n_2423),
.Y(n_3157)
);

NAND2x1p5_ASAP7_75t_L g3158 ( 
.A(n_2581),
.B(n_236),
.Y(n_3158)
);

CKINVDCx8_ASAP7_75t_R g3159 ( 
.A(n_2612),
.Y(n_3159)
);

INVx3_ASAP7_75t_L g3160 ( 
.A(n_2423),
.Y(n_3160)
);

INVx2_ASAP7_75t_SL g3161 ( 
.A(n_2582),
.Y(n_3161)
);

BUFx8_ASAP7_75t_L g3162 ( 
.A(n_2739),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2749),
.Y(n_3163)
);

INVx5_ASAP7_75t_SL g3164 ( 
.A(n_2428),
.Y(n_3164)
);

INVx3_ASAP7_75t_L g3165 ( 
.A(n_2486),
.Y(n_3165)
);

BUFx6f_ASAP7_75t_L g3166 ( 
.A(n_2517),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2577),
.Y(n_3167)
);

BUFx3_ASAP7_75t_L g3168 ( 
.A(n_2582),
.Y(n_3168)
);

INVx5_ASAP7_75t_L g3169 ( 
.A(n_2526),
.Y(n_3169)
);

CKINVDCx5p33_ASAP7_75t_R g3170 ( 
.A(n_2506),
.Y(n_3170)
);

BUFx6f_ASAP7_75t_L g3171 ( 
.A(n_2526),
.Y(n_3171)
);

BUFx12f_ASAP7_75t_L g3172 ( 
.A(n_2346),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2632),
.B(n_237),
.Y(n_3173)
);

INVx4_ASAP7_75t_L g3174 ( 
.A(n_2434),
.Y(n_3174)
);

BUFx6f_ASAP7_75t_L g3175 ( 
.A(n_2526),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2378),
.B(n_237),
.Y(n_3176)
);

INVx4_ASAP7_75t_L g3177 ( 
.A(n_2434),
.Y(n_3177)
);

INVx8_ASAP7_75t_L g3178 ( 
.A(n_2450),
.Y(n_3178)
);

INVx2_ASAP7_75t_SL g3179 ( 
.A(n_2588),
.Y(n_3179)
);

BUFx24_ASAP7_75t_L g3180 ( 
.A(n_2450),
.Y(n_3180)
);

INVx1_ASAP7_75t_SL g3181 ( 
.A(n_2380),
.Y(n_3181)
);

BUFx6f_ASAP7_75t_L g3182 ( 
.A(n_2527),
.Y(n_3182)
);

BUFx2_ASAP7_75t_SL g3183 ( 
.A(n_2527),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2480),
.B(n_238),
.Y(n_3184)
);

INVx5_ASAP7_75t_L g3185 ( 
.A(n_2527),
.Y(n_3185)
);

BUFx3_ASAP7_75t_L g3186 ( 
.A(n_2588),
.Y(n_3186)
);

INVxp67_ASAP7_75t_SL g3187 ( 
.A(n_2519),
.Y(n_3187)
);

BUFx8_ASAP7_75t_L g3188 ( 
.A(n_2346),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2736),
.Y(n_3189)
);

BUFx2_ASAP7_75t_SL g3190 ( 
.A(n_2812),
.Y(n_3190)
);

INVx4_ASAP7_75t_L g3191 ( 
.A(n_2455),
.Y(n_3191)
);

BUFx4f_ASAP7_75t_SL g3192 ( 
.A(n_2721),
.Y(n_3192)
);

HB1xp67_ASAP7_75t_L g3193 ( 
.A(n_2643),
.Y(n_3193)
);

INVx3_ASAP7_75t_L g3194 ( 
.A(n_2486),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2740),
.Y(n_3195)
);

NAND2x1p5_ASAP7_75t_L g3196 ( 
.A(n_2592),
.B(n_239),
.Y(n_3196)
);

BUFx6f_ASAP7_75t_L g3197 ( 
.A(n_2812),
.Y(n_3197)
);

INVx1_ASAP7_75t_SL g3198 ( 
.A(n_2380),
.Y(n_3198)
);

INVx4_ASAP7_75t_L g3199 ( 
.A(n_2455),
.Y(n_3199)
);

AND2x4_ASAP7_75t_L g3200 ( 
.A(n_2772),
.B(n_239),
.Y(n_3200)
);

NOR2x1_ASAP7_75t_L g3201 ( 
.A(n_2547),
.B(n_2770),
.Y(n_3201)
);

INVx5_ASAP7_75t_L g3202 ( 
.A(n_2812),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2672),
.Y(n_3203)
);

INVx8_ASAP7_75t_L g3204 ( 
.A(n_2483),
.Y(n_3204)
);

BUFx3_ASAP7_75t_L g3205 ( 
.A(n_2592),
.Y(n_3205)
);

BUFx3_ASAP7_75t_L g3206 ( 
.A(n_2561),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2580),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_2583),
.Y(n_3208)
);

BUFx5_ASAP7_75t_L g3209 ( 
.A(n_2530),
.Y(n_3209)
);

CKINVDCx14_ASAP7_75t_R g3210 ( 
.A(n_2596),
.Y(n_3210)
);

BUFx2_ASAP7_75t_L g3211 ( 
.A(n_2602),
.Y(n_3211)
);

BUFx4f_ASAP7_75t_SL g3212 ( 
.A(n_2735),
.Y(n_3212)
);

INVx5_ASAP7_75t_L g3213 ( 
.A(n_2823),
.Y(n_3213)
);

NAND2x1p5_ASAP7_75t_L g3214 ( 
.A(n_2547),
.B(n_240),
.Y(n_3214)
);

BUFx6f_ASAP7_75t_L g3215 ( 
.A(n_2823),
.Y(n_3215)
);

BUFx2_ASAP7_75t_L g3216 ( 
.A(n_2803),
.Y(n_3216)
);

INVx8_ASAP7_75t_L g3217 ( 
.A(n_2483),
.Y(n_3217)
);

INVxp67_ASAP7_75t_L g3218 ( 
.A(n_2338),
.Y(n_3218)
);

BUFx12f_ASAP7_75t_L g3219 ( 
.A(n_2490),
.Y(n_3219)
);

BUFx3_ASAP7_75t_L g3220 ( 
.A(n_2484),
.Y(n_3220)
);

INVx2_ASAP7_75t_SL g3221 ( 
.A(n_2484),
.Y(n_3221)
);

INVx2_ASAP7_75t_SL g3222 ( 
.A(n_2485),
.Y(n_3222)
);

AOI22xp5_ASAP7_75t_L g3223 ( 
.A1(n_2496),
.A2(n_243),
.B1(n_240),
.B2(n_241),
.Y(n_3223)
);

NAND2x1p5_ASAP7_75t_L g3224 ( 
.A(n_2485),
.B(n_241),
.Y(n_3224)
);

NAND2x1_ASAP7_75t_L g3225 ( 
.A(n_2823),
.B(n_243),
.Y(n_3225)
);

INVx3_ASAP7_75t_L g3226 ( 
.A(n_2613),
.Y(n_3226)
);

INVx2_ASAP7_75t_SL g3227 ( 
.A(n_2539),
.Y(n_3227)
);

CKINVDCx8_ASAP7_75t_R g3228 ( 
.A(n_2612),
.Y(n_3228)
);

CKINVDCx5p33_ASAP7_75t_R g3229 ( 
.A(n_2718),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2504),
.B(n_244),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2600),
.Y(n_3231)
);

BUFx3_ASAP7_75t_L g3232 ( 
.A(n_2687),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2830),
.B(n_245),
.Y(n_3233)
);

BUFx4f_ASAP7_75t_SL g3234 ( 
.A(n_2464),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_2608),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_2831),
.B(n_245),
.Y(n_3236)
);

NAND2x1p5_ASAP7_75t_L g3237 ( 
.A(n_2508),
.B(n_246),
.Y(n_3237)
);

AND2x2_ASAP7_75t_L g3238 ( 
.A(n_2383),
.B(n_247),
.Y(n_3238)
);

BUFx5_ASAP7_75t_L g3239 ( 
.A(n_2530),
.Y(n_3239)
);

INVx2_ASAP7_75t_SL g3240 ( 
.A(n_2645),
.Y(n_3240)
);

INVx5_ASAP7_75t_L g3241 ( 
.A(n_2612),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2618),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2620),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2711),
.B(n_247),
.Y(n_3244)
);

BUFx3_ASAP7_75t_L g3245 ( 
.A(n_2645),
.Y(n_3245)
);

INVx2_ASAP7_75t_SL g3246 ( 
.A(n_2508),
.Y(n_3246)
);

INVx2_ASAP7_75t_SL g3247 ( 
.A(n_2723),
.Y(n_3247)
);

INVx4_ASAP7_75t_L g3248 ( 
.A(n_2612),
.Y(n_3248)
);

BUFx4f_ASAP7_75t_SL g3249 ( 
.A(n_2806),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_2636),
.Y(n_3250)
);

BUFx3_ASAP7_75t_L g3251 ( 
.A(n_2442),
.Y(n_3251)
);

BUFx12f_ASAP7_75t_L g3252 ( 
.A(n_2824),
.Y(n_3252)
);

BUFx4f_ASAP7_75t_L g3253 ( 
.A(n_2712),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2719),
.B(n_248),
.Y(n_3254)
);

AOI22xp33_ASAP7_75t_L g3255 ( 
.A1(n_2594),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_3255)
);

BUFx2_ASAP7_75t_L g3256 ( 
.A(n_2803),
.Y(n_3256)
);

INVx3_ASAP7_75t_L g3257 ( 
.A(n_2613),
.Y(n_3257)
);

BUFx2_ASAP7_75t_L g3258 ( 
.A(n_2775),
.Y(n_3258)
);

INVx5_ASAP7_75t_L g3259 ( 
.A(n_2712),
.Y(n_3259)
);

INVx3_ASAP7_75t_L g3260 ( 
.A(n_2726),
.Y(n_3260)
);

INVx3_ASAP7_75t_L g3261 ( 
.A(n_2726),
.Y(n_3261)
);

AND2x4_ASAP7_75t_L g3262 ( 
.A(n_2442),
.B(n_249),
.Y(n_3262)
);

CKINVDCx5p33_ASAP7_75t_R g3263 ( 
.A(n_2770),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2791),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2347),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_2462),
.Y(n_3266)
);

BUFx3_ASAP7_75t_L g3267 ( 
.A(n_2626),
.Y(n_3267)
);

INVx3_ASAP7_75t_L g3268 ( 
.A(n_2551),
.Y(n_3268)
);

BUFx6f_ASAP7_75t_L g3269 ( 
.A(n_2692),
.Y(n_3269)
);

NAND2x1p5_ASAP7_75t_L g3270 ( 
.A(n_2775),
.B(n_251),
.Y(n_3270)
);

AND2x4_ASAP7_75t_L g3271 ( 
.A(n_2727),
.B(n_252),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_2734),
.B(n_252),
.Y(n_3272)
);

INVx3_ASAP7_75t_L g3273 ( 
.A(n_2551),
.Y(n_3273)
);

INVx3_ASAP7_75t_SL g3274 ( 
.A(n_2828),
.Y(n_3274)
);

BUFx12f_ASAP7_75t_L g3275 ( 
.A(n_2742),
.Y(n_3275)
);

INVx1_ASAP7_75t_SL g3276 ( 
.A(n_2404),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_2838),
.Y(n_3277)
);

BUFx8_ASAP7_75t_L g3278 ( 
.A(n_2851),
.Y(n_3278)
);

BUFx3_ASAP7_75t_L g3279 ( 
.A(n_3075),
.Y(n_3279)
);

NAND2x1p5_ASAP7_75t_L g3280 ( 
.A(n_2856),
.B(n_2777),
.Y(n_3280)
);

CKINVDCx11_ASAP7_75t_R g3281 ( 
.A(n_2876),
.Y(n_3281)
);

CKINVDCx11_ASAP7_75t_R g3282 ( 
.A(n_2873),
.Y(n_3282)
);

AOI22xp33_ASAP7_75t_L g3283 ( 
.A1(n_2928),
.A2(n_2594),
.B1(n_2627),
.B2(n_3216),
.Y(n_3283)
);

HB1xp67_ASAP7_75t_L g3284 ( 
.A(n_2968),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3024),
.Y(n_3285)
);

AOI22xp33_ASAP7_75t_SL g3286 ( 
.A1(n_3064),
.A2(n_2813),
.B1(n_2809),
.B2(n_2623),
.Y(n_3286)
);

INVx5_ASAP7_75t_L g3287 ( 
.A(n_2874),
.Y(n_3287)
);

AOI22xp33_ASAP7_75t_L g3288 ( 
.A1(n_3256),
.A2(n_2627),
.B1(n_2693),
.B2(n_2334),
.Y(n_3288)
);

BUFx2_ASAP7_75t_L g3289 ( 
.A(n_2850),
.Y(n_3289)
);

BUFx12f_ASAP7_75t_L g3290 ( 
.A(n_2942),
.Y(n_3290)
);

AOI22xp33_ASAP7_75t_L g3291 ( 
.A1(n_3258),
.A2(n_2693),
.B1(n_2836),
.B2(n_2819),
.Y(n_3291)
);

AOI22xp33_ASAP7_75t_SL g3292 ( 
.A1(n_3064),
.A2(n_2673),
.B1(n_2591),
.B2(n_2789),
.Y(n_3292)
);

INVx2_ASAP7_75t_L g3293 ( 
.A(n_2839),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3024),
.Y(n_3294)
);

OAI22x1_ASAP7_75t_L g3295 ( 
.A1(n_3263),
.A2(n_2777),
.B1(n_2782),
.B2(n_2780),
.Y(n_3295)
);

NAND2x1p5_ASAP7_75t_L g3296 ( 
.A(n_2856),
.B(n_2863),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3027),
.Y(n_3297)
);

BUFx2_ASAP7_75t_SL g3298 ( 
.A(n_2900),
.Y(n_3298)
);

CKINVDCx16_ASAP7_75t_R g3299 ( 
.A(n_2975),
.Y(n_3299)
);

AOI22xp33_ASAP7_75t_SL g3300 ( 
.A1(n_3023),
.A2(n_2789),
.B1(n_2780),
.B2(n_2782),
.Y(n_3300)
);

AOI22xp5_ASAP7_75t_L g3301 ( 
.A1(n_3210),
.A2(n_2763),
.B1(n_2654),
.B2(n_2553),
.Y(n_3301)
);

CKINVDCx11_ASAP7_75t_R g3302 ( 
.A(n_2910),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_2861),
.B(n_2507),
.Y(n_3303)
);

CKINVDCx11_ASAP7_75t_R g3304 ( 
.A(n_2912),
.Y(n_3304)
);

BUFx8_ASAP7_75t_SL g3305 ( 
.A(n_2843),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3027),
.Y(n_3306)
);

BUFx8_ASAP7_75t_L g3307 ( 
.A(n_2900),
.Y(n_3307)
);

BUFx2_ASAP7_75t_L g3308 ( 
.A(n_3063),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3045),
.Y(n_3309)
);

AOI22xp33_ASAP7_75t_L g3310 ( 
.A1(n_3073),
.A2(n_2713),
.B1(n_2430),
.B2(n_2790),
.Y(n_3310)
);

INVx3_ASAP7_75t_L g3311 ( 
.A(n_3020),
.Y(n_3311)
);

AOI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_3001),
.A2(n_2691),
.B(n_2774),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3045),
.Y(n_3313)
);

AOI22xp33_ASAP7_75t_L g3314 ( 
.A1(n_3073),
.A2(n_2713),
.B1(n_2790),
.B2(n_2722),
.Y(n_3314)
);

AOI22xp33_ASAP7_75t_L g3315 ( 
.A1(n_3001),
.A2(n_2790),
.B1(n_2714),
.B2(n_2722),
.Y(n_3315)
);

AOI22xp33_ASAP7_75t_SL g3316 ( 
.A1(n_3023),
.A2(n_2712),
.B1(n_2391),
.B2(n_2422),
.Y(n_3316)
);

OAI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_3270),
.A2(n_2723),
.B1(n_2784),
.B2(n_2668),
.Y(n_3317)
);

OAI22xp5_ASAP7_75t_L g3318 ( 
.A1(n_3164),
.A2(n_2699),
.B1(n_2745),
.B2(n_2675),
.Y(n_3318)
);

AOI22xp33_ASAP7_75t_L g3319 ( 
.A1(n_2889),
.A2(n_2790),
.B1(n_2714),
.B2(n_2748),
.Y(n_3319)
);

OAI22xp5_ASAP7_75t_L g3320 ( 
.A1(n_3164),
.A2(n_2940),
.B1(n_3021),
.B2(n_3015),
.Y(n_3320)
);

INVx2_ASAP7_75t_SL g3321 ( 
.A(n_3068),
.Y(n_3321)
);

BUFx4f_ASAP7_75t_SL g3322 ( 
.A(n_2868),
.Y(n_3322)
);

INVx4_ASAP7_75t_L g3323 ( 
.A(n_3052),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3057),
.Y(n_3324)
);

AOI22xp33_ASAP7_75t_L g3325 ( 
.A1(n_3046),
.A2(n_2748),
.B1(n_2728),
.B2(n_2767),
.Y(n_3325)
);

INVxp67_ASAP7_75t_SL g3326 ( 
.A(n_3049),
.Y(n_3326)
);

CKINVDCx6p67_ASAP7_75t_R g3327 ( 
.A(n_2870),
.Y(n_3327)
);

CKINVDCx11_ASAP7_75t_R g3328 ( 
.A(n_2860),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_2867),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3264),
.Y(n_3330)
);

BUFx10_ASAP7_75t_L g3331 ( 
.A(n_3037),
.Y(n_3331)
);

BUFx2_ASAP7_75t_L g3332 ( 
.A(n_3063),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_2842),
.B(n_2538),
.Y(n_3333)
);

AOI22xp33_ASAP7_75t_L g3334 ( 
.A1(n_3162),
.A2(n_2767),
.B1(n_2778),
.B2(n_2800),
.Y(n_3334)
);

OAI22xp5_ASAP7_75t_L g3335 ( 
.A1(n_3056),
.A2(n_2648),
.B1(n_2669),
.B2(n_2756),
.Y(n_3335)
);

OAI22xp5_ASAP7_75t_L g3336 ( 
.A1(n_3020),
.A2(n_2762),
.B1(n_2769),
.B2(n_2738),
.Y(n_3336)
);

INVx1_ASAP7_75t_SL g3337 ( 
.A(n_3069),
.Y(n_3337)
);

CKINVDCx5p33_ASAP7_75t_R g3338 ( 
.A(n_2841),
.Y(n_3338)
);

AOI22xp33_ASAP7_75t_L g3339 ( 
.A1(n_3162),
.A2(n_3013),
.B1(n_3067),
.B2(n_3201),
.Y(n_3339)
);

BUFx2_ASAP7_75t_L g3340 ( 
.A(n_3080),
.Y(n_3340)
);

INVx6_ASAP7_75t_L g3341 ( 
.A(n_2991),
.Y(n_3341)
);

INVx6_ASAP7_75t_L g3342 ( 
.A(n_2991),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_2857),
.B(n_2606),
.Y(n_3343)
);

BUFx6f_ASAP7_75t_L g3344 ( 
.A(n_2859),
.Y(n_3344)
);

AOI22xp5_ASAP7_75t_SL g3345 ( 
.A1(n_3103),
.A2(n_2712),
.B1(n_2769),
.B2(n_2785),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_3167),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_3013),
.A2(n_2778),
.B1(n_2665),
.B2(n_2579),
.Y(n_3347)
);

BUFx3_ASAP7_75t_L g3348 ( 
.A(n_2862),
.Y(n_3348)
);

OAI22xp5_ASAP7_75t_L g3349 ( 
.A1(n_3253),
.A2(n_2681),
.B1(n_2731),
.B2(n_2725),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_3208),
.Y(n_3350)
);

OAI22xp5_ASAP7_75t_L g3351 ( 
.A1(n_3253),
.A2(n_3100),
.B1(n_3082),
.B2(n_3114),
.Y(n_3351)
);

BUFx12f_ASAP7_75t_L g3352 ( 
.A(n_2869),
.Y(n_3352)
);

OAI22xp33_ASAP7_75t_SL g3353 ( 
.A1(n_2874),
.A2(n_2533),
.B1(n_2492),
.B2(n_2787),
.Y(n_3353)
);

INVx6_ASAP7_75t_L g3354 ( 
.A(n_2863),
.Y(n_3354)
);

AND2x4_ASAP7_75t_L g3355 ( 
.A(n_2964),
.B(n_2674),
.Y(n_3355)
);

AOI22xp33_ASAP7_75t_L g3356 ( 
.A1(n_3067),
.A2(n_2603),
.B1(n_2686),
.B2(n_2678),
.Y(n_3356)
);

AOI22xp33_ASAP7_75t_L g3357 ( 
.A1(n_2917),
.A2(n_2701),
.B1(n_2706),
.B2(n_2671),
.Y(n_3357)
);

INVx6_ASAP7_75t_L g3358 ( 
.A(n_2885),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3057),
.Y(n_3359)
);

AOI22xp33_ASAP7_75t_L g3360 ( 
.A1(n_3271),
.A2(n_2443),
.B1(n_2453),
.B2(n_2657),
.Y(n_3360)
);

BUFx10_ASAP7_75t_L g3361 ( 
.A(n_3037),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3058),
.Y(n_3362)
);

OAI21xp5_ASAP7_75t_SL g3363 ( 
.A1(n_2883),
.A2(n_2647),
.B(n_2793),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_2933),
.B(n_2730),
.Y(n_3364)
);

CKINVDCx11_ASAP7_75t_R g3365 ( 
.A(n_2947),
.Y(n_3365)
);

INVx8_ASAP7_75t_L g3366 ( 
.A(n_2886),
.Y(n_3366)
);

OAI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_3114),
.A2(n_3174),
.B1(n_3177),
.B2(n_3139),
.Y(n_3367)
);

AOI22xp33_ASAP7_75t_L g3368 ( 
.A1(n_3271),
.A2(n_2657),
.B1(n_2375),
.B2(n_2768),
.Y(n_3368)
);

INVx6_ASAP7_75t_L g3369 ( 
.A(n_2885),
.Y(n_3369)
);

AND2x2_ASAP7_75t_L g3370 ( 
.A(n_3038),
.B(n_2564),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3058),
.Y(n_3371)
);

AOI22xp33_ASAP7_75t_SL g3372 ( 
.A1(n_3123),
.A2(n_2797),
.B1(n_2792),
.B2(n_2436),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3061),
.Y(n_3373)
);

CKINVDCx14_ASAP7_75t_R g3374 ( 
.A(n_2965),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_3235),
.Y(n_3375)
);

CKINVDCx11_ASAP7_75t_R g3376 ( 
.A(n_2946),
.Y(n_3376)
);

BUFx6f_ASAP7_75t_L g3377 ( 
.A(n_2859),
.Y(n_3377)
);

INVx2_ASAP7_75t_SL g3378 ( 
.A(n_2847),
.Y(n_3378)
);

INVx1_ASAP7_75t_SL g3379 ( 
.A(n_2875),
.Y(n_3379)
);

AOI22xp33_ASAP7_75t_L g3380 ( 
.A1(n_3188),
.A2(n_2768),
.B1(n_2448),
.B2(n_2468),
.Y(n_3380)
);

CKINVDCx11_ASAP7_75t_R g3381 ( 
.A(n_2846),
.Y(n_3381)
);

AOI22xp33_ASAP7_75t_L g3382 ( 
.A1(n_3188),
.A2(n_2768),
.B1(n_2489),
.B2(n_2441),
.Y(n_3382)
);

AOI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_3033),
.A2(n_2715),
.B1(n_2622),
.B2(n_2469),
.Y(n_3383)
);

INVx8_ASAP7_75t_L g3384 ( 
.A(n_3030),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3061),
.Y(n_3385)
);

CKINVDCx11_ASAP7_75t_R g3386 ( 
.A(n_2955),
.Y(n_3386)
);

BUFx10_ASAP7_75t_L g3387 ( 
.A(n_3004),
.Y(n_3387)
);

CKINVDCx5p33_ASAP7_75t_R g3388 ( 
.A(n_2966),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3203),
.Y(n_3389)
);

AOI22xp33_ASAP7_75t_SL g3390 ( 
.A1(n_3123),
.A2(n_2792),
.B1(n_2403),
.B2(n_2376),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_2878),
.Y(n_3391)
);

BUFx8_ASAP7_75t_SL g3392 ( 
.A(n_2934),
.Y(n_3392)
);

INVx4_ASAP7_75t_L g3393 ( 
.A(n_3052),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_2878),
.Y(n_3394)
);

AND2x2_ASAP7_75t_L g3395 ( 
.A(n_2892),
.B(n_2750),
.Y(n_3395)
);

CKINVDCx6p67_ASAP7_75t_R g3396 ( 
.A(n_3180),
.Y(n_3396)
);

BUFx2_ASAP7_75t_L g3397 ( 
.A(n_3080),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_2890),
.Y(n_3398)
);

AOI22xp33_ASAP7_75t_SL g3399 ( 
.A1(n_3178),
.A2(n_2663),
.B1(n_2569),
.B2(n_2796),
.Y(n_3399)
);

OAI22xp33_ASAP7_75t_L g3400 ( 
.A1(n_2945),
.A2(n_2753),
.B1(n_2732),
.B2(n_2628),
.Y(n_3400)
);

INVx4_ASAP7_75t_L g3401 ( 
.A(n_2865),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_2890),
.Y(n_3402)
);

AOI22xp33_ASAP7_75t_L g3403 ( 
.A1(n_3140),
.A2(n_2766),
.B1(n_2360),
.B2(n_2773),
.Y(n_3403)
);

BUFx6f_ASAP7_75t_L g3404 ( 
.A(n_2859),
.Y(n_3404)
);

AOI22xp33_ASAP7_75t_L g3405 ( 
.A1(n_3140),
.A2(n_2773),
.B1(n_2796),
.B2(n_2798),
.Y(n_3405)
);

AOI22xp33_ASAP7_75t_L g3406 ( 
.A1(n_3144),
.A2(n_2801),
.B1(n_2659),
.B2(n_2584),
.Y(n_3406)
);

INVx1_ASAP7_75t_SL g3407 ( 
.A(n_3192),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_2840),
.Y(n_3408)
);

INVx6_ASAP7_75t_L g3409 ( 
.A(n_2992),
.Y(n_3409)
);

OAI22xp5_ASAP7_75t_L g3410 ( 
.A1(n_3139),
.A2(n_3177),
.B1(n_3191),
.B2(n_3174),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_2899),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_2899),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_2840),
.B(n_2381),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_2903),
.Y(n_3414)
);

CKINVDCx5p33_ASAP7_75t_R g3415 ( 
.A(n_2976),
.Y(n_3415)
);

BUFx3_ASAP7_75t_L g3416 ( 
.A(n_2898),
.Y(n_3416)
);

BUFx10_ASAP7_75t_L g3417 ( 
.A(n_3032),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_2903),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_2858),
.B(n_2385),
.Y(n_3419)
);

INVx3_ASAP7_75t_L g3420 ( 
.A(n_2964),
.Y(n_3420)
);

OAI22xp33_ASAP7_75t_L g3421 ( 
.A1(n_2945),
.A2(n_2521),
.B1(n_2595),
.B2(n_2482),
.Y(n_3421)
);

INVx5_ASAP7_75t_L g3422 ( 
.A(n_2865),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3189),
.B(n_2377),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_2986),
.B(n_2355),
.Y(n_3424)
);

OAI22xp5_ASAP7_75t_L g3425 ( 
.A1(n_3191),
.A2(n_2832),
.B1(n_2808),
.B2(n_2788),
.Y(n_3425)
);

AOI22xp33_ASAP7_75t_SL g3426 ( 
.A1(n_3178),
.A2(n_3204),
.B1(n_3217),
.B2(n_3030),
.Y(n_3426)
);

AOI22xp33_ASAP7_75t_L g3427 ( 
.A1(n_3144),
.A2(n_2604),
.B1(n_2611),
.B2(n_2571),
.Y(n_3427)
);

AOI22xp33_ASAP7_75t_L g3428 ( 
.A1(n_3172),
.A2(n_2624),
.B1(n_2651),
.B2(n_2615),
.Y(n_3428)
);

AOI22xp33_ASAP7_75t_L g3429 ( 
.A1(n_3143),
.A2(n_2655),
.B1(n_2379),
.B2(n_2341),
.Y(n_3429)
);

OAI21xp5_ASAP7_75t_SL g3430 ( 
.A1(n_3029),
.A2(n_2656),
.B(n_2786),
.Y(n_3430)
);

AOI22xp33_ASAP7_75t_L g3431 ( 
.A1(n_3106),
.A2(n_2409),
.B1(n_2390),
.B2(n_2513),
.Y(n_3431)
);

OAI22xp5_ASAP7_75t_L g3432 ( 
.A1(n_3199),
.A2(n_2565),
.B1(n_2566),
.B2(n_2737),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_2913),
.Y(n_3433)
);

BUFx12f_ASAP7_75t_L g3434 ( 
.A(n_2931),
.Y(n_3434)
);

INVx3_ASAP7_75t_L g3435 ( 
.A(n_2871),
.Y(n_3435)
);

NAND2x1p5_ASAP7_75t_L g3436 ( 
.A(n_2847),
.B(n_2475),
.Y(n_3436)
);

AOI22xp33_ASAP7_75t_L g3437 ( 
.A1(n_3106),
.A2(n_2562),
.B1(n_2500),
.B2(n_2493),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_2913),
.Y(n_3438)
);

AOI22xp33_ASAP7_75t_L g3439 ( 
.A1(n_3031),
.A2(n_2666),
.B1(n_2680),
.B2(n_2676),
.Y(n_3439)
);

CKINVDCx6p67_ASAP7_75t_R g3440 ( 
.A(n_2904),
.Y(n_3440)
);

OAI21xp33_ASAP7_75t_L g3441 ( 
.A1(n_3255),
.A2(n_2821),
.B(n_2682),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_2938),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_L g3443 ( 
.A1(n_3041),
.A2(n_2688),
.B1(n_2716),
.B2(n_2696),
.Y(n_3443)
);

OAI21xp33_ASAP7_75t_SL g3444 ( 
.A1(n_3248),
.A2(n_2682),
.B(n_2646),
.Y(n_3444)
);

OAI22xp5_ASAP7_75t_L g3445 ( 
.A1(n_3199),
.A2(n_2743),
.B1(n_2746),
.B2(n_2345),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_2938),
.Y(n_3446)
);

AOI22xp5_ASAP7_75t_SL g3447 ( 
.A1(n_2990),
.A2(n_2386),
.B1(n_2473),
.B2(n_2472),
.Y(n_3447)
);

BUFx8_ASAP7_75t_L g3448 ( 
.A(n_2884),
.Y(n_3448)
);

BUFx6f_ASAP7_75t_L g3449 ( 
.A(n_2872),
.Y(n_3449)
);

AOI22xp33_ASAP7_75t_SL g3450 ( 
.A1(n_3204),
.A2(n_3217),
.B1(n_3059),
.B2(n_3009),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3276),
.B(n_2481),
.Y(n_3451)
);

AOI22xp33_ASAP7_75t_L g3452 ( 
.A1(n_3234),
.A2(n_2717),
.B1(n_2548),
.B2(n_2758),
.Y(n_3452)
);

AOI22xp33_ASAP7_75t_L g3453 ( 
.A1(n_3249),
.A2(n_2758),
.B1(n_2610),
.B2(n_2488),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_3074),
.Y(n_3454)
);

INVx6_ASAP7_75t_L g3455 ( 
.A(n_2993),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3189),
.B(n_2491),
.Y(n_3456)
);

OAI22xp5_ASAP7_75t_L g3457 ( 
.A1(n_2997),
.A2(n_2733),
.B1(n_2799),
.B2(n_2779),
.Y(n_3457)
);

CKINVDCx20_ASAP7_75t_R g3458 ( 
.A(n_3054),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_L g3459 ( 
.A(n_3011),
.B(n_2479),
.Y(n_3459)
);

AOI22xp33_ASAP7_75t_L g3460 ( 
.A1(n_3070),
.A2(n_2758),
.B1(n_2518),
.B2(n_2524),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_2926),
.Y(n_3461)
);

INVx6_ASAP7_75t_L g3462 ( 
.A(n_3219),
.Y(n_3462)
);

CKINVDCx11_ASAP7_75t_R g3463 ( 
.A(n_3047),
.Y(n_3463)
);

INVx8_ASAP7_75t_L g3464 ( 
.A(n_2949),
.Y(n_3464)
);

OAI22xp5_ASAP7_75t_L g3465 ( 
.A1(n_3224),
.A2(n_2761),
.B1(n_2366),
.B2(n_2370),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_2853),
.B(n_3085),
.Y(n_3466)
);

CKINVDCx11_ASAP7_75t_R g3467 ( 
.A(n_3275),
.Y(n_3467)
);

OAI22xp33_ASAP7_75t_L g3468 ( 
.A1(n_3214),
.A2(n_2543),
.B1(n_2514),
.B2(n_2425),
.Y(n_3468)
);

OAI22xp5_ASAP7_75t_L g3469 ( 
.A1(n_3133),
.A2(n_2512),
.B1(n_2432),
.B2(n_2435),
.Y(n_3469)
);

CKINVDCx5p33_ASAP7_75t_R g3470 ( 
.A(n_2930),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_2937),
.Y(n_3471)
);

BUFx6f_ASAP7_75t_L g3472 ( 
.A(n_2872),
.Y(n_3472)
);

AOI22xp33_ASAP7_75t_L g3473 ( 
.A1(n_3200),
.A2(n_2759),
.B1(n_2833),
.B2(n_2421),
.Y(n_3473)
);

BUFx4f_ASAP7_75t_L g3474 ( 
.A(n_2849),
.Y(n_3474)
);

BUFx4f_ASAP7_75t_SL g3475 ( 
.A(n_2914),
.Y(n_3475)
);

CKINVDCx11_ASAP7_75t_R g3476 ( 
.A(n_2949),
.Y(n_3476)
);

CKINVDCx11_ASAP7_75t_R g3477 ( 
.A(n_2998),
.Y(n_3477)
);

BUFx6f_ASAP7_75t_L g3478 ( 
.A(n_2872),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_2959),
.Y(n_3479)
);

INVx6_ASAP7_75t_L g3480 ( 
.A(n_2891),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_2962),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3074),
.Y(n_3482)
);

AO22x1_ASAP7_75t_L g3483 ( 
.A1(n_2865),
.A2(n_2646),
.B1(n_2437),
.B2(n_2439),
.Y(n_3483)
);

INVx3_ASAP7_75t_SL g3484 ( 
.A(n_3229),
.Y(n_3484)
);

CKINVDCx11_ASAP7_75t_R g3485 ( 
.A(n_2998),
.Y(n_3485)
);

INVx1_ASAP7_75t_SL g3486 ( 
.A(n_3212),
.Y(n_3486)
);

AOI22xp33_ASAP7_75t_L g3487 ( 
.A1(n_3200),
.A2(n_2759),
.B1(n_2413),
.B2(n_2459),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3081),
.Y(n_3488)
);

OAI22xp5_ASAP7_75t_L g3489 ( 
.A1(n_3158),
.A2(n_2454),
.B1(n_2460),
.B2(n_2774),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3081),
.Y(n_3490)
);

BUFx3_ASAP7_75t_L g3491 ( 
.A(n_2988),
.Y(n_3491)
);

BUFx12f_ASAP7_75t_L g3492 ( 
.A(n_3002),
.Y(n_3492)
);

BUFx2_ASAP7_75t_SL g3493 ( 
.A(n_2849),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_2963),
.Y(n_3494)
);

INVx3_ASAP7_75t_L g3495 ( 
.A(n_2871),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_2967),
.Y(n_3496)
);

OAI22xp5_ASAP7_75t_L g3497 ( 
.A1(n_3196),
.A2(n_2670),
.B1(n_2649),
.B2(n_2759),
.Y(n_3497)
);

CKINVDCx11_ASAP7_75t_R g3498 ( 
.A(n_3026),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_2973),
.Y(n_3499)
);

INVx1_ASAP7_75t_SL g3500 ( 
.A(n_2866),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3195),
.B(n_2764),
.Y(n_3501)
);

OAI22xp33_ASAP7_75t_L g3502 ( 
.A1(n_3237),
.A2(n_2649),
.B1(n_2670),
.B2(n_2683),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3128),
.B(n_2765),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3195),
.B(n_2683),
.Y(n_3504)
);

OAI22xp33_ASAP7_75t_L g3505 ( 
.A1(n_3170),
.A2(n_2741),
.B1(n_2703),
.B2(n_2755),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3088),
.Y(n_3506)
);

INVx3_ASAP7_75t_L g3507 ( 
.A(n_2882),
.Y(n_3507)
);

INVx5_ASAP7_75t_L g3508 ( 
.A(n_2888),
.Y(n_3508)
);

AOI22xp33_ASAP7_75t_L g3509 ( 
.A1(n_3252),
.A2(n_2619),
.B1(n_2820),
.B2(n_2371),
.Y(n_3509)
);

AOI22xp33_ASAP7_75t_L g3510 ( 
.A1(n_3126),
.A2(n_2827),
.B1(n_2755),
.B2(n_2741),
.Y(n_3510)
);

CKINVDCx20_ASAP7_75t_R g3511 ( 
.A(n_2845),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_2977),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3130),
.B(n_2703),
.Y(n_3513)
);

AOI22xp33_ASAP7_75t_L g3514 ( 
.A1(n_3008),
.A2(n_2392),
.B1(n_2535),
.B2(n_2532),
.Y(n_3514)
);

INVx1_ASAP7_75t_SL g3515 ( 
.A(n_3005),
.Y(n_3515)
);

OAI22xp5_ASAP7_75t_L g3516 ( 
.A1(n_3127),
.A2(n_2563),
.B1(n_2572),
.B2(n_2552),
.Y(n_3516)
);

BUFx3_ASAP7_75t_L g3517 ( 
.A(n_2995),
.Y(n_3517)
);

AOI22xp5_ASAP7_75t_L g3518 ( 
.A1(n_3121),
.A2(n_2535),
.B1(n_2552),
.B2(n_2532),
.Y(n_3518)
);

INVx6_ASAP7_75t_L g3519 ( 
.A(n_3026),
.Y(n_3519)
);

OAI22xp33_ASAP7_75t_L g3520 ( 
.A1(n_2929),
.A2(n_2573),
.B1(n_2563),
.B2(n_2572),
.Y(n_3520)
);

INVx1_ASAP7_75t_SL g3521 ( 
.A(n_3022),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3193),
.B(n_3129),
.Y(n_3522)
);

OAI22xp5_ASAP7_75t_L g3523 ( 
.A1(n_3187),
.A2(n_2586),
.B1(n_2573),
.B2(n_2461),
.Y(n_3523)
);

BUFx4f_ASAP7_75t_L g3524 ( 
.A(n_2854),
.Y(n_3524)
);

CKINVDCx20_ASAP7_75t_R g3525 ( 
.A(n_2845),
.Y(n_3525)
);

CKINVDCx11_ASAP7_75t_R g3526 ( 
.A(n_3159),
.Y(n_3526)
);

AOI22xp5_ASAP7_75t_L g3527 ( 
.A1(n_3136),
.A2(n_2586),
.B1(n_2368),
.B2(n_2405),
.Y(n_3527)
);

INVx6_ASAP7_75t_L g3528 ( 
.A(n_3104),
.Y(n_3528)
);

AOI22xp33_ASAP7_75t_L g3529 ( 
.A1(n_3220),
.A2(n_2427),
.B1(n_2438),
.B2(n_2363),
.Y(n_3529)
);

BUFx6f_ASAP7_75t_L g3530 ( 
.A(n_2880),
.Y(n_3530)
);

INVxp67_ASAP7_75t_SL g3531 ( 
.A(n_3149),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3151),
.B(n_2980),
.Y(n_3532)
);

OAI22x1_ASAP7_75t_L g3533 ( 
.A1(n_3248),
.A2(n_3116),
.B1(n_3218),
.B2(n_3241),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_2981),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3092),
.Y(n_3535)
);

CKINVDCx20_ASAP7_75t_R g3536 ( 
.A(n_2877),
.Y(n_3536)
);

INVx1_ASAP7_75t_SL g3537 ( 
.A(n_3028),
.Y(n_3537)
);

BUFx12f_ASAP7_75t_L g3538 ( 
.A(n_2895),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3092),
.Y(n_3539)
);

AOI22xp33_ASAP7_75t_SL g3540 ( 
.A1(n_3152),
.A2(n_2461),
.B1(n_2574),
.B2(n_2551),
.Y(n_3540)
);

BUFx12f_ASAP7_75t_L g3541 ( 
.A(n_2896),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3076),
.B(n_2465),
.Y(n_3542)
);

CKINVDCx11_ASAP7_75t_R g3543 ( 
.A(n_3228),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3207),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3231),
.Y(n_3545)
);

BUFx12f_ASAP7_75t_L g3546 ( 
.A(n_2911),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3242),
.Y(n_3547)
);

AOI22xp5_ASAP7_75t_L g3548 ( 
.A1(n_3221),
.A2(n_2495),
.B1(n_2503),
.B2(n_2466),
.Y(n_3548)
);

INVxp67_ASAP7_75t_SL g3549 ( 
.A(n_3168),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_2922),
.B(n_2523),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_2948),
.B(n_3238),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3141),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3243),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3250),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3266),
.Y(n_3555)
);

CKINVDCx20_ASAP7_75t_R g3556 ( 
.A(n_2996),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_3088),
.Y(n_3557)
);

CKINVDCx5p33_ASAP7_75t_R g3558 ( 
.A(n_2984),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3137),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3137),
.Y(n_3560)
);

INVx8_ASAP7_75t_L g3561 ( 
.A(n_2854),
.Y(n_3561)
);

BUFx6f_ASAP7_75t_L g3562 ( 
.A(n_2880),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3094),
.Y(n_3563)
);

BUFx2_ASAP7_75t_L g3564 ( 
.A(n_2852),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3094),
.Y(n_3565)
);

BUFx6f_ASAP7_75t_L g3566 ( 
.A(n_2880),
.Y(n_3566)
);

AOI22xp33_ASAP7_75t_L g3567 ( 
.A1(n_3245),
.A2(n_2754),
.B1(n_2575),
.B2(n_2574),
.Y(n_3567)
);

CKINVDCx11_ASAP7_75t_R g3568 ( 
.A(n_2907),
.Y(n_3568)
);

BUFx3_ASAP7_75t_L g3569 ( 
.A(n_3035),
.Y(n_3569)
);

CKINVDCx20_ASAP7_75t_R g3570 ( 
.A(n_3087),
.Y(n_3570)
);

INVx6_ASAP7_75t_L g3571 ( 
.A(n_3104),
.Y(n_3571)
);

AO22x1_ASAP7_75t_L g3572 ( 
.A1(n_2888),
.A2(n_2575),
.B1(n_2574),
.B2(n_2692),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_2901),
.Y(n_3573)
);

OAI22xp5_ASAP7_75t_L g3574 ( 
.A1(n_3186),
.A2(n_2575),
.B1(n_2754),
.B2(n_2694),
.Y(n_3574)
);

AOI22xp33_ASAP7_75t_L g3575 ( 
.A1(n_3222),
.A2(n_2754),
.B1(n_2694),
.B2(n_2692),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3006),
.B(n_253),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_2905),
.Y(n_3577)
);

AOI22xp33_ASAP7_75t_SL g3578 ( 
.A1(n_3034),
.A2(n_2694),
.B1(n_256),
.B2(n_254),
.Y(n_3578)
);

AND2x4_ASAP7_75t_L g3579 ( 
.A(n_2999),
.B(n_254),
.Y(n_3579)
);

INVx6_ASAP7_75t_L g3580 ( 
.A(n_3095),
.Y(n_3580)
);

BUFx8_ASAP7_75t_L g3581 ( 
.A(n_3211),
.Y(n_3581)
);

AOI22xp33_ASAP7_75t_L g3582 ( 
.A1(n_3240),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_2908),
.Y(n_3583)
);

BUFx3_ASAP7_75t_L g3584 ( 
.A(n_3051),
.Y(n_3584)
);

AOI22xp33_ASAP7_75t_L g3585 ( 
.A1(n_3265),
.A2(n_259),
.B1(n_255),
.B2(n_257),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3099),
.Y(n_3586)
);

INVx3_ASAP7_75t_L g3587 ( 
.A(n_2882),
.Y(n_3587)
);

BUFx2_ASAP7_75t_L g3588 ( 
.A(n_2925),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3099),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_3006),
.B(n_259),
.Y(n_3590)
);

INVx2_ASAP7_75t_SL g3591 ( 
.A(n_2925),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3102),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3102),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3110),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_2987),
.B(n_260),
.Y(n_3595)
);

INVx6_ASAP7_75t_L g3596 ( 
.A(n_3053),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_3036),
.Y(n_3597)
);

AOI22xp33_ASAP7_75t_L g3598 ( 
.A1(n_3274),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_3598)
);

BUFx3_ASAP7_75t_L g3599 ( 
.A(n_2920),
.Y(n_3599)
);

BUFx2_ASAP7_75t_L g3600 ( 
.A(n_3206),
.Y(n_3600)
);

OAI22xp5_ASAP7_75t_L g3601 ( 
.A1(n_3205),
.A2(n_264),
.B1(n_261),
.B2(n_263),
.Y(n_3601)
);

OAI22xp5_ASAP7_75t_L g3602 ( 
.A1(n_3101),
.A2(n_267),
.B1(n_264),
.B2(n_265),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3110),
.Y(n_3603)
);

AOI22xp33_ASAP7_75t_SL g3604 ( 
.A1(n_3034),
.A2(n_271),
.B1(n_268),
.B2(n_270),
.Y(n_3604)
);

NAND2x1p5_ASAP7_75t_L g3605 ( 
.A(n_2888),
.B(n_270),
.Y(n_3605)
);

CKINVDCx6p67_ASAP7_75t_R g3606 ( 
.A(n_2943),
.Y(n_3606)
);

BUFx2_ASAP7_75t_L g3607 ( 
.A(n_3105),
.Y(n_3607)
);

CKINVDCx11_ASAP7_75t_R g3608 ( 
.A(n_2921),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3131),
.A2(n_272),
.B(n_273),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3118),
.Y(n_3610)
);

INVx2_ASAP7_75t_SL g3611 ( 
.A(n_3117),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3118),
.Y(n_3612)
);

INVx1_ASAP7_75t_SL g3613 ( 
.A(n_2950),
.Y(n_3613)
);

CKINVDCx5p33_ASAP7_75t_R g3614 ( 
.A(n_2936),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3122),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3122),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_SL g3617 ( 
.A(n_2943),
.B(n_272),
.Y(n_3617)
);

AOI22xp33_ASAP7_75t_SL g3618 ( 
.A1(n_3055),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3044),
.Y(n_3619)
);

INVx6_ASAP7_75t_L g3620 ( 
.A(n_3060),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3141),
.Y(n_3621)
);

OR2x2_ASAP7_75t_L g3622 ( 
.A(n_2985),
.B(n_274),
.Y(n_3622)
);

HB1xp67_ASAP7_75t_L g3623 ( 
.A(n_3113),
.Y(n_3623)
);

CKINVDCx20_ASAP7_75t_R g3624 ( 
.A(n_2936),
.Y(n_3624)
);

AOI22xp33_ASAP7_75t_L g3625 ( 
.A1(n_3176),
.A2(n_278),
.B1(n_275),
.B2(n_277),
.Y(n_3625)
);

AOI22xp33_ASAP7_75t_SL g3626 ( 
.A1(n_3055),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_3626)
);

OR2x2_ASAP7_75t_L g3627 ( 
.A(n_2879),
.B(n_280),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3050),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3148),
.Y(n_3629)
);

BUFx6f_ASAP7_75t_SL g3630 ( 
.A(n_3112),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3148),
.Y(n_3631)
);

AOI22xp33_ASAP7_75t_SL g3632 ( 
.A1(n_3115),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_3632)
);

BUFx12f_ASAP7_75t_L g3633 ( 
.A(n_3012),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3154),
.Y(n_3634)
);

BUFx10_ASAP7_75t_L g3635 ( 
.A(n_3040),
.Y(n_3635)
);

AOI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_3134),
.A2(n_281),
.B(n_283),
.Y(n_3636)
);

BUFx3_ASAP7_75t_L g3637 ( 
.A(n_3079),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_3522),
.B(n_3466),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3389),
.Y(n_3639)
);

AOI22xp33_ASAP7_75t_SL g3640 ( 
.A1(n_3345),
.A2(n_3010),
.B1(n_2999),
.B2(n_3000),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3544),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3454),
.Y(n_3642)
);

OAI22xp5_ASAP7_75t_L g3643 ( 
.A1(n_3310),
.A2(n_3283),
.B1(n_3314),
.B2(n_3300),
.Y(n_3643)
);

AOI22xp33_ASAP7_75t_L g3644 ( 
.A1(n_3295),
.A2(n_3112),
.B1(n_2971),
.B2(n_3135),
.Y(n_3644)
);

HB1xp67_ASAP7_75t_L g3645 ( 
.A(n_3284),
.Y(n_3645)
);

AOI22xp33_ASAP7_75t_L g3646 ( 
.A1(n_3288),
.A2(n_3135),
.B1(n_2881),
.B2(n_2893),
.Y(n_3646)
);

INVxp67_ASAP7_75t_L g3647 ( 
.A(n_3279),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3545),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3482),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3547),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3553),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_3451),
.B(n_3040),
.Y(n_3652)
);

OAI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3316),
.A2(n_2999),
.B1(n_3010),
.B2(n_3000),
.Y(n_3653)
);

BUFx4f_ASAP7_75t_L g3654 ( 
.A(n_3396),
.Y(n_3654)
);

INVx4_ASAP7_75t_L g3655 ( 
.A(n_3614),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3488),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3554),
.Y(n_3657)
);

AOI22xp33_ASAP7_75t_L g3658 ( 
.A1(n_3291),
.A2(n_2970),
.B1(n_2956),
.B2(n_2894),
.Y(n_3658)
);

AOI22xp33_ASAP7_75t_L g3659 ( 
.A1(n_3317),
.A2(n_2894),
.B1(n_3161),
.B2(n_3150),
.Y(n_3659)
);

BUFx2_ASAP7_75t_L g3660 ( 
.A(n_3624),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3503),
.B(n_3551),
.Y(n_3661)
);

AOI22xp33_ASAP7_75t_L g3662 ( 
.A1(n_3336),
.A2(n_3246),
.B1(n_3179),
.B2(n_3262),
.Y(n_3662)
);

NAND3xp33_ASAP7_75t_L g3663 ( 
.A(n_3509),
.B(n_2915),
.C(n_2939),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3490),
.Y(n_3664)
);

OAI21xp5_ASAP7_75t_SL g3665 ( 
.A1(n_3286),
.A2(n_3003),
.B(n_2972),
.Y(n_3665)
);

OAI21xp33_ASAP7_75t_L g3666 ( 
.A1(n_3441),
.A2(n_3223),
.B(n_3184),
.Y(n_3666)
);

AOI22xp33_ASAP7_75t_L g3667 ( 
.A1(n_3287),
.A2(n_3262),
.B1(n_3267),
.B2(n_3007),
.Y(n_3667)
);

AOI22xp33_ASAP7_75t_L g3668 ( 
.A1(n_3287),
.A2(n_3016),
.B1(n_2864),
.B2(n_3153),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3285),
.Y(n_3669)
);

AOI22xp33_ASAP7_75t_SL g3670 ( 
.A1(n_3630),
.A2(n_3010),
.B1(n_3014),
.B2(n_3000),
.Y(n_3670)
);

AND2x2_ASAP7_75t_L g3671 ( 
.A(n_3370),
.B(n_2887),
.Y(n_3671)
);

AOI22xp33_ASAP7_75t_L g3672 ( 
.A1(n_3287),
.A2(n_2864),
.B1(n_3259),
.B2(n_3241),
.Y(n_3672)
);

AOI22xp33_ASAP7_75t_L g3673 ( 
.A1(n_3630),
.A2(n_3259),
.B1(n_3241),
.B2(n_3017),
.Y(n_3673)
);

AOI22xp33_ASAP7_75t_L g3674 ( 
.A1(n_3372),
.A2(n_3259),
.B1(n_2943),
.B2(n_3042),
.Y(n_3674)
);

INVx3_ASAP7_75t_L g3675 ( 
.A(n_3528),
.Y(n_3675)
);

AND2x2_ASAP7_75t_L g3676 ( 
.A(n_3576),
.B(n_3590),
.Y(n_3676)
);

OAI21xp5_ASAP7_75t_SL g3677 ( 
.A1(n_3292),
.A2(n_3227),
.B(n_3119),
.Y(n_3677)
);

OAI21xp5_ASAP7_75t_SL g3678 ( 
.A1(n_3280),
.A2(n_3119),
.B(n_3107),
.Y(n_3678)
);

OAI22xp33_ASAP7_75t_L g3679 ( 
.A1(n_3301),
.A2(n_3014),
.B1(n_3042),
.B2(n_3012),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3294),
.Y(n_3680)
);

AOI22xp33_ASAP7_75t_SL g3681 ( 
.A1(n_3353),
.A2(n_3014),
.B1(n_3042),
.B2(n_2944),
.Y(n_3681)
);

AOI22xp33_ASAP7_75t_SL g3682 ( 
.A1(n_3447),
.A2(n_2944),
.B1(n_2969),
.B2(n_2951),
.Y(n_3682)
);

AOI22xp33_ASAP7_75t_L g3683 ( 
.A1(n_3395),
.A2(n_2906),
.B1(n_2927),
.B2(n_3072),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_3408),
.B(n_3333),
.Y(n_3684)
);

AOI22xp33_ASAP7_75t_SL g3685 ( 
.A1(n_3635),
.A2(n_2951),
.B1(n_2974),
.B2(n_2969),
.Y(n_3685)
);

BUFx4f_ASAP7_75t_SL g3686 ( 
.A(n_3278),
.Y(n_3686)
);

INVx4_ASAP7_75t_L g3687 ( 
.A(n_3384),
.Y(n_3687)
);

AOI22xp33_ASAP7_75t_L g3688 ( 
.A1(n_3400),
.A2(n_2902),
.B1(n_3109),
.B2(n_3091),
.Y(n_3688)
);

AOI22xp5_ASAP7_75t_L g3689 ( 
.A1(n_3349),
.A2(n_2844),
.B1(n_3236),
.B2(n_3233),
.Y(n_3689)
);

AOI22xp33_ASAP7_75t_SL g3690 ( 
.A1(n_3635),
.A2(n_3457),
.B1(n_3318),
.B2(n_3564),
.Y(n_3690)
);

NOR2xp33_ASAP7_75t_L g3691 ( 
.A(n_3379),
.B(n_3458),
.Y(n_3691)
);

INVx3_ASAP7_75t_L g3692 ( 
.A(n_3528),
.Y(n_3692)
);

AOI22xp33_ASAP7_75t_L g3693 ( 
.A1(n_3445),
.A2(n_2855),
.B1(n_3043),
.B2(n_3019),
.Y(n_3693)
);

CKINVDCx5p33_ASAP7_75t_R g3694 ( 
.A(n_3386),
.Y(n_3694)
);

HB1xp67_ASAP7_75t_L g3695 ( 
.A(n_3588),
.Y(n_3695)
);

AOI22xp33_ASAP7_75t_L g3696 ( 
.A1(n_3432),
.A2(n_3425),
.B1(n_3465),
.B2(n_3421),
.Y(n_3696)
);

AOI22xp33_ASAP7_75t_SL g3697 ( 
.A1(n_3335),
.A2(n_2989),
.B1(n_2974),
.B2(n_3107),
.Y(n_3697)
);

AOI22xp33_ASAP7_75t_L g3698 ( 
.A1(n_3360),
.A2(n_3230),
.B1(n_3232),
.B2(n_2848),
.Y(n_3698)
);

AOI22xp33_ASAP7_75t_L g3699 ( 
.A1(n_3424),
.A2(n_3244),
.B1(n_3272),
.B2(n_3254),
.Y(n_3699)
);

AOI22xp33_ASAP7_75t_SL g3700 ( 
.A1(n_3320),
.A2(n_2989),
.B1(n_2960),
.B2(n_2983),
.Y(n_3700)
);

AOI222xp33_ASAP7_75t_L g3701 ( 
.A1(n_3303),
.A2(n_3124),
.B1(n_3173),
.B2(n_3247),
.C1(n_3163),
.C2(n_3154),
.Y(n_3701)
);

OAI22xp5_ASAP7_75t_L g3702 ( 
.A1(n_3319),
.A2(n_3083),
.B1(n_3089),
.B2(n_3066),
.Y(n_3702)
);

AOI22xp33_ASAP7_75t_L g3703 ( 
.A1(n_3429),
.A2(n_3163),
.B1(n_2941),
.B2(n_2952),
.Y(n_3703)
);

AOI22xp33_ASAP7_75t_SL g3704 ( 
.A1(n_3355),
.A2(n_2960),
.B1(n_2983),
.B2(n_2932),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3297),
.Y(n_3705)
);

AOI22xp33_ASAP7_75t_L g3706 ( 
.A1(n_3383),
.A2(n_2961),
.B1(n_3062),
.B2(n_2994),
.Y(n_3706)
);

AOI22xp33_ASAP7_75t_L g3707 ( 
.A1(n_3406),
.A2(n_2994),
.B1(n_2932),
.B2(n_2909),
.Y(n_3707)
);

AOI22xp33_ASAP7_75t_L g3708 ( 
.A1(n_3427),
.A2(n_2909),
.B1(n_2916),
.B2(n_2897),
.Y(n_3708)
);

OAI22xp5_ASAP7_75t_SL g3709 ( 
.A1(n_3374),
.A2(n_2916),
.B1(n_2897),
.B2(n_3181),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3506),
.Y(n_3710)
);

AOI22xp33_ASAP7_75t_L g3711 ( 
.A1(n_3469),
.A2(n_3093),
.B1(n_3097),
.B2(n_3090),
.Y(n_3711)
);

CKINVDCx5p33_ASAP7_75t_R g3712 ( 
.A(n_3467),
.Y(n_3712)
);

AOI22xp33_ASAP7_75t_L g3713 ( 
.A1(n_3405),
.A2(n_3120),
.B1(n_3111),
.B2(n_3086),
.Y(n_3713)
);

OAI22xp5_ASAP7_75t_L g3714 ( 
.A1(n_3368),
.A2(n_3198),
.B1(n_3086),
.B2(n_3160),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3306),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3557),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3309),
.Y(n_3717)
);

OAI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_3315),
.A2(n_3160),
.B1(n_3165),
.B2(n_3157),
.Y(n_3718)
);

OAI22xp5_ASAP7_75t_L g3719 ( 
.A1(n_3334),
.A2(n_3165),
.B1(n_3194),
.B2(n_3157),
.Y(n_3719)
);

AOI22xp33_ASAP7_75t_L g3720 ( 
.A1(n_3403),
.A2(n_3194),
.B1(n_3261),
.B2(n_3260),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3555),
.B(n_2954),
.Y(n_3721)
);

INVx8_ASAP7_75t_L g3722 ( 
.A(n_3384),
.Y(n_3722)
);

BUFx12f_ASAP7_75t_L g3723 ( 
.A(n_3278),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_3346),
.B(n_284),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3560),
.Y(n_3725)
);

AOI22xp33_ASAP7_75t_SL g3726 ( 
.A1(n_3355),
.A2(n_3261),
.B1(n_3260),
.B2(n_3226),
.Y(n_3726)
);

AOI22xp33_ASAP7_75t_L g3727 ( 
.A1(n_3347),
.A2(n_3251),
.B1(n_3257),
.B2(n_3226),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3313),
.Y(n_3728)
);

AOI22xp33_ASAP7_75t_L g3729 ( 
.A1(n_3468),
.A2(n_3428),
.B1(n_3437),
.B2(n_3356),
.Y(n_3729)
);

AND2x2_ASAP7_75t_L g3730 ( 
.A(n_3350),
.B(n_285),
.Y(n_3730)
);

NOR2xp33_ASAP7_75t_L g3731 ( 
.A(n_3568),
.B(n_3608),
.Y(n_3731)
);

AO22x1_ASAP7_75t_L g3732 ( 
.A1(n_3307),
.A2(n_3185),
.B1(n_3202),
.B2(n_3169),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3535),
.B(n_2958),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3539),
.B(n_3257),
.Y(n_3734)
);

AOI22xp33_ASAP7_75t_L g3735 ( 
.A1(n_3431),
.A2(n_3225),
.B1(n_3108),
.B2(n_3209),
.Y(n_3735)
);

BUFx3_ASAP7_75t_L g3736 ( 
.A(n_3556),
.Y(n_3736)
);

AOI22xp33_ASAP7_75t_L g3737 ( 
.A1(n_3439),
.A2(n_3108),
.B1(n_3209),
.B2(n_3098),
.Y(n_3737)
);

OAI22xp5_ASAP7_75t_L g3738 ( 
.A1(n_3325),
.A2(n_3084),
.B1(n_3185),
.B2(n_3169),
.Y(n_3738)
);

OAI21xp5_ASAP7_75t_SL g3739 ( 
.A1(n_3363),
.A2(n_3147),
.B(n_3145),
.Y(n_3739)
);

AOI22xp33_ASAP7_75t_SL g3740 ( 
.A1(n_3311),
.A2(n_3239),
.B1(n_3108),
.B2(n_3209),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3324),
.B(n_3098),
.Y(n_3741)
);

AOI22xp33_ASAP7_75t_L g3742 ( 
.A1(n_3443),
.A2(n_3489),
.B1(n_3632),
.B2(n_3602),
.Y(n_3742)
);

AOI22xp33_ASAP7_75t_SL g3743 ( 
.A1(n_3311),
.A2(n_3239),
.B1(n_3108),
.B2(n_3209),
.Y(n_3743)
);

OAI21xp33_ASAP7_75t_L g3744 ( 
.A1(n_3444),
.A2(n_3147),
.B(n_3145),
.Y(n_3744)
);

AOI22xp33_ASAP7_75t_L g3745 ( 
.A1(n_3601),
.A2(n_3239),
.B1(n_3098),
.B2(n_3096),
.Y(n_3745)
);

OAI22xp5_ASAP7_75t_L g3746 ( 
.A1(n_3399),
.A2(n_3084),
.B1(n_3185),
.B2(n_3169),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3359),
.Y(n_3747)
);

AOI22xp33_ASAP7_75t_L g3748 ( 
.A1(n_3357),
.A2(n_3239),
.B1(n_3098),
.B2(n_3096),
.Y(n_3748)
);

CKINVDCx11_ASAP7_75t_R g3749 ( 
.A(n_3290),
.Y(n_3749)
);

OAI22xp5_ASAP7_75t_L g3750 ( 
.A1(n_3390),
.A2(n_3084),
.B1(n_3213),
.B2(n_3202),
.Y(n_3750)
);

AOI22xp33_ASAP7_75t_SL g3751 ( 
.A1(n_3579),
.A2(n_3183),
.B1(n_3190),
.B2(n_3077),
.Y(n_3751)
);

AOI22xp33_ASAP7_75t_L g3752 ( 
.A1(n_3343),
.A2(n_3183),
.B1(n_3190),
.B2(n_3077),
.Y(n_3752)
);

AND2x4_ASAP7_75t_L g3753 ( 
.A(n_3420),
.B(n_3422),
.Y(n_3753)
);

HB1xp67_ASAP7_75t_L g3754 ( 
.A(n_3500),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3375),
.Y(n_3755)
);

OAI22xp5_ASAP7_75t_L g3756 ( 
.A1(n_3380),
.A2(n_3213),
.B1(n_3202),
.B2(n_3273),
.Y(n_3756)
);

BUFx12f_ASAP7_75t_L g3757 ( 
.A(n_3463),
.Y(n_3757)
);

AOI22xp33_ASAP7_75t_SL g3758 ( 
.A1(n_3579),
.A2(n_3213),
.B1(n_3273),
.B2(n_3268),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3362),
.Y(n_3759)
);

INVx4_ASAP7_75t_L g3760 ( 
.A(n_3422),
.Y(n_3760)
);

AOI22xp33_ASAP7_75t_L g3761 ( 
.A1(n_3598),
.A2(n_3268),
.B1(n_2919),
.B2(n_2923),
.Y(n_3761)
);

INVxp67_ASAP7_75t_SL g3762 ( 
.A(n_3326),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3371),
.Y(n_3763)
);

OAI22xp5_ASAP7_75t_L g3764 ( 
.A1(n_3382),
.A2(n_3578),
.B1(n_3450),
.B2(n_3339),
.Y(n_3764)
);

AOI22xp33_ASAP7_75t_L g3765 ( 
.A1(n_3459),
.A2(n_3487),
.B1(n_3502),
.B2(n_3625),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3373),
.B(n_2918),
.Y(n_3766)
);

CKINVDCx5p33_ASAP7_75t_R g3767 ( 
.A(n_3281),
.Y(n_3767)
);

AND2x2_ASAP7_75t_L g3768 ( 
.A(n_3599),
.B(n_285),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3385),
.B(n_2918),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3461),
.B(n_2918),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3471),
.B(n_2919),
.Y(n_3771)
);

OAI222xp33_ASAP7_75t_L g3772 ( 
.A1(n_3604),
.A2(n_289),
.B1(n_291),
.B2(n_286),
.C1(n_288),
.C2(n_290),
.Y(n_3772)
);

OAI22xp5_ASAP7_75t_L g3773 ( 
.A1(n_3618),
.A2(n_3215),
.B1(n_3197),
.B2(n_2923),
.Y(n_3773)
);

AOI22xp33_ASAP7_75t_L g3774 ( 
.A1(n_3298),
.A2(n_2923),
.B1(n_2924),
.B2(n_2919),
.Y(n_3774)
);

AND2x2_ASAP7_75t_L g3775 ( 
.A(n_3289),
.B(n_286),
.Y(n_3775)
);

OAI21xp5_ASAP7_75t_SL g3776 ( 
.A1(n_3426),
.A2(n_2935),
.B(n_2924),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3479),
.Y(n_3777)
);

CKINVDCx11_ASAP7_75t_R g3778 ( 
.A(n_3302),
.Y(n_3778)
);

AOI22xp33_ASAP7_75t_L g3779 ( 
.A1(n_3364),
.A2(n_2935),
.B1(n_2953),
.B2(n_2924),
.Y(n_3779)
);

AOI22xp33_ASAP7_75t_SL g3780 ( 
.A1(n_3571),
.A2(n_2953),
.B1(n_2957),
.B2(n_2935),
.Y(n_3780)
);

AOI22xp33_ASAP7_75t_L g3781 ( 
.A1(n_3626),
.A2(n_2957),
.B1(n_2978),
.B2(n_2953),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3481),
.Y(n_3782)
);

AOI22xp33_ASAP7_75t_SL g3783 ( 
.A1(n_3571),
.A2(n_2978),
.B1(n_2979),
.B2(n_2957),
.Y(n_3783)
);

AND2x2_ASAP7_75t_L g3784 ( 
.A(n_3277),
.B(n_288),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3494),
.B(n_2978),
.Y(n_3785)
);

OAI22xp5_ASAP7_75t_L g3786 ( 
.A1(n_3605),
.A2(n_3155),
.B1(n_3156),
.B2(n_3146),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3329),
.Y(n_3787)
);

AOI22xp33_ASAP7_75t_L g3788 ( 
.A1(n_3452),
.A2(n_2982),
.B1(n_3018),
.B2(n_2979),
.Y(n_3788)
);

NOR2xp33_ASAP7_75t_SL g3789 ( 
.A(n_3388),
.B(n_2979),
.Y(n_3789)
);

HB1xp67_ASAP7_75t_L g3790 ( 
.A(n_3613),
.Y(n_3790)
);

BUFx3_ASAP7_75t_L g3791 ( 
.A(n_3570),
.Y(n_3791)
);

INVx1_ASAP7_75t_SL g3792 ( 
.A(n_3476),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3496),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3573),
.Y(n_3794)
);

BUFx4f_ASAP7_75t_L g3795 ( 
.A(n_3296),
.Y(n_3795)
);

BUFx2_ASAP7_75t_L g3796 ( 
.A(n_3581),
.Y(n_3796)
);

INVx4_ASAP7_75t_L g3797 ( 
.A(n_3422),
.Y(n_3797)
);

OAI22xp33_ASAP7_75t_SL g3798 ( 
.A1(n_3519),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_3798)
);

AOI22xp33_ASAP7_75t_SL g3799 ( 
.A1(n_3367),
.A2(n_3410),
.B1(n_3549),
.B2(n_3531),
.Y(n_3799)
);

OAI21xp5_ASAP7_75t_SL g3800 ( 
.A1(n_3430),
.A2(n_3018),
.B(n_2982),
.Y(n_3800)
);

OAI22x1_ASAP7_75t_SL g3801 ( 
.A1(n_3415),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_3801)
);

CKINVDCx5p33_ASAP7_75t_R g3802 ( 
.A(n_3365),
.Y(n_3802)
);

INVx2_ASAP7_75t_L g3803 ( 
.A(n_3577),
.Y(n_3803)
);

AOI211xp5_ASAP7_75t_L g3804 ( 
.A1(n_3505),
.A2(n_3018),
.B(n_3025),
.C(n_2982),
.Y(n_3804)
);

INVx1_ASAP7_75t_SL g3805 ( 
.A(n_3480),
.Y(n_3805)
);

INVx3_ASAP7_75t_L g3806 ( 
.A(n_3508),
.Y(n_3806)
);

OAI22xp5_ASAP7_75t_L g3807 ( 
.A1(n_3453),
.A2(n_3215),
.B1(n_3197),
.B2(n_3039),
.Y(n_3807)
);

AOI22xp33_ASAP7_75t_L g3808 ( 
.A1(n_3515),
.A2(n_3039),
.B1(n_3048),
.B2(n_3025),
.Y(n_3808)
);

OAI222xp33_ASAP7_75t_L g3809 ( 
.A1(n_3497),
.A2(n_296),
.B1(n_298),
.B2(n_292),
.C1(n_294),
.C2(n_297),
.Y(n_3809)
);

AOI22xp33_ASAP7_75t_L g3810 ( 
.A1(n_3521),
.A2(n_3039),
.B1(n_3048),
.B2(n_3025),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3499),
.B(n_3048),
.Y(n_3811)
);

OAI22xp5_ASAP7_75t_SL g3812 ( 
.A1(n_3299),
.A2(n_3071),
.B1(n_3078),
.B2(n_3065),
.Y(n_3812)
);

AOI22xp33_ASAP7_75t_L g3813 ( 
.A1(n_3537),
.A2(n_3071),
.B1(n_3078),
.B2(n_3065),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3512),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_3293),
.B(n_296),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3532),
.B(n_3330),
.Y(n_3816)
);

INVx4_ASAP7_75t_L g3817 ( 
.A(n_3508),
.Y(n_3817)
);

OAI22xp5_ASAP7_75t_L g3818 ( 
.A1(n_3473),
.A2(n_3071),
.B1(n_3078),
.B2(n_3065),
.Y(n_3818)
);

BUFx2_ASAP7_75t_L g3819 ( 
.A(n_3581),
.Y(n_3819)
);

AOI22xp33_ASAP7_75t_SL g3820 ( 
.A1(n_3323),
.A2(n_3132),
.B1(n_3138),
.B2(n_3125),
.Y(n_3820)
);

HB1xp67_ASAP7_75t_L g3821 ( 
.A(n_3623),
.Y(n_3821)
);

AOI22xp33_ASAP7_75t_L g3822 ( 
.A1(n_3526),
.A2(n_3132),
.B1(n_3138),
.B2(n_3125),
.Y(n_3822)
);

AOI22xp33_ASAP7_75t_L g3823 ( 
.A1(n_3543),
.A2(n_3132),
.B1(n_3138),
.B2(n_3125),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3534),
.B(n_3142),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3559),
.Y(n_3825)
);

OAI22xp33_ASAP7_75t_SL g3826 ( 
.A1(n_3519),
.A2(n_300),
.B1(n_297),
.B2(n_299),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3563),
.Y(n_3827)
);

AOI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3419),
.A2(n_3146),
.B1(n_3155),
.B2(n_3142),
.Y(n_3828)
);

BUFx6f_ASAP7_75t_L g3829 ( 
.A(n_3354),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3565),
.Y(n_3830)
);

NOR2xp33_ASAP7_75t_L g3831 ( 
.A(n_3462),
.B(n_299),
.Y(n_3831)
);

AOI22xp33_ASAP7_75t_SL g3832 ( 
.A1(n_3323),
.A2(n_3146),
.B1(n_3155),
.B2(n_3142),
.Y(n_3832)
);

OAI22xp33_ASAP7_75t_L g3833 ( 
.A1(n_3393),
.A2(n_3166),
.B1(n_3171),
.B2(n_3156),
.Y(n_3833)
);

AOI22xp33_ASAP7_75t_SL g3834 ( 
.A1(n_3393),
.A2(n_3166),
.B1(n_3171),
.B2(n_3156),
.Y(n_3834)
);

NOR2xp33_ASAP7_75t_L g3835 ( 
.A(n_3462),
.B(n_300),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3583),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3597),
.Y(n_3837)
);

OAI22xp5_ASAP7_75t_L g3838 ( 
.A1(n_3460),
.A2(n_3171),
.B1(n_3175),
.B2(n_3166),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3586),
.Y(n_3839)
);

AND2x2_ASAP7_75t_L g3840 ( 
.A(n_3637),
.B(n_301),
.Y(n_3840)
);

AOI22xp33_ASAP7_75t_SL g3841 ( 
.A1(n_3420),
.A2(n_3182),
.B1(n_3197),
.B2(n_3175),
.Y(n_3841)
);

HB1xp67_ASAP7_75t_L g3842 ( 
.A(n_3589),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3592),
.B(n_3175),
.Y(n_3843)
);

BUFx2_ASAP7_75t_SL g3844 ( 
.A(n_3511),
.Y(n_3844)
);

AOI22xp33_ASAP7_75t_SL g3845 ( 
.A1(n_3351),
.A2(n_3215),
.B1(n_3182),
.B2(n_3269),
.Y(n_3845)
);

INVx4_ASAP7_75t_L g3846 ( 
.A(n_3508),
.Y(n_3846)
);

OAI21xp5_ASAP7_75t_SL g3847 ( 
.A1(n_3312),
.A2(n_3182),
.B(n_3269),
.Y(n_3847)
);

INVx4_ASAP7_75t_L g3848 ( 
.A(n_3464),
.Y(n_3848)
);

OAI21xp5_ASAP7_75t_SL g3849 ( 
.A1(n_3321),
.A2(n_3269),
.B(n_302),
.Y(n_3849)
);

NOR2xp33_ASAP7_75t_L g3850 ( 
.A(n_3354),
.B(n_3409),
.Y(n_3850)
);

AOI22xp5_ASAP7_75t_L g3851 ( 
.A1(n_3413),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_3851)
);

AOI22xp33_ASAP7_75t_L g3852 ( 
.A1(n_3585),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_3852)
);

OAI22xp5_ASAP7_75t_L g3853 ( 
.A1(n_3518),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_3853)
);

NOR3xp33_ASAP7_75t_SL g3854 ( 
.A(n_3558),
.B(n_308),
.C(n_309),
.Y(n_3854)
);

AOI211xp5_ASAP7_75t_L g3855 ( 
.A1(n_3483),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_3855)
);

BUFx6f_ASAP7_75t_L g3856 ( 
.A(n_3344),
.Y(n_3856)
);

CKINVDCx20_ASAP7_75t_R g3857 ( 
.A(n_3392),
.Y(n_3857)
);

AOI22xp33_ASAP7_75t_L g3858 ( 
.A1(n_3627),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_3858)
);

OAI22xp5_ASAP7_75t_L g3859 ( 
.A1(n_3527),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.Y(n_3859)
);

AOI22xp33_ASAP7_75t_SL g3860 ( 
.A1(n_3435),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_3860)
);

OAI21xp5_ASAP7_75t_SL g3861 ( 
.A1(n_3540),
.A2(n_316),
.B(n_317),
.Y(n_3861)
);

OAI22xp33_ASAP7_75t_L g3862 ( 
.A1(n_3622),
.A2(n_322),
.B1(n_319),
.B2(n_321),
.Y(n_3862)
);

OAI22xp5_ASAP7_75t_L g3863 ( 
.A1(n_3358),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_3863)
);

INVx4_ASAP7_75t_L g3864 ( 
.A(n_3464),
.Y(n_3864)
);

AOI22xp33_ASAP7_75t_L g3865 ( 
.A1(n_3582),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_3865)
);

AOI22xp5_ASAP7_75t_L g3866 ( 
.A1(n_3456),
.A2(n_3423),
.B1(n_3536),
.B2(n_3485),
.Y(n_3866)
);

AOI22xp33_ASAP7_75t_L g3867 ( 
.A1(n_3609),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_3867)
);

AOI22xp33_ASAP7_75t_L g3868 ( 
.A1(n_3636),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3619),
.Y(n_3869)
);

INVx2_ASAP7_75t_L g3870 ( 
.A(n_3628),
.Y(n_3870)
);

OAI22xp33_ASAP7_75t_L g3871 ( 
.A1(n_3440),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_3871)
);

AOI22xp33_ASAP7_75t_SL g3872 ( 
.A1(n_3435),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_3872)
);

OAI21xp5_ASAP7_75t_SL g3873 ( 
.A1(n_3337),
.A2(n_332),
.B(n_334),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3593),
.Y(n_3874)
);

CKINVDCx5p33_ASAP7_75t_R g3875 ( 
.A(n_3305),
.Y(n_3875)
);

BUFx2_ASAP7_75t_L g3876 ( 
.A(n_3448),
.Y(n_3876)
);

AOI22xp33_ASAP7_75t_L g3877 ( 
.A1(n_3307),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_3877)
);

AOI22xp33_ASAP7_75t_SL g3878 ( 
.A1(n_3495),
.A2(n_3587),
.B1(n_3507),
.B2(n_3342),
.Y(n_3878)
);

OAI22xp5_ASAP7_75t_L g3879 ( 
.A1(n_3358),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_3879)
);

AOI22xp33_ASAP7_75t_SL g3880 ( 
.A1(n_3495),
.A2(n_3587),
.B1(n_3507),
.B2(n_3342),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3594),
.B(n_339),
.Y(n_3881)
);

INVx3_ASAP7_75t_L g3882 ( 
.A(n_3401),
.Y(n_3882)
);

INVx3_ASAP7_75t_L g3883 ( 
.A(n_3401),
.Y(n_3883)
);

BUFx12f_ASAP7_75t_L g3884 ( 
.A(n_3282),
.Y(n_3884)
);

AOI22xp33_ASAP7_75t_L g3885 ( 
.A1(n_3477),
.A2(n_342),
.B1(n_339),
.B2(n_341),
.Y(n_3885)
);

AOI22xp5_ASAP7_75t_L g3886 ( 
.A1(n_3498),
.A2(n_344),
.B1(n_341),
.B2(n_342),
.Y(n_3886)
);

AOI22xp33_ASAP7_75t_L g3887 ( 
.A1(n_3607),
.A2(n_3552),
.B1(n_3541),
.B2(n_3546),
.Y(n_3887)
);

AND2x2_ASAP7_75t_L g3888 ( 
.A(n_3591),
.B(n_3600),
.Y(n_3888)
);

INVx3_ASAP7_75t_L g3889 ( 
.A(n_3369),
.Y(n_3889)
);

OAI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3369),
.A2(n_347),
.B1(n_344),
.B2(n_345),
.Y(n_3890)
);

OAI22xp5_ASAP7_75t_L g3891 ( 
.A1(n_3606),
.A2(n_3510),
.B1(n_3436),
.B2(n_3620),
.Y(n_3891)
);

OAI22xp5_ASAP7_75t_L g3892 ( 
.A1(n_3620),
.A2(n_348),
.B1(n_345),
.B2(n_347),
.Y(n_3892)
);

OAI222xp33_ASAP7_75t_L g3893 ( 
.A1(n_3617),
.A2(n_350),
.B1(n_352),
.B2(n_348),
.C1(n_349),
.C2(n_351),
.Y(n_3893)
);

AOI22xp33_ASAP7_75t_SL g3894 ( 
.A1(n_3341),
.A2(n_353),
.B1(n_349),
.B2(n_350),
.Y(n_3894)
);

BUFx4f_ASAP7_75t_SL g3895 ( 
.A(n_3327),
.Y(n_3895)
);

AOI22xp33_ASAP7_75t_L g3896 ( 
.A1(n_3552),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_3896)
);

AOI22xp33_ASAP7_75t_SL g3897 ( 
.A1(n_3341),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_3897)
);

BUFx2_ASAP7_75t_L g3898 ( 
.A(n_3448),
.Y(n_3898)
);

AOI22xp33_ASAP7_75t_L g3899 ( 
.A1(n_3538),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_3899)
);

AOI22xp33_ASAP7_75t_SL g3900 ( 
.A1(n_3493),
.A2(n_362),
.B1(n_359),
.B2(n_361),
.Y(n_3900)
);

OAI21xp5_ASAP7_75t_SL g3901 ( 
.A1(n_3520),
.A2(n_362),
.B(n_364),
.Y(n_3901)
);

AOI22xp33_ASAP7_75t_L g3902 ( 
.A1(n_3595),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_3902)
);

INVx4_ASAP7_75t_SL g3903 ( 
.A(n_3344),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3603),
.B(n_365),
.Y(n_3904)
);

HB1xp67_ASAP7_75t_L g3905 ( 
.A(n_3610),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_L g3906 ( 
.A(n_3409),
.B(n_368),
.Y(n_3906)
);

AOI22xp33_ASAP7_75t_SL g3907 ( 
.A1(n_3366),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_3907)
);

INVx2_ASAP7_75t_L g3908 ( 
.A(n_3612),
.Y(n_3908)
);

HB1xp67_ASAP7_75t_L g3909 ( 
.A(n_3615),
.Y(n_3909)
);

INVx3_ASAP7_75t_L g3910 ( 
.A(n_3474),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3616),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3391),
.B(n_369),
.Y(n_3912)
);

OAI22xp33_ASAP7_75t_L g3913 ( 
.A1(n_3322),
.A2(n_3366),
.B1(n_3525),
.B2(n_3524),
.Y(n_3913)
);

AOI22xp33_ASAP7_75t_SL g3914 ( 
.A1(n_3561),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_3914)
);

OAI21xp5_ASAP7_75t_SL g3915 ( 
.A1(n_3407),
.A2(n_3486),
.B(n_3332),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3394),
.B(n_371),
.Y(n_3916)
);

NOR2xp33_ASAP7_75t_L g3917 ( 
.A(n_3455),
.B(n_372),
.Y(n_3917)
);

OAI22xp33_ASAP7_75t_L g3918 ( 
.A1(n_3474),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3398),
.B(n_3402),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3411),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3412),
.Y(n_3921)
);

AND2x2_ASAP7_75t_L g3922 ( 
.A(n_3491),
.B(n_839),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3414),
.B(n_375),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3418),
.Y(n_3924)
);

NOR2xp33_ASAP7_75t_L g3925 ( 
.A(n_3455),
.B(n_376),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3433),
.B(n_376),
.Y(n_3926)
);

CKINVDCx5p33_ASAP7_75t_R g3927 ( 
.A(n_3304),
.Y(n_3927)
);

BUFx12f_ASAP7_75t_L g3928 ( 
.A(n_3376),
.Y(n_3928)
);

OAI21xp5_ASAP7_75t_SL g3929 ( 
.A1(n_3308),
.A2(n_377),
.B(n_378),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3438),
.Y(n_3930)
);

AOI22xp33_ASAP7_75t_L g3931 ( 
.A1(n_3643),
.A2(n_3446),
.B1(n_3442),
.B2(n_3621),
.Y(n_3931)
);

AOI22xp5_ASAP7_75t_L g3932 ( 
.A1(n_3901),
.A2(n_3633),
.B1(n_3516),
.B2(n_3397),
.Y(n_3932)
);

AOI22xp33_ASAP7_75t_L g3933 ( 
.A1(n_3696),
.A2(n_3340),
.B1(n_3631),
.B2(n_3629),
.Y(n_3933)
);

AOI22xp33_ASAP7_75t_L g3934 ( 
.A1(n_3729),
.A2(n_3634),
.B1(n_3513),
.B2(n_3533),
.Y(n_3934)
);

AOI22xp33_ASAP7_75t_L g3935 ( 
.A1(n_3690),
.A2(n_3381),
.B1(n_3596),
.B2(n_3378),
.Y(n_3935)
);

AOI22xp33_ASAP7_75t_SL g3936 ( 
.A1(n_3709),
.A2(n_3561),
.B1(n_3524),
.B2(n_3480),
.Y(n_3936)
);

OAI221xp5_ASAP7_75t_L g3937 ( 
.A1(n_3665),
.A2(n_3611),
.B1(n_3501),
.B2(n_3529),
.C(n_3584),
.Y(n_3937)
);

AOI221xp5_ASAP7_75t_L g3938 ( 
.A1(n_3871),
.A2(n_3504),
.B1(n_3550),
.B2(n_3542),
.C(n_3348),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3816),
.B(n_3517),
.Y(n_3939)
);

OAI22xp5_ASAP7_75t_L g3940 ( 
.A1(n_3901),
.A2(n_3514),
.B1(n_3567),
.B2(n_3580),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_SL g3941 ( 
.A(n_3682),
.B(n_3878),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3684),
.B(n_3569),
.Y(n_3942)
);

AOI22xp33_ASAP7_75t_L g3943 ( 
.A1(n_3701),
.A2(n_3663),
.B1(n_3764),
.B2(n_3661),
.Y(n_3943)
);

AOI22xp33_ASAP7_75t_SL g3944 ( 
.A1(n_3654),
.A2(n_3596),
.B1(n_3331),
.B2(n_3361),
.Y(n_3944)
);

AOI22xp33_ASAP7_75t_L g3945 ( 
.A1(n_3663),
.A2(n_3638),
.B1(n_3644),
.B2(n_3646),
.Y(n_3945)
);

OAI221xp5_ASAP7_75t_L g3946 ( 
.A1(n_3665),
.A2(n_3416),
.B1(n_3580),
.B2(n_3484),
.C(n_3548),
.Y(n_3946)
);

OAI22xp5_ASAP7_75t_L g3947 ( 
.A1(n_3929),
.A2(n_3575),
.B1(n_3523),
.B2(n_3475),
.Y(n_3947)
);

AOI22xp33_ASAP7_75t_L g3948 ( 
.A1(n_3742),
.A2(n_3331),
.B1(n_3361),
.B2(n_3574),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3639),
.B(n_3344),
.Y(n_3949)
);

AOI22xp33_ASAP7_75t_L g3950 ( 
.A1(n_3658),
.A2(n_3328),
.B1(n_3404),
.B2(n_3377),
.Y(n_3950)
);

AOI22xp33_ASAP7_75t_L g3951 ( 
.A1(n_3662),
.A2(n_3404),
.B1(n_3449),
.B2(n_3377),
.Y(n_3951)
);

AOI22xp33_ASAP7_75t_SL g3952 ( 
.A1(n_3654),
.A2(n_3404),
.B1(n_3449),
.B2(n_3377),
.Y(n_3952)
);

OAI21xp33_ASAP7_75t_L g3953 ( 
.A1(n_3849),
.A2(n_3338),
.B(n_3470),
.Y(n_3953)
);

AOI22xp33_ASAP7_75t_L g3954 ( 
.A1(n_3666),
.A2(n_3449),
.B1(n_3478),
.B2(n_3472),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3641),
.B(n_3472),
.Y(n_3955)
);

AOI22xp33_ASAP7_75t_L g3956 ( 
.A1(n_3652),
.A2(n_3472),
.B1(n_3530),
.B2(n_3478),
.Y(n_3956)
);

OAI211xp5_ASAP7_75t_SL g3957 ( 
.A1(n_3866),
.A2(n_3387),
.B(n_3417),
.C(n_3352),
.Y(n_3957)
);

NOR3xp33_ASAP7_75t_L g3958 ( 
.A(n_3929),
.B(n_3572),
.C(n_3387),
.Y(n_3958)
);

AOI22xp33_ASAP7_75t_L g3959 ( 
.A1(n_3765),
.A2(n_3900),
.B1(n_3671),
.B2(n_3693),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_SL g3960 ( 
.A1(n_3762),
.A2(n_3478),
.B1(n_3562),
.B2(n_3530),
.Y(n_3960)
);

OAI22xp5_ASAP7_75t_L g3961 ( 
.A1(n_3861),
.A2(n_3530),
.B1(n_3566),
.B2(n_3562),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3648),
.B(n_3562),
.Y(n_3962)
);

BUFx2_ASAP7_75t_L g3963 ( 
.A(n_3695),
.Y(n_3963)
);

AOI22xp33_ASAP7_75t_L g3964 ( 
.A1(n_3918),
.A2(n_3566),
.B1(n_3417),
.B2(n_3492),
.Y(n_3964)
);

AOI22xp33_ASAP7_75t_L g3965 ( 
.A1(n_3688),
.A2(n_3566),
.B1(n_3434),
.B2(n_380),
.Y(n_3965)
);

AOI22xp33_ASAP7_75t_SL g3966 ( 
.A1(n_3702),
.A2(n_381),
.B1(n_378),
.B2(n_379),
.Y(n_3966)
);

OAI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_3861),
.A2(n_383),
.B1(n_379),
.B2(n_382),
.Y(n_3967)
);

AOI22xp33_ASAP7_75t_L g3968 ( 
.A1(n_3914),
.A2(n_385),
.B1(n_382),
.B2(n_383),
.Y(n_3968)
);

NOR3xp33_ASAP7_75t_SL g3969 ( 
.A(n_3849),
.B(n_386),
.C(n_387),
.Y(n_3969)
);

AOI22xp33_ASAP7_75t_L g3970 ( 
.A1(n_3676),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_3970)
);

AOI22xp33_ASAP7_75t_L g3971 ( 
.A1(n_3860),
.A2(n_392),
.B1(n_389),
.B2(n_390),
.Y(n_3971)
);

AOI221xp5_ASAP7_75t_L g3972 ( 
.A1(n_3862),
.A2(n_396),
.B1(n_393),
.B2(n_394),
.C(n_397),
.Y(n_3972)
);

OAI22xp5_ASAP7_75t_L g3973 ( 
.A1(n_3697),
.A2(n_398),
.B1(n_393),
.B2(n_397),
.Y(n_3973)
);

AOI22xp33_ASAP7_75t_L g3974 ( 
.A1(n_3872),
.A2(n_402),
.B1(n_399),
.B2(n_400),
.Y(n_3974)
);

AOI22xp33_ASAP7_75t_L g3975 ( 
.A1(n_3659),
.A2(n_403),
.B1(n_400),
.B2(n_402),
.Y(n_3975)
);

OAI22xp5_ASAP7_75t_L g3976 ( 
.A1(n_3685),
.A2(n_406),
.B1(n_403),
.B2(n_404),
.Y(n_3976)
);

AOI22xp33_ASAP7_75t_L g3977 ( 
.A1(n_3859),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3842),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3821),
.B(n_829),
.Y(n_3979)
);

AOI22xp33_ASAP7_75t_L g3980 ( 
.A1(n_3703),
.A2(n_411),
.B1(n_408),
.B2(n_410),
.Y(n_3980)
);

AOI22xp33_ASAP7_75t_L g3981 ( 
.A1(n_3853),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_3981)
);

AOI22xp33_ASAP7_75t_L g3982 ( 
.A1(n_3894),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_3982)
);

AOI22xp33_ASAP7_75t_L g3983 ( 
.A1(n_3897),
.A2(n_417),
.B1(n_413),
.B2(n_415),
.Y(n_3983)
);

AOI22xp33_ASAP7_75t_SL g3984 ( 
.A1(n_3891),
.A2(n_419),
.B1(n_415),
.B2(n_418),
.Y(n_3984)
);

AOI22xp33_ASAP7_75t_L g3985 ( 
.A1(n_3863),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_3985)
);

AOI22xp33_ASAP7_75t_L g3986 ( 
.A1(n_3879),
.A2(n_3890),
.B1(n_3892),
.B2(n_3907),
.Y(n_3986)
);

OAI222xp33_ASAP7_75t_L g3987 ( 
.A1(n_3799),
.A2(n_423),
.B1(n_425),
.B2(n_420),
.C1(n_422),
.C2(n_424),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_3642),
.Y(n_3988)
);

OAI22xp5_ASAP7_75t_L g3989 ( 
.A1(n_3667),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.Y(n_3989)
);

AOI22xp33_ASAP7_75t_SL g3990 ( 
.A1(n_3773),
.A2(n_429),
.B1(n_425),
.B2(n_426),
.Y(n_3990)
);

AOI22xp33_ASAP7_75t_L g3991 ( 
.A1(n_3877),
.A2(n_431),
.B1(n_426),
.B2(n_430),
.Y(n_3991)
);

AOI21xp5_ASAP7_75t_SL g3992 ( 
.A1(n_3653),
.A2(n_431),
.B(n_432),
.Y(n_3992)
);

AOI22xp33_ASAP7_75t_L g3993 ( 
.A1(n_3754),
.A2(n_436),
.B1(n_433),
.B2(n_435),
.Y(n_3993)
);

AOI22xp33_ASAP7_75t_L g3994 ( 
.A1(n_3645),
.A2(n_438),
.B1(n_435),
.B2(n_437),
.Y(n_3994)
);

AOI22xp33_ASAP7_75t_SL g3995 ( 
.A1(n_3812),
.A2(n_440),
.B1(n_437),
.B2(n_439),
.Y(n_3995)
);

AOI22xp33_ASAP7_75t_L g3996 ( 
.A1(n_3698),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_3996)
);

OAI22xp5_ASAP7_75t_L g3997 ( 
.A1(n_3855),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_3997)
);

INVx3_ASAP7_75t_L g3998 ( 
.A(n_3760),
.Y(n_3998)
);

OAI22xp33_ASAP7_75t_L g3999 ( 
.A1(n_3873),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.Y(n_3999)
);

AOI22xp33_ASAP7_75t_L g4000 ( 
.A1(n_3683),
.A2(n_447),
.B1(n_445),
.B2(n_446),
.Y(n_4000)
);

AOI22xp33_ASAP7_75t_L g4001 ( 
.A1(n_3899),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3649),
.Y(n_4002)
);

OAI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_3880),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.Y(n_4003)
);

OAI22xp5_ASAP7_75t_L g4004 ( 
.A1(n_3700),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_4004)
);

AND2x2_ASAP7_75t_L g4005 ( 
.A(n_3790),
.B(n_452),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3650),
.B(n_454),
.Y(n_4006)
);

AOI22xp33_ASAP7_75t_SL g4007 ( 
.A1(n_3876),
.A2(n_456),
.B1(n_454),
.B2(n_455),
.Y(n_4007)
);

AOI22xp33_ASAP7_75t_L g4008 ( 
.A1(n_3885),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3651),
.B(n_458),
.Y(n_4009)
);

AOI22xp33_ASAP7_75t_L g4010 ( 
.A1(n_3775),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_4010)
);

OAI22xp5_ASAP7_75t_L g4011 ( 
.A1(n_3677),
.A2(n_3668),
.B1(n_3704),
.B2(n_3726),
.Y(n_4011)
);

AND2x2_ASAP7_75t_L g4012 ( 
.A(n_3888),
.B(n_459),
.Y(n_4012)
);

OAI21xp5_ASAP7_75t_SL g4013 ( 
.A1(n_3915),
.A2(n_460),
.B(n_461),
.Y(n_4013)
);

AOI22xp33_ASAP7_75t_L g4014 ( 
.A1(n_3798),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_4014)
);

OAI222xp33_ASAP7_75t_L g4015 ( 
.A1(n_3681),
.A2(n_465),
.B1(n_467),
.B2(n_462),
.C1(n_463),
.C2(n_466),
.Y(n_4015)
);

AOI22xp5_ASAP7_75t_L g4016 ( 
.A1(n_3689),
.A2(n_468),
.B1(n_465),
.B2(n_466),
.Y(n_4016)
);

AOI21xp33_ASAP7_75t_L g4017 ( 
.A1(n_3677),
.A2(n_469),
.B(n_470),
.Y(n_4017)
);

OA21x2_ASAP7_75t_L g4018 ( 
.A1(n_3847),
.A2(n_823),
.B(n_469),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3657),
.B(n_472),
.Y(n_4019)
);

AOI22xp33_ASAP7_75t_SL g4020 ( 
.A1(n_3898),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_4020)
);

AOI22xp33_ASAP7_75t_L g4021 ( 
.A1(n_3826),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_SL g4022 ( 
.A(n_3804),
.B(n_476),
.Y(n_4022)
);

AOI22xp33_ASAP7_75t_L g4023 ( 
.A1(n_3840),
.A2(n_3699),
.B1(n_3852),
.B2(n_3713),
.Y(n_4023)
);

AOI22xp33_ASAP7_75t_SL g4024 ( 
.A1(n_3895),
.A2(n_479),
.B1(n_477),
.B2(n_478),
.Y(n_4024)
);

AOI22xp33_ASAP7_75t_L g4025 ( 
.A1(n_3865),
.A2(n_481),
.B1(n_478),
.B2(n_480),
.Y(n_4025)
);

AOI22xp5_ASAP7_75t_L g4026 ( 
.A1(n_3886),
.A2(n_487),
.B1(n_484),
.B2(n_486),
.Y(n_4026)
);

OAI22xp5_ASAP7_75t_L g4027 ( 
.A1(n_3707),
.A2(n_487),
.B1(n_484),
.B2(n_486),
.Y(n_4027)
);

AOI22xp33_ASAP7_75t_L g4028 ( 
.A1(n_3858),
.A2(n_490),
.B1(n_488),
.B2(n_489),
.Y(n_4028)
);

AOI22xp33_ASAP7_75t_L g4029 ( 
.A1(n_3905),
.A2(n_491),
.B1(n_488),
.B2(n_490),
.Y(n_4029)
);

AOI22xp33_ASAP7_75t_L g4030 ( 
.A1(n_3909),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3777),
.Y(n_4031)
);

AOI22xp33_ASAP7_75t_L g4032 ( 
.A1(n_3796),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_4032)
);

AOI22xp33_ASAP7_75t_L g4033 ( 
.A1(n_3819),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.Y(n_4033)
);

AOI22xp33_ASAP7_75t_SL g4034 ( 
.A1(n_3722),
.A2(n_499),
.B1(n_496),
.B2(n_497),
.Y(n_4034)
);

AOI221xp5_ASAP7_75t_L g4035 ( 
.A1(n_3801),
.A2(n_501),
.B1(n_499),
.B2(n_500),
.C(n_502),
.Y(n_4035)
);

AOI22xp5_ASAP7_75t_L g4036 ( 
.A1(n_3706),
.A2(n_503),
.B1(n_500),
.B2(n_502),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3782),
.B(n_503),
.Y(n_4037)
);

OAI21xp5_ASAP7_75t_SL g4038 ( 
.A1(n_3915),
.A2(n_505),
.B(n_506),
.Y(n_4038)
);

NAND3xp33_ASAP7_75t_L g4039 ( 
.A(n_3854),
.B(n_507),
.C(n_508),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3793),
.B(n_507),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3814),
.B(n_509),
.Y(n_4041)
);

AOI22xp33_ASAP7_75t_L g4042 ( 
.A1(n_3660),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3669),
.Y(n_4043)
);

AOI22xp33_ASAP7_75t_L g4044 ( 
.A1(n_3768),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.Y(n_4044)
);

OAI221xp5_ASAP7_75t_SL g4045 ( 
.A1(n_3800),
.A2(n_515),
.B1(n_513),
.B2(n_514),
.C(n_516),
.Y(n_4045)
);

BUFx3_ASAP7_75t_L g4046 ( 
.A(n_3722),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_3711),
.A2(n_516),
.B1(n_514),
.B2(n_515),
.Y(n_4047)
);

AOI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_3922),
.A2(n_519),
.B1(n_517),
.B2(n_518),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_3755),
.B(n_815),
.Y(n_4049)
);

AOI22xp33_ASAP7_75t_L g4050 ( 
.A1(n_3867),
.A2(n_519),
.B1(n_517),
.B2(n_518),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3787),
.B(n_809),
.Y(n_4051)
);

AOI22xp33_ASAP7_75t_L g4052 ( 
.A1(n_3868),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_4052)
);

OAI221xp5_ASAP7_75t_L g4053 ( 
.A1(n_3708),
.A2(n_524),
.B1(n_521),
.B2(n_523),
.C(n_525),
.Y(n_4053)
);

OAI22xp5_ASAP7_75t_L g4054 ( 
.A1(n_3781),
.A2(n_525),
.B1(n_523),
.B2(n_524),
.Y(n_4054)
);

AOI22xp33_ASAP7_75t_L g4055 ( 
.A1(n_3737),
.A2(n_528),
.B1(n_526),
.B2(n_527),
.Y(n_4055)
);

OAI222xp33_ASAP7_75t_L g4056 ( 
.A1(n_3686),
.A2(n_529),
.B1(n_530),
.B2(n_531),
.C1(n_532),
.C2(n_533),
.Y(n_4056)
);

INVx2_ASAP7_75t_L g4057 ( 
.A(n_3656),
.Y(n_4057)
);

OAI22xp5_ASAP7_75t_L g4058 ( 
.A1(n_3678),
.A2(n_534),
.B1(n_529),
.B2(n_531),
.Y(n_4058)
);

OAI222xp33_ASAP7_75t_L g4059 ( 
.A1(n_3640),
.A2(n_534),
.B1(n_535),
.B2(n_536),
.C1(n_537),
.C2(n_538),
.Y(n_4059)
);

AOI22xp33_ASAP7_75t_L g4060 ( 
.A1(n_3902),
.A2(n_538),
.B1(n_535),
.B2(n_536),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3680),
.Y(n_4061)
);

AOI22xp33_ASAP7_75t_L g4062 ( 
.A1(n_3896),
.A2(n_542),
.B1(n_539),
.B2(n_541),
.Y(n_4062)
);

AOI22xp33_ASAP7_75t_SL g4063 ( 
.A1(n_3722),
.A2(n_543),
.B1(n_539),
.B2(n_541),
.Y(n_4063)
);

AOI22xp33_ASAP7_75t_L g4064 ( 
.A1(n_3724),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3705),
.Y(n_4065)
);

AOI221xp5_ASAP7_75t_L g4066 ( 
.A1(n_3772),
.A2(n_547),
.B1(n_545),
.B2(n_546),
.C(n_548),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_3715),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3717),
.Y(n_4068)
);

OAI222xp33_ASAP7_75t_L g4069 ( 
.A1(n_3647),
.A2(n_548),
.B1(n_550),
.B2(n_551),
.C1(n_553),
.C2(n_554),
.Y(n_4069)
);

AOI22xp5_ASAP7_75t_L g4070 ( 
.A1(n_3678),
.A2(n_555),
.B1(n_551),
.B2(n_553),
.Y(n_4070)
);

OAI22xp5_ASAP7_75t_L g4071 ( 
.A1(n_3776),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.Y(n_4071)
);

AOI22xp33_ASAP7_75t_L g4072 ( 
.A1(n_3730),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3794),
.B(n_806),
.Y(n_4073)
);

AOI22xp33_ASAP7_75t_L g4074 ( 
.A1(n_3784),
.A2(n_561),
.B1(n_558),
.B2(n_560),
.Y(n_4074)
);

AOI22xp33_ASAP7_75t_SL g4075 ( 
.A1(n_3882),
.A2(n_563),
.B1(n_560),
.B2(n_561),
.Y(n_4075)
);

OAI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_3893),
.A2(n_563),
.B(n_564),
.Y(n_4076)
);

AOI22xp33_ASAP7_75t_L g4077 ( 
.A1(n_3815),
.A2(n_566),
.B1(n_564),
.B2(n_565),
.Y(n_4077)
);

OAI21xp5_ASAP7_75t_SL g4078 ( 
.A1(n_3800),
.A2(n_565),
.B(n_566),
.Y(n_4078)
);

AOI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_3761),
.A2(n_572),
.B1(n_568),
.B2(n_571),
.Y(n_4079)
);

OAI222xp33_ASAP7_75t_L g4080 ( 
.A1(n_3845),
.A2(n_568),
.B1(n_571),
.B2(n_573),
.C1(n_574),
.C2(n_575),
.Y(n_4080)
);

AOI22xp33_ASAP7_75t_SL g4081 ( 
.A1(n_3882),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3908),
.B(n_576),
.Y(n_4082)
);

AND2x2_ASAP7_75t_L g4083 ( 
.A(n_3803),
.B(n_806),
.Y(n_4083)
);

AOI22xp33_ASAP7_75t_L g4084 ( 
.A1(n_3719),
.A2(n_579),
.B1(n_577),
.B2(n_578),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3911),
.B(n_577),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3825),
.B(n_578),
.Y(n_4086)
);

AOI22xp33_ASAP7_75t_L g4087 ( 
.A1(n_3851),
.A2(n_3714),
.B1(n_3835),
.B2(n_3831),
.Y(n_4087)
);

AOI22xp33_ASAP7_75t_L g4088 ( 
.A1(n_3906),
.A2(n_582),
.B1(n_580),
.B2(n_581),
.Y(n_4088)
);

AOI22xp33_ASAP7_75t_L g4089 ( 
.A1(n_3917),
.A2(n_582),
.B1(n_580),
.B2(n_581),
.Y(n_4089)
);

OAI22xp5_ASAP7_75t_L g4090 ( 
.A1(n_3776),
.A2(n_585),
.B1(n_583),
.B2(n_584),
.Y(n_4090)
);

AOI22xp33_ASAP7_75t_L g4091 ( 
.A1(n_3925),
.A2(n_585),
.B1(n_583),
.B2(n_584),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_3827),
.B(n_586),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3830),
.B(n_3839),
.Y(n_4093)
);

AOI22xp33_ASAP7_75t_L g4094 ( 
.A1(n_3745),
.A2(n_3691),
.B1(n_3748),
.B2(n_3727),
.Y(n_4094)
);

OAI22xp33_ASAP7_75t_L g4095 ( 
.A1(n_3687),
.A2(n_589),
.B1(n_586),
.B2(n_587),
.Y(n_4095)
);

AOI22xp33_ASAP7_75t_L g4096 ( 
.A1(n_3718),
.A2(n_591),
.B1(n_587),
.B2(n_590),
.Y(n_4096)
);

AOI22xp5_ASAP7_75t_L g4097 ( 
.A1(n_3795),
.A2(n_592),
.B1(n_590),
.B2(n_591),
.Y(n_4097)
);

OAI22xp5_ASAP7_75t_L g4098 ( 
.A1(n_3751),
.A2(n_595),
.B1(n_592),
.B2(n_593),
.Y(n_4098)
);

AOI22xp33_ASAP7_75t_L g4099 ( 
.A1(n_3889),
.A2(n_3675),
.B1(n_3692),
.B2(n_3883),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3874),
.B(n_593),
.Y(n_4100)
);

OAI22xp5_ASAP7_75t_L g4101 ( 
.A1(n_3670),
.A2(n_3720),
.B1(n_3887),
.B2(n_3795),
.Y(n_4101)
);

NAND3xp33_ASAP7_75t_L g4102 ( 
.A(n_3739),
.B(n_596),
.C(n_597),
.Y(n_4102)
);

AOI22xp33_ASAP7_75t_L g4103 ( 
.A1(n_3889),
.A2(n_598),
.B1(n_596),
.B2(n_597),
.Y(n_4103)
);

AOI22xp33_ASAP7_75t_L g4104 ( 
.A1(n_3675),
.A2(n_600),
.B1(n_598),
.B2(n_599),
.Y(n_4104)
);

OAI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_3674),
.A2(n_602),
.B1(n_600),
.B2(n_601),
.Y(n_4105)
);

AOI22xp33_ASAP7_75t_L g4106 ( 
.A1(n_3692),
.A2(n_603),
.B1(n_601),
.B2(n_602),
.Y(n_4106)
);

OAI22xp5_ASAP7_75t_L g4107 ( 
.A1(n_3758),
.A2(n_607),
.B1(n_604),
.B2(n_605),
.Y(n_4107)
);

AOI22xp33_ASAP7_75t_SL g4108 ( 
.A1(n_3883),
.A2(n_608),
.B1(n_605),
.B2(n_607),
.Y(n_4108)
);

OAI22xp33_ASAP7_75t_L g4109 ( 
.A1(n_3687),
.A2(n_611),
.B1(n_608),
.B2(n_609),
.Y(n_4109)
);

AOI22xp33_ASAP7_75t_SL g4110 ( 
.A1(n_3753),
.A2(n_612),
.B1(n_609),
.B2(n_611),
.Y(n_4110)
);

OAI221xp5_ASAP7_75t_L g4111 ( 
.A1(n_3739),
.A2(n_613),
.B1(n_614),
.B2(n_615),
.C(n_616),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3728),
.B(n_613),
.Y(n_4112)
);

OAI22xp5_ASAP7_75t_L g4113 ( 
.A1(n_3672),
.A2(n_618),
.B1(n_614),
.B2(n_617),
.Y(n_4113)
);

AOI22xp5_ASAP7_75t_L g4114 ( 
.A1(n_3913),
.A2(n_620),
.B1(n_617),
.B2(n_619),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_3747),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_3759),
.B(n_621),
.Y(n_4116)
);

AOI22xp5_ASAP7_75t_L g4117 ( 
.A1(n_3850),
.A2(n_625),
.B1(n_622),
.B2(n_623),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_3664),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3763),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_3920),
.Y(n_4120)
);

AOI22xp33_ASAP7_75t_L g4121 ( 
.A1(n_3921),
.A2(n_625),
.B1(n_622),
.B2(n_623),
.Y(n_4121)
);

AND2x2_ASAP7_75t_L g4122 ( 
.A(n_3963),
.B(n_3930),
.Y(n_4122)
);

AOI22xp33_ASAP7_75t_L g4123 ( 
.A1(n_3943),
.A2(n_3838),
.B1(n_3735),
.B2(n_3753),
.Y(n_4123)
);

NAND3xp33_ASAP7_75t_L g4124 ( 
.A(n_3943),
.B(n_3733),
.C(n_3721),
.Y(n_4124)
);

NAND3xp33_ASAP7_75t_L g4125 ( 
.A(n_3945),
.B(n_3916),
.C(n_3912),
.Y(n_4125)
);

OAI22xp5_ASAP7_75t_L g4126 ( 
.A1(n_3945),
.A2(n_3743),
.B1(n_3740),
.B2(n_3841),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_3978),
.B(n_3924),
.Y(n_4127)
);

OAI22xp5_ASAP7_75t_L g4128 ( 
.A1(n_3931),
.A2(n_3673),
.B1(n_3832),
.B2(n_3820),
.Y(n_4128)
);

NOR3xp33_ASAP7_75t_L g4129 ( 
.A(n_3999),
.B(n_3809),
.C(n_3848),
.Y(n_4129)
);

OAI221xp5_ASAP7_75t_L g4130 ( 
.A1(n_4013),
.A2(n_3805),
.B1(n_3904),
.B2(n_3881),
.C(n_3792),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_4043),
.B(n_3919),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_4061),
.B(n_3710),
.Y(n_4132)
);

AND2x2_ASAP7_75t_L g4133 ( 
.A(n_3939),
.B(n_3716),
.Y(n_4133)
);

OAI221xp5_ASAP7_75t_SL g4134 ( 
.A1(n_4038),
.A2(n_3847),
.B1(n_3923),
.B2(n_3926),
.C(n_3788),
.Y(n_4134)
);

OAI221xp5_ASAP7_75t_L g4135 ( 
.A1(n_3935),
.A2(n_3731),
.B1(n_3864),
.B2(n_3848),
.C(n_3789),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3931),
.B(n_3725),
.Y(n_4136)
);

NAND3xp33_ASAP7_75t_L g4137 ( 
.A(n_3969),
.B(n_3779),
.C(n_3828),
.Y(n_4137)
);

AND2x2_ASAP7_75t_L g4138 ( 
.A(n_4031),
.B(n_3836),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_4065),
.B(n_3837),
.Y(n_4139)
);

AOI22xp33_ASAP7_75t_L g4140 ( 
.A1(n_4111),
.A2(n_3829),
.B1(n_3752),
.B2(n_3797),
.Y(n_4140)
);

AND2x2_ASAP7_75t_SL g4141 ( 
.A(n_3958),
.B(n_3864),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_4067),
.B(n_3869),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_4068),
.B(n_3870),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_SL g4144 ( 
.A(n_3953),
.B(n_3829),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_4115),
.B(n_3770),
.Y(n_4145)
);

OAI221xp5_ASAP7_75t_SL g4146 ( 
.A1(n_3959),
.A2(n_3679),
.B1(n_3734),
.B2(n_3823),
.C(n_3822),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_4119),
.B(n_4120),
.Y(n_4147)
);

OAI21xp33_ASAP7_75t_L g4148 ( 
.A1(n_3969),
.A2(n_4078),
.B(n_3934),
.Y(n_4148)
);

NAND2xp33_ASAP7_75t_SL g4149 ( 
.A(n_3941),
.B(n_3857),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_4093),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_3988),
.B(n_3741),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_4002),
.B(n_3771),
.Y(n_4152)
);

OA21x2_ASAP7_75t_L g4153 ( 
.A1(n_3954),
.A2(n_3744),
.B(n_3785),
.Y(n_4153)
);

NAND3xp33_ASAP7_75t_L g4154 ( 
.A(n_4087),
.B(n_3829),
.C(n_3810),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_4057),
.B(n_3811),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_4118),
.B(n_3766),
.Y(n_4156)
);

AND2x2_ASAP7_75t_L g4157 ( 
.A(n_3942),
.B(n_3824),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_4012),
.B(n_3769),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_3933),
.B(n_3843),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_3979),
.B(n_3806),
.Y(n_4160)
);

NAND4xp25_ASAP7_75t_L g4161 ( 
.A(n_4035),
.B(n_3736),
.C(n_3791),
.D(n_3774),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_4005),
.B(n_3806),
.Y(n_4162)
);

NOR3xp33_ASAP7_75t_L g4163 ( 
.A(n_3999),
.B(n_3738),
.C(n_3732),
.Y(n_4163)
);

AOI22xp33_ASAP7_75t_SL g4164 ( 
.A1(n_4011),
.A2(n_3723),
.B1(n_3797),
.B2(n_3760),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_3949),
.B(n_3807),
.Y(n_4165)
);

OAI21xp33_ASAP7_75t_L g4166 ( 
.A1(n_4032),
.A2(n_3783),
.B(n_3780),
.Y(n_4166)
);

AND2x2_ASAP7_75t_L g4167 ( 
.A(n_3956),
.B(n_3808),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_L g4168 ( 
.A(n_3955),
.B(n_3813),
.Y(n_4168)
);

AOI22xp5_ASAP7_75t_L g4169 ( 
.A1(n_3967),
.A2(n_3910),
.B1(n_3756),
.B2(n_3750),
.Y(n_4169)
);

AND2x2_ASAP7_75t_L g4170 ( 
.A(n_3962),
.B(n_3655),
.Y(n_4170)
);

AND2x2_ASAP7_75t_L g4171 ( 
.A(n_3950),
.B(n_3655),
.Y(n_4171)
);

AND2x2_ASAP7_75t_L g4172 ( 
.A(n_3998),
.B(n_3817),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_4049),
.B(n_4051),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_3998),
.B(n_3817),
.Y(n_4174)
);

AND2x2_ASAP7_75t_L g4175 ( 
.A(n_4094),
.B(n_3846),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_4073),
.Y(n_4176)
);

OAI22xp5_ASAP7_75t_L g4177 ( 
.A1(n_4102),
.A2(n_3834),
.B1(n_3846),
.B2(n_3786),
.Y(n_4177)
);

AND2x2_ASAP7_75t_L g4178 ( 
.A(n_4083),
.B(n_3844),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4018),
.B(n_3818),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_SL g4180 ( 
.A(n_3936),
.B(n_3833),
.Y(n_4180)
);

AND2x2_ASAP7_75t_L g4181 ( 
.A(n_4099),
.B(n_3856),
.Y(n_4181)
);

AND2x2_ASAP7_75t_L g4182 ( 
.A(n_3960),
.B(n_3856),
.Y(n_4182)
);

AND2x2_ASAP7_75t_L g4183 ( 
.A(n_3948),
.B(n_3856),
.Y(n_4183)
);

AND2x2_ASAP7_75t_L g4184 ( 
.A(n_3951),
.B(n_3903),
.Y(n_4184)
);

NOR3xp33_ASAP7_75t_L g4185 ( 
.A(n_3987),
.B(n_3746),
.C(n_3749),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_4006),
.B(n_627),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_4018),
.B(n_3903),
.Y(n_4187)
);

OAI221xp5_ASAP7_75t_L g4188 ( 
.A1(n_4024),
.A2(n_3910),
.B1(n_3927),
.B2(n_3767),
.C(n_3802),
.Y(n_4188)
);

OAI22xp5_ASAP7_75t_L g4189 ( 
.A1(n_4045),
.A2(n_3712),
.B1(n_3694),
.B2(n_3757),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_4018),
.B(n_3903),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4009),
.Y(n_4191)
);

NAND3xp33_ASAP7_75t_L g4192 ( 
.A(n_3990),
.B(n_3778),
.C(n_3875),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4019),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_L g4194 ( 
.A(n_4037),
.B(n_4040),
.Y(n_4194)
);

OAI22xp5_ASAP7_75t_L g4195 ( 
.A1(n_4029),
.A2(n_3928),
.B1(n_3884),
.B2(n_630),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_3932),
.B(n_628),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_4023),
.B(n_628),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_SL g4198 ( 
.A(n_3961),
.B(n_629),
.Y(n_4198)
);

NOR3xp33_ASAP7_75t_L g4199 ( 
.A(n_4056),
.B(n_629),
.C(n_631),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_4046),
.B(n_632),
.Y(n_4200)
);

NOR2xp33_ASAP7_75t_L g4201 ( 
.A(n_3957),
.B(n_632),
.Y(n_4201)
);

AND2x2_ASAP7_75t_L g4202 ( 
.A(n_4041),
.B(n_4086),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_L g4203 ( 
.A(n_4092),
.B(n_633),
.Y(n_4203)
);

NAND4xp25_ASAP7_75t_L g4204 ( 
.A(n_4032),
.B(n_633),
.C(n_634),
.D(n_635),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_4100),
.B(n_634),
.Y(n_4205)
);

NOR3xp33_ASAP7_75t_L g4206 ( 
.A(n_4017),
.B(n_636),
.C(n_637),
.Y(n_4206)
);

NAND3xp33_ASAP7_75t_L g4207 ( 
.A(n_3984),
.B(n_636),
.C(n_637),
.Y(n_4207)
);

NOR3xp33_ASAP7_75t_L g4208 ( 
.A(n_4015),
.B(n_639),
.C(n_640),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_4112),
.B(n_804),
.Y(n_4209)
);

AND2x2_ASAP7_75t_L g4210 ( 
.A(n_4116),
.B(n_639),
.Y(n_4210)
);

OAI21xp33_ASAP7_75t_L g4211 ( 
.A1(n_4033),
.A2(n_640),
.B(n_641),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_4082),
.B(n_642),
.Y(n_4212)
);

INVx1_ASAP7_75t_SL g4213 ( 
.A(n_4200),
.Y(n_4213)
);

AOI22xp33_ASAP7_75t_L g4214 ( 
.A1(n_4129),
.A2(n_4071),
.B1(n_4090),
.B2(n_4076),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_4122),
.B(n_3964),
.Y(n_4215)
);

AO21x2_ASAP7_75t_L g4216 ( 
.A1(n_4179),
.A2(n_4022),
.B(n_4085),
.Y(n_4216)
);

CKINVDCx20_ASAP7_75t_R g4217 ( 
.A(n_4149),
.Y(n_4217)
);

BUFx3_ASAP7_75t_L g4218 ( 
.A(n_4172),
.Y(n_4218)
);

NOR2xp33_ASAP7_75t_L g4219 ( 
.A(n_4135),
.B(n_3946),
.Y(n_4219)
);

NOR3xp33_ASAP7_75t_L g4220 ( 
.A(n_4195),
.B(n_4080),
.C(n_4059),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4147),
.Y(n_4221)
);

NOR2x1_ASAP7_75t_L g4222 ( 
.A(n_4180),
.B(n_3992),
.Y(n_4222)
);

NOR3xp33_ASAP7_75t_L g4223 ( 
.A(n_4195),
.B(n_4109),
.C(n_4095),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_4133),
.B(n_3940),
.Y(n_4224)
);

NOR3xp33_ASAP7_75t_L g4225 ( 
.A(n_4189),
.B(n_4109),
.C(n_4095),
.Y(n_4225)
);

AOI22xp33_ASAP7_75t_L g4226 ( 
.A1(n_4148),
.A2(n_3986),
.B1(n_4058),
.B2(n_4066),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_4127),
.Y(n_4227)
);

NAND3xp33_ASAP7_75t_L g4228 ( 
.A(n_4164),
.B(n_3995),
.C(n_4029),
.Y(n_4228)
);

NOR3xp33_ASAP7_75t_L g4229 ( 
.A(n_4189),
.B(n_4069),
.C(n_3937),
.Y(n_4229)
);

INVx2_ASAP7_75t_SL g4230 ( 
.A(n_4174),
.Y(n_4230)
);

HB1xp67_ASAP7_75t_L g4231 ( 
.A(n_4157),
.Y(n_4231)
);

OAI211xp5_ASAP7_75t_SL g4232 ( 
.A1(n_4188),
.A2(n_4033),
.B(n_4007),
.C(n_4020),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_4150),
.B(n_3938),
.Y(n_4233)
);

NOR2xp33_ASAP7_75t_L g4234 ( 
.A(n_4192),
.B(n_4101),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_4158),
.B(n_3947),
.Y(n_4235)
);

AOI221xp5_ASAP7_75t_L g4236 ( 
.A1(n_4126),
.A2(n_4042),
.B1(n_3989),
.B2(n_4053),
.C(n_4039),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_4162),
.B(n_3952),
.Y(n_4237)
);

NAND4xp75_ASAP7_75t_L g4238 ( 
.A(n_4141),
.B(n_4070),
.C(n_4114),
.D(n_4026),
.Y(n_4238)
);

AOI22xp5_ASAP7_75t_L g4239 ( 
.A1(n_4185),
.A2(n_3997),
.B1(n_4030),
.B2(n_4042),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_4138),
.Y(n_4240)
);

OR2x2_ASAP7_75t_L g4241 ( 
.A(n_4127),
.B(n_4030),
.Y(n_4241)
);

NAND4xp75_ASAP7_75t_L g4242 ( 
.A(n_4175),
.B(n_4097),
.C(n_4117),
.D(n_4016),
.Y(n_4242)
);

NOR3xp33_ASAP7_75t_SL g4243 ( 
.A(n_4146),
.B(n_3973),
.C(n_4004),
.Y(n_4243)
);

NAND3xp33_ASAP7_75t_L g4244 ( 
.A(n_4163),
.B(n_4110),
.C(n_4063),
.Y(n_4244)
);

NAND3xp33_ASAP7_75t_L g4245 ( 
.A(n_4126),
.B(n_4034),
.C(n_4075),
.Y(n_4245)
);

NOR3xp33_ASAP7_75t_L g4246 ( 
.A(n_4161),
.B(n_3976),
.C(n_4003),
.Y(n_4246)
);

OR2x2_ASAP7_75t_L g4247 ( 
.A(n_4131),
.B(n_4121),
.Y(n_4247)
);

AOI22xp33_ASAP7_75t_L g4248 ( 
.A1(n_4199),
.A2(n_3966),
.B1(n_4098),
.B2(n_3972),
.Y(n_4248)
);

NAND3xp33_ASAP7_75t_L g4249 ( 
.A(n_4177),
.B(n_4108),
.C(n_4081),
.Y(n_4249)
);

NOR2xp33_ASAP7_75t_L g4250 ( 
.A(n_4191),
.B(n_3944),
.Y(n_4250)
);

OR2x2_ASAP7_75t_L g4251 ( 
.A(n_4131),
.B(n_4121),
.Y(n_4251)
);

OA211x2_ASAP7_75t_L g4252 ( 
.A1(n_4166),
.A2(n_4014),
.B(n_4021),
.C(n_4084),
.Y(n_4252)
);

OR2x2_ASAP7_75t_L g4253 ( 
.A(n_4156),
.B(n_4054),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4132),
.Y(n_4254)
);

NOR2xp33_ASAP7_75t_SL g4255 ( 
.A(n_4124),
.B(n_4107),
.Y(n_4255)
);

AND2x2_ASAP7_75t_L g4256 ( 
.A(n_4170),
.B(n_3965),
.Y(n_4256)
);

NAND4xp75_ASAP7_75t_L g4257 ( 
.A(n_4144),
.B(n_4036),
.C(n_3970),
.D(n_4010),
.Y(n_4257)
);

AND2x2_ASAP7_75t_L g4258 ( 
.A(n_4178),
.B(n_4096),
.Y(n_4258)
);

NOR3xp33_ASAP7_75t_L g4259 ( 
.A(n_4177),
.B(n_4128),
.C(n_4130),
.Y(n_4259)
);

AND2x2_ASAP7_75t_L g4260 ( 
.A(n_4145),
.B(n_4079),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4132),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4139),
.Y(n_4262)
);

OR2x2_ASAP7_75t_L g4263 ( 
.A(n_4156),
.B(n_4027),
.Y(n_4263)
);

OA211x2_ASAP7_75t_L g4264 ( 
.A1(n_4198),
.A2(n_3968),
.B(n_4048),
.C(n_3983),
.Y(n_4264)
);

INVx2_ASAP7_75t_SL g4265 ( 
.A(n_4160),
.Y(n_4265)
);

AO21x2_ASAP7_75t_L g4266 ( 
.A1(n_4179),
.A2(n_4196),
.B(n_4136),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4193),
.B(n_3994),
.Y(n_4267)
);

AOI22xp5_ASAP7_75t_L g4268 ( 
.A1(n_4204),
.A2(n_4105),
.B1(n_3996),
.B2(n_4113),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4142),
.Y(n_4269)
);

NOR3xp33_ASAP7_75t_L g4270 ( 
.A(n_4128),
.B(n_3982),
.C(n_4088),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_4152),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_4176),
.B(n_4044),
.Y(n_4272)
);

INVx2_ASAP7_75t_SL g4273 ( 
.A(n_4155),
.Y(n_4273)
);

AND2x2_ASAP7_75t_L g4274 ( 
.A(n_4181),
.B(n_3975),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4143),
.Y(n_4275)
);

AND2x2_ASAP7_75t_L g4276 ( 
.A(n_4183),
.B(n_4055),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4151),
.Y(n_4277)
);

AND2x2_ASAP7_75t_L g4278 ( 
.A(n_4182),
.B(n_4064),
.Y(n_4278)
);

NOR3xp33_ASAP7_75t_L g4279 ( 
.A(n_4201),
.B(n_4091),
.C(n_4089),
.Y(n_4279)
);

AND2x2_ASAP7_75t_L g4280 ( 
.A(n_4167),
.B(n_4072),
.Y(n_4280)
);

NOR4xp25_ASAP7_75t_L g4281 ( 
.A(n_4134),
.B(n_3993),
.C(n_4000),
.D(n_3980),
.Y(n_4281)
);

NAND4xp75_ASAP7_75t_L g4282 ( 
.A(n_4171),
.B(n_4074),
.C(n_4077),
.D(n_4008),
.Y(n_4282)
);

INVx3_ASAP7_75t_L g4283 ( 
.A(n_4218),
.Y(n_4283)
);

NOR3xp33_ASAP7_75t_SL g4284 ( 
.A(n_4245),
.B(n_4154),
.C(n_4125),
.Y(n_4284)
);

NOR3xp33_ASAP7_75t_L g4285 ( 
.A(n_4259),
.B(n_4211),
.C(n_4208),
.Y(n_4285)
);

XNOR2xp5_ASAP7_75t_L g4286 ( 
.A(n_4217),
.B(n_4202),
.Y(n_4286)
);

NAND4xp75_ASAP7_75t_L g4287 ( 
.A(n_4222),
.B(n_4197),
.C(n_4169),
.D(n_4184),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_4254),
.Y(n_4288)
);

AND2x2_ASAP7_75t_L g4289 ( 
.A(n_4230),
.B(n_4187),
.Y(n_4289)
);

NAND4xp75_ASAP7_75t_L g4290 ( 
.A(n_4252),
.B(n_4190),
.C(n_4194),
.D(n_4210),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4261),
.Y(n_4291)
);

XNOR2x2_ASAP7_75t_L g4292 ( 
.A(n_4234),
.B(n_4137),
.Y(n_4292)
);

AND2x2_ASAP7_75t_L g4293 ( 
.A(n_4231),
.B(n_4153),
.Y(n_4293)
);

XOR2x2_ASAP7_75t_L g4294 ( 
.A(n_4229),
.B(n_4207),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4271),
.Y(n_4295)
);

BUFx2_ASAP7_75t_SL g4296 ( 
.A(n_4213),
.Y(n_4296)
);

CKINVDCx5p33_ASAP7_75t_R g4297 ( 
.A(n_4250),
.Y(n_4297)
);

NAND4xp75_ASAP7_75t_SL g4298 ( 
.A(n_4219),
.B(n_4153),
.C(n_4140),
.D(n_4123),
.Y(n_4298)
);

NAND4xp75_ASAP7_75t_L g4299 ( 
.A(n_4264),
.B(n_4168),
.C(n_4173),
.D(n_4159),
.Y(n_4299)
);

INVx3_ASAP7_75t_L g4300 ( 
.A(n_4240),
.Y(n_4300)
);

XOR2x1_ASAP7_75t_L g4301 ( 
.A(n_4235),
.B(n_4206),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_4266),
.B(n_4173),
.Y(n_4302)
);

INVx2_ASAP7_75t_SL g4303 ( 
.A(n_4273),
.Y(n_4303)
);

XNOR2x1_ASAP7_75t_L g4304 ( 
.A(n_4282),
.B(n_4186),
.Y(n_4304)
);

XNOR2xp5_ASAP7_75t_L g4305 ( 
.A(n_4215),
.B(n_4203),
.Y(n_4305)
);

CKINVDCx5p33_ASAP7_75t_R g4306 ( 
.A(n_4265),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4227),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4262),
.Y(n_4308)
);

NAND4xp75_ASAP7_75t_L g4309 ( 
.A(n_4239),
.B(n_4243),
.C(n_4236),
.D(n_4278),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4269),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4275),
.Y(n_4311)
);

OR2x2_ASAP7_75t_L g4312 ( 
.A(n_4277),
.B(n_4165),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_4266),
.B(n_4212),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_4224),
.B(n_4212),
.Y(n_4314)
);

XNOR2xp5_ASAP7_75t_L g4315 ( 
.A(n_4237),
.B(n_4205),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4221),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4233),
.Y(n_4317)
);

AOI22xp5_ASAP7_75t_L g4318 ( 
.A1(n_4225),
.A2(n_4209),
.B1(n_4047),
.B2(n_4028),
.Y(n_4318)
);

XNOR2xp5_ASAP7_75t_L g4319 ( 
.A(n_4245),
.B(n_3991),
.Y(n_4319)
);

NAND4xp75_ASAP7_75t_SL g4320 ( 
.A(n_4280),
.B(n_3974),
.C(n_3971),
.D(n_4028),
.Y(n_4320)
);

NAND4xp75_ASAP7_75t_SL g4321 ( 
.A(n_4276),
.B(n_4274),
.C(n_4220),
.D(n_4249),
.Y(n_4321)
);

OAI22x1_ASAP7_75t_L g4322 ( 
.A1(n_4244),
.A2(n_4106),
.B1(n_4104),
.B2(n_4103),
.Y(n_4322)
);

INVx2_ASAP7_75t_SL g4323 ( 
.A(n_4256),
.Y(n_4323)
);

INVx4_ASAP7_75t_L g4324 ( 
.A(n_4216),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_4241),
.B(n_4247),
.Y(n_4325)
);

NAND4xp75_ASAP7_75t_L g4326 ( 
.A(n_4239),
.B(n_3985),
.C(n_3981),
.D(n_3977),
.Y(n_4326)
);

BUFx2_ASAP7_75t_L g4327 ( 
.A(n_4216),
.Y(n_4327)
);

INVx2_ASAP7_75t_SL g4328 ( 
.A(n_4258),
.Y(n_4328)
);

NAND4xp75_ASAP7_75t_L g4329 ( 
.A(n_4267),
.B(n_4001),
.C(n_4060),
.D(n_4052),
.Y(n_4329)
);

AOI22xp5_ASAP7_75t_L g4330 ( 
.A1(n_4255),
.A2(n_4050),
.B1(n_4062),
.B2(n_4025),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4251),
.Y(n_4331)
);

NOR3xp33_ASAP7_75t_L g4332 ( 
.A(n_4249),
.B(n_642),
.C(n_643),
.Y(n_4332)
);

OR2x2_ASAP7_75t_L g4333 ( 
.A(n_4263),
.B(n_644),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_4253),
.B(n_644),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4272),
.Y(n_4335)
);

INVx4_ASAP7_75t_L g4336 ( 
.A(n_4260),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_4226),
.B(n_646),
.Y(n_4337)
);

NOR3xp33_ASAP7_75t_L g4338 ( 
.A(n_4244),
.B(n_647),
.C(n_648),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4223),
.Y(n_4339)
);

INVx2_ASAP7_75t_L g4340 ( 
.A(n_4242),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_4270),
.B(n_647),
.Y(n_4341)
);

BUFx2_ASAP7_75t_L g4342 ( 
.A(n_4228),
.Y(n_4342)
);

BUFx2_ASAP7_75t_L g4343 ( 
.A(n_4228),
.Y(n_4343)
);

NAND4xp75_ASAP7_75t_L g4344 ( 
.A(n_4268),
.B(n_649),
.C(n_650),
.D(n_651),
.Y(n_4344)
);

OR2x2_ASAP7_75t_L g4345 ( 
.A(n_4331),
.B(n_4281),
.Y(n_4345)
);

AOI22xp5_ASAP7_75t_L g4346 ( 
.A1(n_4309),
.A2(n_4246),
.B1(n_4214),
.B2(n_4238),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4300),
.Y(n_4347)
);

INVxp67_ASAP7_75t_L g4348 ( 
.A(n_4296),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4295),
.Y(n_4349)
);

AND2x2_ASAP7_75t_L g4350 ( 
.A(n_4283),
.B(n_4281),
.Y(n_4350)
);

INVx1_ASAP7_75t_SL g4351 ( 
.A(n_4283),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_4331),
.B(n_4279),
.Y(n_4352)
);

HB1xp67_ASAP7_75t_L g4353 ( 
.A(n_4300),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4295),
.Y(n_4354)
);

NOR2xp33_ASAP7_75t_L g4355 ( 
.A(n_4342),
.B(n_4232),
.Y(n_4355)
);

XOR2x2_ASAP7_75t_L g4356 ( 
.A(n_4321),
.B(n_4257),
.Y(n_4356)
);

INVx4_ASAP7_75t_L g4357 ( 
.A(n_4306),
.Y(n_4357)
);

XNOR2x1_ASAP7_75t_L g4358 ( 
.A(n_4299),
.B(n_4268),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4291),
.Y(n_4359)
);

INVx2_ASAP7_75t_L g4360 ( 
.A(n_4288),
.Y(n_4360)
);

INVxp67_ASAP7_75t_L g4361 ( 
.A(n_4340),
.Y(n_4361)
);

XNOR2x1_ASAP7_75t_L g4362 ( 
.A(n_4290),
.B(n_650),
.Y(n_4362)
);

XOR2x2_ASAP7_75t_L g4363 ( 
.A(n_4286),
.B(n_4304),
.Y(n_4363)
);

AO22x1_ASAP7_75t_L g4364 ( 
.A1(n_4343),
.A2(n_4248),
.B1(n_653),
.B2(n_654),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4307),
.Y(n_4365)
);

CKINVDCx16_ASAP7_75t_R g4366 ( 
.A(n_4333),
.Y(n_4366)
);

XNOR2xp5_ASAP7_75t_L g4367 ( 
.A(n_4301),
.B(n_652),
.Y(n_4367)
);

INVx1_ASAP7_75t_SL g4368 ( 
.A(n_4303),
.Y(n_4368)
);

XOR2x2_ASAP7_75t_L g4369 ( 
.A(n_4292),
.B(n_652),
.Y(n_4369)
);

INVx2_ASAP7_75t_L g4370 ( 
.A(n_4308),
.Y(n_4370)
);

AO22x2_ASAP7_75t_L g4371 ( 
.A1(n_4339),
.A2(n_654),
.B1(n_656),
.B2(n_657),
.Y(n_4371)
);

XOR2x2_ASAP7_75t_L g4372 ( 
.A(n_4294),
.B(n_656),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4316),
.Y(n_4373)
);

INVx2_ASAP7_75t_L g4374 ( 
.A(n_4310),
.Y(n_4374)
);

AND2x2_ASAP7_75t_L g4375 ( 
.A(n_4323),
.B(n_658),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_4328),
.B(n_659),
.Y(n_4376)
);

XOR2x2_ASAP7_75t_L g4377 ( 
.A(n_4305),
.B(n_660),
.Y(n_4377)
);

XNOR2xp5_ASAP7_75t_L g4378 ( 
.A(n_4287),
.B(n_660),
.Y(n_4378)
);

AND2x2_ASAP7_75t_L g4379 ( 
.A(n_4336),
.B(n_661),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_4336),
.B(n_661),
.Y(n_4380)
);

XOR2x2_ASAP7_75t_L g4381 ( 
.A(n_4315),
.B(n_662),
.Y(n_4381)
);

OA22x2_ASAP7_75t_L g4382 ( 
.A1(n_4297),
.A2(n_662),
.B1(n_663),
.B2(n_664),
.Y(n_4382)
);

INVx4_ASAP7_75t_L g4383 ( 
.A(n_4324),
.Y(n_4383)
);

AOI22xp5_ASAP7_75t_L g4384 ( 
.A1(n_4319),
.A2(n_663),
.B1(n_665),
.B2(n_666),
.Y(n_4384)
);

INVx2_ASAP7_75t_SL g4385 ( 
.A(n_4289),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4370),
.Y(n_4386)
);

BUFx3_ASAP7_75t_L g4387 ( 
.A(n_4357),
.Y(n_4387)
);

OAI22xp33_ASAP7_75t_SL g4388 ( 
.A1(n_4345),
.A2(n_4324),
.B1(n_4313),
.B2(n_4302),
.Y(n_4388)
);

INVx2_ASAP7_75t_SL g4389 ( 
.A(n_4357),
.Y(n_4389)
);

XNOR2xp5_ASAP7_75t_L g4390 ( 
.A(n_4363),
.B(n_4298),
.Y(n_4390)
);

XOR2x2_ASAP7_75t_L g4391 ( 
.A(n_4356),
.B(n_4320),
.Y(n_4391)
);

AOI22x1_ASAP7_75t_SL g4392 ( 
.A1(n_4383),
.A2(n_4317),
.B1(n_4284),
.B2(n_4335),
.Y(n_4392)
);

XOR2x2_ASAP7_75t_L g4393 ( 
.A(n_4372),
.B(n_4369),
.Y(n_4393)
);

OAI22xp5_ASAP7_75t_L g4394 ( 
.A1(n_4361),
.A2(n_4325),
.B1(n_4312),
.B2(n_4293),
.Y(n_4394)
);

AOI22xp5_ASAP7_75t_L g4395 ( 
.A1(n_4346),
.A2(n_4285),
.B1(n_4332),
.B2(n_4338),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4374),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4373),
.Y(n_4397)
);

OA22x2_ASAP7_75t_L g4398 ( 
.A1(n_4350),
.A2(n_4341),
.B1(n_4327),
.B2(n_4318),
.Y(n_4398)
);

AOI22xp5_ASAP7_75t_L g4399 ( 
.A1(n_4358),
.A2(n_4329),
.B1(n_4326),
.B2(n_4337),
.Y(n_4399)
);

INVx3_ASAP7_75t_L g4400 ( 
.A(n_4351),
.Y(n_4400)
);

INVx2_ASAP7_75t_L g4401 ( 
.A(n_4353),
.Y(n_4401)
);

BUFx2_ASAP7_75t_L g4402 ( 
.A(n_4383),
.Y(n_4402)
);

NAND2x1_ASAP7_75t_L g4403 ( 
.A(n_4349),
.B(n_4354),
.Y(n_4403)
);

BUFx2_ASAP7_75t_L g4404 ( 
.A(n_4348),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4373),
.Y(n_4405)
);

INVx2_ASAP7_75t_L g4406 ( 
.A(n_4360),
.Y(n_4406)
);

XNOR2xp5_ASAP7_75t_L g4407 ( 
.A(n_4381),
.B(n_4322),
.Y(n_4407)
);

BUFx3_ASAP7_75t_L g4408 ( 
.A(n_4368),
.Y(n_4408)
);

BUFx2_ASAP7_75t_L g4409 ( 
.A(n_4367),
.Y(n_4409)
);

INVx3_ASAP7_75t_L g4410 ( 
.A(n_4379),
.Y(n_4410)
);

BUFx2_ASAP7_75t_L g4411 ( 
.A(n_4352),
.Y(n_4411)
);

AOI22x1_ASAP7_75t_L g4412 ( 
.A1(n_4378),
.A2(n_4311),
.B1(n_4344),
.B2(n_4334),
.Y(n_4412)
);

OA22x2_ASAP7_75t_L g4413 ( 
.A1(n_4380),
.A2(n_4314),
.B1(n_4330),
.B2(n_669),
.Y(n_4413)
);

OA22x2_ASAP7_75t_L g4414 ( 
.A1(n_4384),
.A2(n_667),
.B1(n_668),
.B2(n_669),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4359),
.Y(n_4415)
);

AO22x2_ASAP7_75t_L g4416 ( 
.A1(n_4362),
.A2(n_667),
.B1(n_668),
.B2(n_670),
.Y(n_4416)
);

XNOR2x1_ASAP7_75t_L g4417 ( 
.A(n_4377),
.B(n_671),
.Y(n_4417)
);

INVx3_ASAP7_75t_SL g4418 ( 
.A(n_4382),
.Y(n_4418)
);

OAI22x1_ASAP7_75t_L g4419 ( 
.A1(n_4355),
.A2(n_671),
.B1(n_672),
.B2(n_674),
.Y(n_4419)
);

AOI22x1_ASAP7_75t_SL g4420 ( 
.A1(n_4364),
.A2(n_4366),
.B1(n_4347),
.B2(n_4365),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_4349),
.Y(n_4421)
);

BUFx6f_ASAP7_75t_L g4422 ( 
.A(n_4375),
.Y(n_4422)
);

OA22x2_ASAP7_75t_L g4423 ( 
.A1(n_4384),
.A2(n_674),
.B1(n_676),
.B2(n_677),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4359),
.Y(n_4424)
);

INVx2_ASAP7_75t_L g4425 ( 
.A(n_4354),
.Y(n_4425)
);

HB1xp67_ASAP7_75t_L g4426 ( 
.A(n_4365),
.Y(n_4426)
);

INVx3_ASAP7_75t_L g4427 ( 
.A(n_4385),
.Y(n_4427)
);

XNOR2x1_ASAP7_75t_L g4428 ( 
.A(n_4371),
.B(n_676),
.Y(n_4428)
);

OAI322xp33_ASAP7_75t_L g4429 ( 
.A1(n_4398),
.A2(n_4366),
.A3(n_4376),
.B1(n_4371),
.B2(n_682),
.C1(n_683),
.C2(n_684),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_4404),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_4404),
.Y(n_4431)
);

HB1xp67_ASAP7_75t_L g4432 ( 
.A(n_4408),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4426),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4402),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4402),
.Y(n_4435)
);

BUFx4f_ASAP7_75t_SL g4436 ( 
.A(n_4387),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_4400),
.Y(n_4437)
);

OAI22xp5_ASAP7_75t_L g4438 ( 
.A1(n_4399),
.A2(n_678),
.B1(n_680),
.B2(n_681),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_4397),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4405),
.Y(n_4440)
);

OAI322xp33_ASAP7_75t_L g4441 ( 
.A1(n_4395),
.A2(n_681),
.A3(n_682),
.B1(n_683),
.B2(n_684),
.C1(n_685),
.C2(n_686),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4415),
.Y(n_4442)
);

INVx2_ASAP7_75t_SL g4443 ( 
.A(n_4389),
.Y(n_4443)
);

XOR2x2_ASAP7_75t_L g4444 ( 
.A(n_4393),
.B(n_685),
.Y(n_4444)
);

INVxp33_ASAP7_75t_SL g4445 ( 
.A(n_4407),
.Y(n_4445)
);

INVx2_ASAP7_75t_L g4446 ( 
.A(n_4401),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4424),
.Y(n_4447)
);

OA22x2_ASAP7_75t_L g4448 ( 
.A1(n_4390),
.A2(n_686),
.B1(n_687),
.B2(n_688),
.Y(n_4448)
);

OAI322xp33_ASAP7_75t_L g4449 ( 
.A1(n_4413),
.A2(n_688),
.A3(n_690),
.B1(n_694),
.B2(n_695),
.C1(n_696),
.C2(n_697),
.Y(n_4449)
);

INVxp67_ASAP7_75t_SL g4450 ( 
.A(n_4428),
.Y(n_4450)
);

CKINVDCx16_ASAP7_75t_R g4451 ( 
.A(n_4409),
.Y(n_4451)
);

INVx2_ASAP7_75t_L g4452 ( 
.A(n_4406),
.Y(n_4452)
);

CKINVDCx5p33_ASAP7_75t_R g4453 ( 
.A(n_4409),
.Y(n_4453)
);

HB1xp67_ASAP7_75t_L g4454 ( 
.A(n_4386),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4396),
.Y(n_4455)
);

INVx2_ASAP7_75t_L g4456 ( 
.A(n_4403),
.Y(n_4456)
);

INVx2_ASAP7_75t_L g4457 ( 
.A(n_4403),
.Y(n_4457)
);

INVx2_ASAP7_75t_SL g4458 ( 
.A(n_4427),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4432),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4432),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4430),
.Y(n_4461)
);

AOI22xp5_ASAP7_75t_L g4462 ( 
.A1(n_4443),
.A2(n_4418),
.B1(n_4392),
.B2(n_4420),
.Y(n_4462)
);

OAI22xp33_ASAP7_75t_L g4463 ( 
.A1(n_4458),
.A2(n_4411),
.B1(n_4394),
.B2(n_4410),
.Y(n_4463)
);

NAND4xp25_ASAP7_75t_L g4464 ( 
.A(n_4445),
.B(n_4411),
.C(n_4391),
.D(n_4392),
.Y(n_4464)
);

AO22x2_ASAP7_75t_L g4465 ( 
.A1(n_4434),
.A2(n_4420),
.B1(n_4417),
.B2(n_4425),
.Y(n_4465)
);

BUFx4_ASAP7_75t_R g4466 ( 
.A(n_4437),
.Y(n_4466)
);

AOI32xp33_ASAP7_75t_L g4467 ( 
.A1(n_4450),
.A2(n_4416),
.A3(n_4388),
.B1(n_4412),
.B2(n_4421),
.Y(n_4467)
);

AOI211xp5_ASAP7_75t_SL g4468 ( 
.A1(n_4429),
.A2(n_4416),
.B(n_4419),
.C(n_4423),
.Y(n_4468)
);

OAI322xp33_ASAP7_75t_L g4469 ( 
.A1(n_4431),
.A2(n_4414),
.A3(n_4422),
.B1(n_696),
.B2(n_698),
.C1(n_699),
.C2(n_700),
.Y(n_4469)
);

AOI211xp5_ASAP7_75t_SL g4470 ( 
.A1(n_4436),
.A2(n_4422),
.B(n_695),
.C(n_698),
.Y(n_4470)
);

AO22x2_ASAP7_75t_L g4471 ( 
.A1(n_4435),
.A2(n_4422),
.B1(n_699),
.B2(n_700),
.Y(n_4471)
);

BUFx6f_ASAP7_75t_L g4472 ( 
.A(n_4453),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4454),
.Y(n_4473)
);

AOI211x1_ASAP7_75t_L g4474 ( 
.A1(n_4433),
.A2(n_694),
.B(n_701),
.C(n_702),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4454),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4446),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4446),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4455),
.Y(n_4478)
);

OAI322xp33_ASAP7_75t_L g4479 ( 
.A1(n_4451),
.A2(n_703),
.A3(n_704),
.B1(n_705),
.B2(n_706),
.C1(n_707),
.C2(n_708),
.Y(n_4479)
);

AOI221xp5_ASAP7_75t_L g4480 ( 
.A1(n_4450),
.A2(n_705),
.B1(n_709),
.B2(n_710),
.C(n_711),
.Y(n_4480)
);

AO22x2_ASAP7_75t_L g4481 ( 
.A1(n_4456),
.A2(n_710),
.B1(n_711),
.B2(n_713),
.Y(n_4481)
);

OAI22x1_ASAP7_75t_L g4482 ( 
.A1(n_4462),
.A2(n_4436),
.B1(n_4456),
.B2(n_4457),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4459),
.Y(n_4483)
);

NOR2x1_ASAP7_75t_L g4484 ( 
.A(n_4464),
.B(n_4449),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_4460),
.Y(n_4485)
);

OAI211xp5_ASAP7_75t_SL g4486 ( 
.A1(n_4467),
.A2(n_4438),
.B(n_4444),
.C(n_4448),
.Y(n_4486)
);

HB1xp67_ASAP7_75t_SL g4487 ( 
.A(n_4472),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4476),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4477),
.Y(n_4489)
);

OAI22xp5_ASAP7_75t_L g4490 ( 
.A1(n_4465),
.A2(n_4452),
.B1(n_4447),
.B2(n_4442),
.Y(n_4490)
);

OAI22xp5_ASAP7_75t_L g4491 ( 
.A1(n_4463),
.A2(n_4461),
.B1(n_4475),
.B2(n_4473),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4471),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4481),
.Y(n_4493)
);

O2A1O1Ixp33_ASAP7_75t_SL g4494 ( 
.A1(n_4468),
.A2(n_4440),
.B(n_4439),
.C(n_4448),
.Y(n_4494)
);

AOI22xp5_ASAP7_75t_L g4495 ( 
.A1(n_4472),
.A2(n_4452),
.B1(n_4441),
.B2(n_716),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_4478),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4466),
.Y(n_4497)
);

OAI22x1_ASAP7_75t_L g4498 ( 
.A1(n_4469),
.A2(n_714),
.B1(n_715),
.B2(n_716),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4479),
.Y(n_4499)
);

O2A1O1Ixp33_ASAP7_75t_SL g4500 ( 
.A1(n_4470),
.A2(n_714),
.B(n_715),
.C(n_717),
.Y(n_4500)
);

O2A1O1Ixp33_ASAP7_75t_SL g4501 ( 
.A1(n_4480),
.A2(n_719),
.B(n_720),
.C(n_721),
.Y(n_4501)
);

NOR2x1_ASAP7_75t_L g4502 ( 
.A(n_4497),
.B(n_4474),
.Y(n_4502)
);

AO22x1_ASAP7_75t_L g4503 ( 
.A1(n_4484),
.A2(n_719),
.B1(n_721),
.B2(n_723),
.Y(n_4503)
);

OAI221xp5_ASAP7_75t_L g4504 ( 
.A1(n_4490),
.A2(n_724),
.B1(n_725),
.B2(n_726),
.C(n_727),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4488),
.Y(n_4505)
);

INVx2_ASAP7_75t_L g4506 ( 
.A(n_4489),
.Y(n_4506)
);

NOR2xp33_ASAP7_75t_L g4507 ( 
.A(n_4487),
.B(n_724),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4483),
.Y(n_4508)
);

NAND4xp25_ASAP7_75t_SL g4509 ( 
.A(n_4499),
.B(n_725),
.C(n_726),
.D(n_727),
.Y(n_4509)
);

AO22x2_ASAP7_75t_L g4510 ( 
.A1(n_4492),
.A2(n_728),
.B1(n_729),
.B2(n_730),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4485),
.Y(n_4511)
);

AO22x1_ASAP7_75t_L g4512 ( 
.A1(n_4493),
.A2(n_4491),
.B1(n_4496),
.B2(n_4494),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4500),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4482),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4498),
.Y(n_4515)
);

NOR3xp33_ASAP7_75t_L g4516 ( 
.A(n_4503),
.B(n_4486),
.C(n_4495),
.Y(n_4516)
);

HB1xp67_ASAP7_75t_L g4517 ( 
.A(n_4506),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4510),
.Y(n_4518)
);

NOR2xp33_ASAP7_75t_L g4519 ( 
.A(n_4509),
.B(n_4501),
.Y(n_4519)
);

OA22x2_ASAP7_75t_L g4520 ( 
.A1(n_4514),
.A2(n_804),
.B1(n_730),
.B2(n_731),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4510),
.Y(n_4521)
);

AOI22xp5_ASAP7_75t_L g4522 ( 
.A1(n_4507),
.A2(n_728),
.B1(n_731),
.B2(n_732),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_4513),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4515),
.Y(n_4524)
);

NOR2x1_ASAP7_75t_L g4525 ( 
.A(n_4504),
.B(n_732),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4505),
.Y(n_4526)
);

CKINVDCx20_ASAP7_75t_R g4527 ( 
.A(n_4522),
.Y(n_4527)
);

AO211x2_ASAP7_75t_L g4528 ( 
.A1(n_4516),
.A2(n_4511),
.B(n_4508),
.C(n_4512),
.Y(n_4528)
);

AOI22xp5_ASAP7_75t_L g4529 ( 
.A1(n_4519),
.A2(n_4502),
.B1(n_734),
.B2(n_735),
.Y(n_4529)
);

AOI22xp5_ASAP7_75t_L g4530 ( 
.A1(n_4523),
.A2(n_733),
.B1(n_734),
.B2(n_736),
.Y(n_4530)
);

AND4x1_ASAP7_75t_L g4531 ( 
.A(n_4525),
.B(n_733),
.C(n_737),
.D(n_738),
.Y(n_4531)
);

NAND2xp5_ASAP7_75t_L g4532 ( 
.A(n_4518),
.B(n_737),
.Y(n_4532)
);

AO22x2_ASAP7_75t_L g4533 ( 
.A1(n_4521),
.A2(n_739),
.B1(n_740),
.B2(n_741),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4533),
.Y(n_4534)
);

AO22x2_ASAP7_75t_L g4535 ( 
.A1(n_4532),
.A2(n_4524),
.B1(n_4526),
.B2(n_4520),
.Y(n_4535)
);

OAI22xp5_ASAP7_75t_L g4536 ( 
.A1(n_4529),
.A2(n_4517),
.B1(n_741),
.B2(n_742),
.Y(n_4536)
);

INVx2_ASAP7_75t_L g4537 ( 
.A(n_4535),
.Y(n_4537)
);

AO22x2_ASAP7_75t_L g4538 ( 
.A1(n_4534),
.A2(n_4528),
.B1(n_4531),
.B2(n_4533),
.Y(n_4538)
);

INVxp67_ASAP7_75t_L g4539 ( 
.A(n_4537),
.Y(n_4539)
);

AOI22xp5_ASAP7_75t_L g4540 ( 
.A1(n_4539),
.A2(n_4527),
.B1(n_4538),
.B2(n_4536),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4540),
.Y(n_4541)
);

AOI22xp5_ASAP7_75t_L g4542 ( 
.A1(n_4541),
.A2(n_4530),
.B1(n_742),
.B2(n_743),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4542),
.Y(n_4543)
);

AOI221xp5_ASAP7_75t_L g4544 ( 
.A1(n_4543),
.A2(n_740),
.B1(n_743),
.B2(n_744),
.C(n_746),
.Y(n_4544)
);

AOI211xp5_ASAP7_75t_L g4545 ( 
.A1(n_4544),
.A2(n_747),
.B(n_748),
.C(n_749),
.Y(n_4545)
);


endmodule