module fake_jpeg_26018_n_90 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

BUFx10_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_52),
.Y(n_64)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_1),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_5),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_43),
.C(n_46),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_2),
.B(n_3),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_70),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_6),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_74),
.B(n_7),
.Y(n_77)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_69),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_77),
.B1(n_66),
.B2(n_59),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_SL g78 ( 
.A(n_73),
.B(n_71),
.C(n_9),
.Y(n_78)
);

AOI221xp5_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.C(n_14),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_80),
.B1(n_15),
.B2(n_17),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_65),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_56),
.B1(n_20),
.B2(n_21),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_86),
.B(n_23),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_89),
.B(n_32),
.CI(n_33),
.CON(n_90),
.SN(n_90)
);


endmodule