module real_jpeg_20879_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_1),
.A2(n_69),
.B1(n_70),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_1),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_1),
.A2(n_42),
.B1(n_49),
.B2(n_136),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_136),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_136),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_2),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_48),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_48),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_3),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_3),
.B(n_75),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_31),
.B(n_34),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_134),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_188),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_89),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_3),
.A2(n_49),
.B(n_219),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_69),
.B1(n_70),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_4),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_4),
.A2(n_42),
.B1(n_49),
.B2(n_116),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_116),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_116),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_5),
.A2(n_69),
.B1(n_70),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_5),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_42),
.B1(n_49),
.B2(n_77),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_77),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_77),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_69),
.B1(n_70),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_6),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_6),
.A2(n_42),
.B1(n_49),
.B2(n_94),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_94),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_94),
.Y(n_222)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_8),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_8),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_8),
.A2(n_42),
.B1(n_49),
.B2(n_71),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_71),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_71),
.Y(n_206)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_11),
.A2(n_42),
.B1(n_49),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_51),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_14),
.A2(n_30),
.A3(n_49),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_15),
.A2(n_42),
.B1(n_49),
.B2(n_73),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_118),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_117),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_97),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_22),
.B(n_97),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_79),
.B2(n_96),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_53),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_40),
.B(n_52),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_40),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_27),
.A2(n_33),
.B1(n_36),
.B2(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_27),
.A2(n_33),
.B1(n_63),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_27),
.A2(n_33),
.B1(n_84),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_27),
.A2(n_33),
.B1(n_109),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_27),
.A2(n_33),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_27),
.A2(n_33),
.B1(n_184),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_27),
.A2(n_33),
.B1(n_204),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_27),
.A2(n_33),
.B1(n_127),
.B2(n_222),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_29),
.B(n_43),
.Y(n_214)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_30),
.A2(n_32),
.B(n_134),
.C(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_31),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_33),
.B(n_134),
.Y(n_189)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

NAND2x1_ASAP7_75t_SL g56 ( 
.A(n_34),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_35),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_40)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_41),
.A2(n_45),
.B1(n_87),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_41),
.A2(n_45),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_41),
.A2(n_45),
.B1(n_112),
.B2(n_131),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_41),
.A2(n_45),
.B1(n_158),
.B2(n_218),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.Y(n_44)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_42),
.A2(n_74),
.B1(n_133),
.B2(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_42),
.B(n_134),
.Y(n_215)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_49),
.B(n_73),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_64),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_62),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_65),
.B1(n_66),
.B2(n_78),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_62),
.B1(n_78),
.B2(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_58),
.B(n_61),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_56),
.A2(n_57),
.B1(n_82),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_56),
.A2(n_60),
.B1(n_107),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_56),
.A2(n_60),
.B1(n_148),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_56),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_56),
.A2(n_57),
.B1(n_174),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_56),
.A2(n_57),
.B1(n_176),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_56),
.A2(n_58),
.B1(n_163),
.B2(n_206),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_57),
.B(n_134),
.Y(n_192)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_59),
.A2(n_172),
.B1(n_173),
.B2(n_175),
.Y(n_171)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_62),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_73),
.B(n_74),
.C(n_75),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_73),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_70),
.B(n_134),
.CON(n_133),
.SN(n_133)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_72),
.A2(n_75),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.C(n_90),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_81),
.B(n_83),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_88),
.A2(n_89),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_92),
.A2(n_95),
.B1(n_115),
.B2(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.C(n_104),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_102),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_104),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_110),
.C(n_113),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_105),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_260),
.B(n_265),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_164),
.B(n_247),
.C(n_259),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_149),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_121),
.B(n_149),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_137),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_123),
.B(n_124),
.C(n_137),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.C(n_132),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_139),
.B(n_143),
.C(n_144),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_147),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_154),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_150),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.C(n_161),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_156),
.B(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_160),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_246),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_241),
.B(n_245),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_227),
.B(n_240),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_208),
.B(n_226),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_196),
.B(n_207),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_185),
.B(n_195),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_177),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_181),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_190),
.B(n_194),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_189),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_198),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_203),
.C(n_205),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_210),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_216),
.B1(n_224),
.B2(n_225),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_211),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_213),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_216),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_220),
.B1(n_221),
.B2(n_223),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_217),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_223),
.C(n_224),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_229),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_237),
.C(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_236),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_237),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_249),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_258),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_250),
.Y(n_258)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_256),
.C(n_258),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);


endmodule