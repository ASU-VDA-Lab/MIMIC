module fake_jpeg_28447_n_108 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_2),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_7),
.B(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_53),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_37),
.B1(n_36),
.B2(n_48),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_17),
.B1(n_31),
.B2(n_30),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_44),
.C(n_37),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_41),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_0),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_36),
.B1(n_46),
.B2(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_75),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_81),
.C(n_4),
.Y(n_82)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_46),
.B(n_1),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_81),
.C(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_35),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_46),
.B(n_55),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_77),
.B(n_80),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_32),
.B1(n_14),
.B2(n_18),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_79),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_29),
.B1(n_13),
.B2(n_22),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_86),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_10),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_93),
.C(n_82),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_23),
.B(n_28),
.C(n_11),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_87),
.C(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_100),
.B(n_101),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_83),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_102),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_94),
.B(n_96),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_96),
.B(n_91),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_92),
.Y(n_108)
);


endmodule