module fake_jpeg_24978_n_86 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_1),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_2),
.B(n_3),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_12),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_42),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_59),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_51),
.B1(n_49),
.B2(n_20),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_18),
.C(n_19),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_54),
.C(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_78),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_77),
.A2(n_75),
.B(n_74),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_70),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_68),
.C(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_82),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_65),
.Y(n_86)
);


endmodule