module fake_jpeg_21224_n_68 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_SL g42 ( 
.A(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_31),
.B(n_1),
.C(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_30),
.Y(n_50)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_52),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_53),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_8),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_54),
.A2(n_55),
.B(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_44),
.B(n_11),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_16),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_18),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_61),
.C(n_56),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_57),
.B(n_51),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_19),
.C(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_25),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);


endmodule