module real_aes_9965_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_707, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_707;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_87;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
AOI22xp33_ASAP7_75t_SL g569 ( .A1(n_0), .A2(n_20), .B1(n_558), .B2(n_559), .Y(n_569) );
INVxp67_ASAP7_75t_SL g641 ( .A(n_0), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_1), .B(n_56), .Y(n_506) );
AND2x2_ASAP7_75t_L g529 ( .A(n_1), .B(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_1), .Y(n_555) );
INVx1_ASAP7_75t_L g575 ( .A(n_1), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_2), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_3), .B(n_115), .Y(n_161) );
INVx2_ASAP7_75t_L g590 ( .A(n_4), .Y(n_590) );
OR2x2_ASAP7_75t_L g605 ( .A(n_4), .B(n_588), .Y(n_605) );
OR2x2_ASAP7_75t_L g505 ( .A(n_5), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g528 ( .A(n_5), .Y(n_528) );
BUFx2_ASAP7_75t_L g552 ( .A(n_5), .Y(n_552) );
BUFx2_ASAP7_75t_L g584 ( .A(n_5), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_6), .B(n_122), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_7), .B(n_107), .Y(n_126) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_8), .A2(n_51), .B1(n_558), .B2(n_559), .Y(n_557) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_8), .A2(n_73), .B1(n_643), .B2(n_644), .C(n_647), .Y(n_642) );
NAND2x1p5_ASAP7_75t_L g202 ( .A(n_9), .B(n_107), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_10), .B(n_157), .Y(n_233) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_11), .A2(n_27), .B1(n_563), .B2(n_565), .Y(n_568) );
INVxp33_ASAP7_75t_SL g664 ( .A(n_11), .Y(n_664) );
AND2x2_ASAP7_75t_L g176 ( .A(n_12), .B(n_177), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_13), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_14), .A2(n_493), .B1(n_494), .B2(n_688), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_14), .Y(n_688) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_15), .Y(n_92) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_16), .B(n_239), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_17), .B(n_165), .Y(n_164) );
NAND2xp33_ASAP7_75t_L g195 ( .A(n_18), .B(n_114), .Y(n_195) );
NAND2xp33_ASAP7_75t_L g123 ( .A(n_19), .B(n_114), .Y(n_123) );
INVxp33_ASAP7_75t_L g661 ( .A(n_20), .Y(n_661) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_21), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_22), .Y(n_134) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_23), .Y(n_490) );
INVx1_ASAP7_75t_L g588 ( .A(n_24), .Y(n_588) );
INVx1_ASAP7_75t_L g635 ( .A(n_24), .Y(n_635) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_25), .Y(n_507) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_25), .A2(n_60), .B1(n_607), .B2(n_612), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_26), .Y(n_480) );
INVxp67_ASAP7_75t_SL g599 ( .A(n_27), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_28), .B(n_201), .Y(n_200) );
OAI21x1_ASAP7_75t_L g109 ( .A1(n_29), .A2(n_46), .B(n_110), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_30), .A2(n_140), .B(n_182), .C(n_183), .Y(n_181) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_30), .Y(n_701) );
NAND2xp33_ASAP7_75t_L g236 ( .A(n_31), .B(n_144), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_32), .B(n_138), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_33), .Y(n_255) );
AND2x6_ASAP7_75t_L g82 ( .A(n_34), .B(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_34), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_34), .B(n_675), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_35), .B(n_137), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_36), .B(n_121), .Y(n_120) );
NAND2xp33_ASAP7_75t_L g162 ( .A(n_37), .B(n_144), .Y(n_162) );
INVx1_ASAP7_75t_L g83 ( .A(n_38), .Y(n_83) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_38), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_39), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_40), .B(n_144), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_41), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_42), .Y(n_251) );
AND2x2_ASAP7_75t_L g185 ( .A(n_43), .B(n_165), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_44), .B(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g513 ( .A(n_45), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_47), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_48), .Y(n_535) );
NAND2xp33_ASAP7_75t_L g218 ( .A(n_49), .B(n_89), .Y(n_218) );
INVxp33_ASAP7_75t_SL g540 ( .A(n_50), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_50), .A2(n_65), .B1(n_618), .B2(n_621), .C(n_625), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_51), .A2(n_58), .B1(n_652), .B2(n_654), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_52), .B(n_194), .Y(n_235) );
BUFx10_ASAP7_75t_L g684 ( .A(n_53), .Y(n_684) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_54), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_55), .B(n_88), .Y(n_116) );
INVx2_ASAP7_75t_L g530 ( .A(n_56), .Y(n_530) );
INVx1_ASAP7_75t_L g556 ( .A(n_56), .Y(n_556) );
NAND2xp33_ASAP7_75t_L g223 ( .A(n_57), .B(n_122), .Y(n_223) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_58), .A2(n_73), .B1(n_563), .B2(n_565), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g113 ( .A(n_59), .B(n_114), .Y(n_113) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_59), .Y(n_485) );
INVxp67_ASAP7_75t_SL g514 ( .A(n_60), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_61), .Y(n_184) );
INVx1_ASAP7_75t_L g531 ( .A(n_62), .Y(n_531) );
INVx2_ASAP7_75t_L g110 ( .A(n_63), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_64), .Y(n_143) );
INVxp33_ASAP7_75t_SL g521 ( .A(n_65), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_66), .B(n_201), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_67), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_68), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g175 ( .A(n_69), .Y(n_175) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_69), .Y(n_699) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_70), .Y(n_136) );
AND2x2_ASAP7_75t_L g149 ( .A(n_71), .B(n_107), .Y(n_149) );
INVx2_ASAP7_75t_L g503 ( .A(n_72), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_74), .B(n_165), .Y(n_224) );
BUFx3_ASAP7_75t_L g593 ( .A(n_75), .Y(n_593) );
INVx1_ASAP7_75t_L g624 ( .A(n_75), .Y(n_624) );
BUFx3_ASAP7_75t_L g595 ( .A(n_76), .Y(n_595) );
INVx1_ASAP7_75t_L g603 ( .A(n_76), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_93), .B(n_475), .Y(n_77) );
AND2x2_ASAP7_75t_L g78 ( .A(n_79), .B(n_84), .Y(n_78) );
HB1xp67_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx8_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_81), .A2(n_132), .B(n_141), .Y(n_131) );
NOR2xp67_ASAP7_75t_L g170 ( .A(n_81), .B(n_171), .Y(n_170) );
INVx8_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
BUFx2_ASAP7_75t_L g237 ( .A(n_82), .Y(n_237) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_85), .Y(n_84) );
AO21x1_ASAP7_75t_L g703 ( .A1(n_85), .A2(n_704), .B(n_705), .Y(n_703) );
NAND2xp33_ASAP7_75t_L g85 ( .A(n_86), .B(n_91), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g252 ( .A(n_88), .Y(n_252) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx2_ASAP7_75t_L g157 ( .A(n_89), .Y(n_157) );
INVx2_ASAP7_75t_L g220 ( .A(n_89), .Y(n_220) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_90), .Y(n_122) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_90), .Y(n_147) );
INVx1_ASAP7_75t_L g179 ( .A(n_90), .Y(n_179) );
INVx1_ASAP7_75t_L g124 ( .A(n_91), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_91), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21x1_ASAP7_75t_L g231 ( .A1(n_91), .A2(n_232), .B(n_233), .Y(n_231) );
INVx5_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
BUFx12f_ASAP7_75t_L g118 ( .A(n_92), .Y(n_118) );
INVx5_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_92), .A2(n_251), .B(n_252), .C(n_253), .Y(n_250) );
HB1xp67_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx2_ASAP7_75t_SL g95 ( .A(n_96), .Y(n_95) );
BUFx3_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
NAND2x1p5_ASAP7_75t_L g97 ( .A(n_98), .B(n_392), .Y(n_97) );
AND5x1_ASAP7_75t_L g98 ( .A(n_99), .B(n_295), .C(n_334), .D(n_360), .E(n_375), .Y(n_98) );
NOR2xp33_ASAP7_75t_L g99 ( .A(n_100), .B(n_262), .Y(n_99) );
OAI221xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_186), .B1(n_203), .B2(n_213), .C(n_241), .Y(n_100) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_127), .Y(n_101) );
INVx1_ASAP7_75t_L g359 ( .A(n_102), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_102), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_102), .B(n_244), .Y(n_443) );
AOI322xp5_ASAP7_75t_L g456 ( .A1(n_102), .A2(n_325), .A3(n_378), .B1(n_457), .B2(n_459), .C1(n_460), .C2(n_463), .Y(n_456) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g344 ( .A(n_103), .B(n_211), .Y(n_344) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_104), .Y(n_212) );
INVx1_ASAP7_75t_L g279 ( .A(n_104), .Y(n_279) );
AND2x2_ASAP7_75t_L g284 ( .A(n_104), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g294 ( .A(n_104), .B(n_208), .Y(n_294) );
AND2x2_ASAP7_75t_L g302 ( .A(n_104), .B(n_150), .Y(n_302) );
INVx1_ASAP7_75t_L g316 ( .A(n_104), .Y(n_316) );
OAI21x1_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_111), .B(n_126), .Y(n_104) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_105), .A2(n_230), .B(n_238), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_105), .A2(n_230), .B(n_238), .Y(n_258) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx4_ASAP7_75t_L g130 ( .A(n_107), .Y(n_130) );
BUFx4f_ASAP7_75t_L g152 ( .A(n_107), .Y(n_152) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_107), .A2(n_216), .B(n_224), .Y(n_215) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_107), .A2(n_216), .B(n_224), .Y(n_261) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_107), .A2(n_216), .B(n_224), .Y(n_266) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g240 ( .A(n_108), .Y(n_240) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g166 ( .A(n_109), .Y(n_166) );
OAI21x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_119), .B(n_125), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_116), .B(n_117), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_114), .B(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g144 ( .A(n_115), .Y(n_144) );
INVx1_ASAP7_75t_L g201 ( .A(n_115), .Y(n_201) );
OAI21xp33_ASAP7_75t_L g141 ( .A1(n_117), .A2(n_142), .B(n_145), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx3_ASAP7_75t_L g159 ( .A(n_118), .Y(n_159) );
BUFx2_ASAP7_75t_L g180 ( .A(n_118), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_118), .A2(n_235), .B(n_236), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_123), .B(n_124), .Y(n_119) );
INVx2_ASAP7_75t_L g182 ( .A(n_121), .Y(n_182) );
INVx2_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_122), .B(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g194 ( .A(n_122), .Y(n_194) );
INVx2_ASAP7_75t_L g199 ( .A(n_122), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g153 ( .A1(n_125), .A2(n_154), .B(n_160), .Y(n_153) );
OAI21x1_ASAP7_75t_L g191 ( .A1(n_125), .A2(n_192), .B(n_196), .Y(n_191) );
OAI21x1_ASAP7_75t_L g216 ( .A1(n_125), .A2(n_217), .B(n_221), .Y(n_216) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_125), .A2(n_250), .B(n_254), .Y(n_249) );
INVx1_ASAP7_75t_L g445 ( .A(n_127), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_167), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_150), .Y(n_128) );
INVx1_ASAP7_75t_L g283 ( .A(n_129), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_129), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_SL g327 ( .A(n_129), .Y(n_327) );
AO21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B(n_149), .Y(n_129) );
INVx3_ASAP7_75t_L g171 ( .A(n_130), .Y(n_171) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_130), .A2(n_131), .B(n_149), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_135), .B(n_139), .Y(n_132) );
NOR2xp67_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
INVx5_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
CKINVDCx6p67_ASAP7_75t_R g163 ( .A(n_140), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
NOR2xp33_ASAP7_75t_SL g145 ( .A(n_146), .B(n_148), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_146), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OR2x2_ASAP7_75t_L g278 ( .A(n_150), .B(n_279), .Y(n_278) );
BUFx3_ASAP7_75t_L g332 ( .A(n_150), .Y(n_332) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g211 ( .A(n_151), .Y(n_211) );
AND2x2_ASAP7_75t_L g309 ( .A(n_151), .B(n_208), .Y(n_309) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_164), .Y(n_151) );
OAI21x1_ASAP7_75t_L g190 ( .A1(n_152), .A2(n_191), .B(n_202), .Y(n_190) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_152), .A2(n_249), .B(n_257), .Y(n_248) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_152), .A2(n_249), .B(n_257), .Y(n_271) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_152), .A2(n_191), .B(n_202), .Y(n_290) );
O2A1O1Ixp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_158), .C(n_159), .Y(n_154) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
O2A1O1Ixp5_ASAP7_75t_L g196 ( .A1(n_159), .A2(n_197), .B(n_198), .C(n_200), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_159), .A2(n_198), .B(n_255), .C(n_256), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_163), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_163), .A2(n_193), .B(n_195), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_163), .A2(n_218), .B(n_219), .Y(n_217) );
BUFx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_167), .B(n_211), .Y(n_472) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_168), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_168), .B(n_211), .Y(n_317) );
INVx1_ASAP7_75t_L g342 ( .A(n_168), .Y(n_342) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g207 ( .A(n_169), .Y(n_207) );
AOI21x1_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_172), .B(n_185), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_181), .Y(n_172) );
OAI21x1_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_176), .B(n_180), .Y(n_173) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_186), .A2(n_429), .B1(n_432), .B2(n_433), .Y(n_428) );
INVx1_ASAP7_75t_L g432 ( .A(n_186), .Y(n_432) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2x1_ASAP7_75t_L g312 ( .A(n_187), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g260 ( .A(n_188), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g300 ( .A(n_188), .B(n_261), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_188), .B(n_289), .Y(n_338) );
OR2x2_ASAP7_75t_L g390 ( .A(n_188), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g272 ( .A(n_189), .B(n_228), .Y(n_272) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g227 ( .A(n_190), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_209), .Y(n_204) );
INVx1_ASAP7_75t_L g384 ( .A(n_205), .Y(n_384) );
NAND2xp67_ASAP7_75t_L g415 ( .A(n_205), .B(n_302), .Y(n_415) );
INVx1_ASAP7_75t_L g458 ( .A(n_205), .Y(n_458) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_208), .Y(n_205) );
INVx1_ASAP7_75t_L g293 ( .A(n_206), .Y(n_293) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g244 ( .A(n_207), .B(n_208), .Y(n_244) );
INVx1_ASAP7_75t_L g285 ( .A(n_207), .Y(n_285) );
AND2x2_ASAP7_75t_L g326 ( .A(n_207), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g346 ( .A(n_210), .B(n_243), .Y(n_346) );
OR2x2_ASAP7_75t_L g374 ( .A(n_210), .B(n_275), .Y(n_374) );
OR2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
INVx2_ASAP7_75t_L g351 ( .A(n_211), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_211), .B(n_283), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_225), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_214), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g331 ( .A(n_214), .B(n_332), .Y(n_331) );
NAND4xp25_ASAP7_75t_L g358 ( .A(n_214), .B(n_275), .C(n_281), .D(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g376 ( .A(n_214), .B(n_268), .Y(n_376) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g287 ( .A(n_215), .Y(n_287) );
AND2x2_ASAP7_75t_L g468 ( .A(n_215), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g412 ( .A(n_225), .Y(n_412) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g281 ( .A(n_227), .B(n_269), .Y(n_281) );
BUFx2_ASAP7_75t_L g306 ( .A(n_227), .Y(n_306) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_227), .B(n_367), .Y(n_407) );
INVx2_ASAP7_75t_L g289 ( .A(n_228), .Y(n_289) );
OR2x2_ASAP7_75t_L g403 ( .A(n_228), .B(n_248), .Y(n_403) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OAI21x1_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_234), .B(n_237), .Y(n_230) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_245), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_242), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_244), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g361 ( .A(n_244), .B(n_277), .Y(n_361) );
AND2x2_ASAP7_75t_L g454 ( .A(n_244), .B(n_430), .Y(n_454) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_259), .Y(n_245) );
INVx2_ASAP7_75t_L g461 ( .A(n_246), .Y(n_461) );
BUFx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_247), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_258), .Y(n_247) );
INVx1_ASAP7_75t_L g305 ( .A(n_248), .Y(n_305) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp33_ASAP7_75t_R g349 ( .A(n_260), .B(n_304), .Y(n_349) );
INVx1_ASAP7_75t_L g448 ( .A(n_260), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_261), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g355 ( .A(n_261), .Y(n_355) );
OAI21xp33_ASAP7_75t_SL g262 ( .A1(n_263), .A2(n_273), .B(n_280), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
O2A1O1Ixp5_ASAP7_75t_L g334 ( .A1(n_264), .A2(n_335), .B(n_339), .C(n_345), .Y(n_334) );
NOR2x1p5_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g311 ( .A(n_266), .Y(n_311) );
BUFx2_ASAP7_75t_L g322 ( .A(n_266), .Y(n_322) );
INVx2_ASAP7_75t_SL g391 ( .A(n_266), .Y(n_391) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
AND2x4_ASAP7_75t_L g297 ( .A(n_269), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g313 ( .A(n_271), .Y(n_313) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_271), .Y(n_337) );
AND2x2_ASAP7_75t_L g320 ( .A(n_272), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g467 ( .A(n_272), .Y(n_467) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g450 ( .A(n_275), .Y(n_450) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g371 ( .A(n_278), .Y(n_371) );
INVx1_ASAP7_75t_SL g381 ( .A(n_278), .Y(n_381) );
OR2x2_ASAP7_75t_L g417 ( .A(n_278), .B(n_341), .Y(n_417) );
OR2x2_ASAP7_75t_L g439 ( .A(n_278), .B(n_427), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B1(n_286), .B2(n_291), .Y(n_280) );
INVx2_ASAP7_75t_L g373 ( .A(n_281), .Y(n_373) );
INVx1_ASAP7_75t_L g323 ( .A(n_282), .Y(n_323) );
AND2x4_ASAP7_75t_L g405 ( .A(n_282), .B(n_351), .Y(n_405) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
BUFx2_ASAP7_75t_SL g434 ( .A(n_283), .Y(n_434) );
AND2x4_ASAP7_75t_L g308 ( .A(n_284), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g399 ( .A(n_284), .Y(n_399) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
OR2x6_ASAP7_75t_SL g402 ( .A(n_287), .B(n_403), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g452 ( .A1(n_287), .A2(n_453), .B(n_456), .C(n_464), .Y(n_452) );
AND2x2_ASAP7_75t_L g459 ( .A(n_287), .B(n_407), .Y(n_459) );
INVx2_ASAP7_75t_L g368 ( .A(n_288), .Y(n_368) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx2_ASAP7_75t_L g298 ( .A(n_289), .Y(n_298) );
INVx2_ASAP7_75t_L g356 ( .A(n_290), .Y(n_356) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g377 ( .A(n_293), .Y(n_377) );
INVxp67_ASAP7_75t_SL g333 ( .A(n_294), .Y(n_333) );
INVx2_ASAP7_75t_L g352 ( .A(n_294), .Y(n_352) );
OR2x2_ASAP7_75t_L g409 ( .A(n_294), .B(n_342), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_318), .Y(n_295) );
OAI332xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_299), .A3(n_301), .B1(n_303), .B2(n_306), .B3(n_307), .C1(n_310), .C2(n_314), .Y(n_296) );
INVx2_ASAP7_75t_L g369 ( .A(n_297), .Y(n_369) );
AND2x4_ASAP7_75t_SL g329 ( .A(n_298), .B(n_313), .Y(n_329) );
BUFx2_ASAP7_75t_L g436 ( .A(n_298), .Y(n_436) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI311xp33_ASAP7_75t_L g345 ( .A1(n_300), .A2(n_346), .A3(n_347), .B1(n_348), .C1(n_358), .Y(n_345) );
AND2x2_ASAP7_75t_L g362 ( .A(n_300), .B(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_301), .A2(n_365), .B1(n_369), .B2(n_370), .Y(n_364) );
AND2x4_ASAP7_75t_L g325 ( .A(n_302), .B(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g367 ( .A(n_305), .Y(n_367) );
NAND3xp33_ASAP7_75t_L g330 ( .A(n_306), .B(n_331), .C(n_333), .Y(n_330) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_306), .A2(n_357), .B1(n_407), .B2(n_408), .Y(n_406) );
INVx2_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
OR2x2_ASAP7_75t_L g401 ( .A(n_311), .B(n_368), .Y(n_401) );
BUFx2_ASAP7_75t_L g347 ( .A(n_313), .Y(n_347) );
INVx1_ASAP7_75t_L g363 ( .A(n_313), .Y(n_363) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
OR2x2_ASAP7_75t_L g474 ( .A(n_315), .B(n_472), .Y(n_474) );
INVx1_ASAP7_75t_L g431 ( .A(n_316), .Y(n_431) );
INVx1_ASAP7_75t_L g387 ( .A(n_317), .Y(n_387) );
OAI221xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_323), .B1(n_324), .B2(n_328), .C(n_330), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g357 ( .A(n_326), .B(n_332), .Y(n_357) );
AND2x2_ASAP7_75t_L g380 ( .A(n_326), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g440 ( .A(n_326), .Y(n_440) );
INVx2_ASAP7_75t_L g413 ( .A(n_329), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_329), .A2(n_436), .B1(n_454), .B2(n_455), .Y(n_453) );
AND2x2_ASAP7_75t_L g470 ( .A(n_333), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_337), .Y(n_389) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_337), .Y(n_447) );
INVx1_ASAP7_75t_L g469 ( .A(n_338), .Y(n_469) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B1(n_353), .B2(n_357), .Y(n_348) );
INVx3_ASAP7_75t_L g451 ( .A(n_350), .Y(n_451) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AOI321xp33_ASAP7_75t_L g375 ( .A1(n_351), .A2(n_376), .A3(n_377), .B1(n_378), .B2(n_380), .C(n_382), .Y(n_375) );
OR2x2_ASAP7_75t_L g383 ( .A(n_351), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g424 ( .A(n_351), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g386 ( .A(n_352), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g379 ( .A(n_354), .Y(n_379) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_354), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AOI211xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B(n_364), .C(n_372), .Y(n_360) );
AOI222xp33_ASAP7_75t_L g464 ( .A1(n_361), .A2(n_465), .B1(n_468), .B2(n_470), .C1(n_473), .C2(n_707), .Y(n_464) );
NAND2x1_ASAP7_75t_L g404 ( .A(n_362), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g378 ( .A(n_363), .B(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI32xp33_ASAP7_75t_L g449 ( .A1(n_368), .A2(n_403), .A3(n_439), .B1(n_450), .B2(n_451), .Y(n_449) );
NOR2xp67_ASAP7_75t_SL g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g463 ( .A(n_374), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_377), .B(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_379), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .B(n_388), .Y(n_382) );
INVx1_ASAP7_75t_L g455 ( .A(n_383), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_385), .A2(n_417), .B1(n_418), .B2(n_421), .Y(n_416) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
INVx1_ASAP7_75t_L g427 ( .A(n_391), .Y(n_427) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_393), .B(n_452), .Y(n_392) );
NAND4xp75_ASAP7_75t_L g393 ( .A(n_394), .B(n_410), .C(n_423), .D(n_441), .Y(n_393) );
AND3x1_ASAP7_75t_L g394 ( .A(n_395), .B(n_404), .C(n_406), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_400), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
NAND2xp33_ASAP7_75t_SL g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx2_ASAP7_75t_L g419 ( .A(n_403), .Y(n_419) );
OR2x2_ASAP7_75t_L g426 ( .A(n_403), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_414), .B(n_416), .Y(n_410) );
NAND2xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2x1_ASAP7_75t_SL g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI21x1_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_428), .B(n_435), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NOR2x1_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR2x1_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_446), .B(n_449), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OAI221xp5_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_671), .B1(n_687), .B2(n_689), .C(n_694), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B1(n_493), .B2(n_494), .Y(n_476) );
CKINVDCx14_ASAP7_75t_R g477 ( .A(n_478), .Y(n_477) );
XNOR2xp5_ASAP7_75t_SL g478 ( .A(n_479), .B(n_484), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_482), .B2(n_483), .Y(n_479) );
INVx1_ASAP7_75t_L g482 ( .A(n_480), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_481), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_487), .B2(n_492), .Y(n_484) );
INVx1_ASAP7_75t_L g492 ( .A(n_485), .Y(n_492) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_487) );
INVx1_ASAP7_75t_L g491 ( .A(n_488), .Y(n_491) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_493), .A2(n_494), .B1(n_699), .B2(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_576), .Y(n_495) );
AND4x1_ASAP7_75t_L g496 ( .A(n_497), .B(n_520), .C(n_534), .D(n_547), .Y(n_496) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_507), .B1(n_508), .B2(n_514), .C(n_515), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_504), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g518 ( .A(n_503), .Y(n_518) );
AND2x4_ASAP7_75t_L g526 ( .A(n_503), .B(n_519), .Y(n_526) );
AND2x2_ASAP7_75t_L g539 ( .A(n_503), .B(n_513), .Y(n_539) );
INVx2_ASAP7_75t_L g544 ( .A(n_503), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_503), .B(n_513), .Y(n_581) );
AND2x4_ASAP7_75t_L g510 ( .A(n_504), .B(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_L g515 ( .A(n_504), .B(n_516), .Y(n_515) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g579 ( .A(n_505), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g519 ( .A(n_513), .Y(n_519) );
INVx1_ASAP7_75t_L g546 ( .A(n_513), .Y(n_546) );
BUFx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx3_ASAP7_75t_L g533 ( .A(n_517), .Y(n_533) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_517), .Y(n_561) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B1(n_531), .B2(n_532), .Y(n_520) );
BUFx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_526), .Y(n_567) );
AND2x6_ASAP7_75t_L g532 ( .A(n_527), .B(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g536 ( .A(n_527), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g541 ( .A(n_527), .B(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g572 ( .A(n_528), .Y(n_572) );
INVx1_ASAP7_75t_L g574 ( .A(n_530), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_531), .A2(n_535), .B1(n_626), .B2(n_630), .C(n_633), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B1(n_540), .B2(n_541), .Y(n_534) );
BUFx3_ASAP7_75t_L g558 ( .A(n_537), .Y(n_558) );
INVx2_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_543), .Y(n_564) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI33xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_557), .A3(n_562), .B1(n_568), .B2(n_569), .B3(n_570), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx2_ASAP7_75t_L g670 ( .A(n_552), .Y(n_670) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
BUFx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
INVx6_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x6_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_596), .B(n_597), .Y(n_576) );
INVx5_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_591), .Y(n_585) );
AND2x4_ASAP7_75t_L g608 ( .A(n_586), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g613 ( .A(n_586), .Y(n_613) );
AND2x4_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g634 ( .A(n_589), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g650 ( .A(n_590), .B(n_635), .Y(n_650) );
INVx2_ASAP7_75t_L g653 ( .A(n_591), .Y(n_653) );
AND2x4_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
INVx1_ASAP7_75t_L g616 ( .A(n_592), .Y(n_616) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g602 ( .A(n_593), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g640 ( .A(n_593), .B(n_595), .Y(n_640) );
INVx1_ASAP7_75t_L g611 ( .A(n_594), .Y(n_611) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g623 ( .A(n_595), .B(n_624), .Y(n_623) );
AOI31xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_636), .A3(n_660), .B(n_668), .Y(n_597) );
AOI211xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B(n_606), .C(n_617), .Y(n_598) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_602), .Y(n_620) );
INVx1_ASAP7_75t_L g629 ( .A(n_603), .Y(n_629) );
AND2x4_ASAP7_75t_L g638 ( .A(n_604), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g663 ( .A(n_605), .B(n_632), .Y(n_663) );
OR2x2_ASAP7_75t_L g666 ( .A(n_605), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_SL g686 ( .A(n_608), .Y(n_686) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g682 ( .A(n_610), .Y(n_682) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_SL g657 ( .A(n_613), .Y(n_657) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx3_ASAP7_75t_L g643 ( .A(n_620), .Y(n_643) );
BUFx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_623), .Y(n_655) );
INVx2_ASAP7_75t_L g667 ( .A(n_623), .Y(n_667) );
INVx1_ASAP7_75t_L g628 ( .A(n_624), .Y(n_628) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
OR2x2_ASAP7_75t_L g632 ( .A(n_628), .B(n_629), .Y(n_632) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_641), .B1(n_642), .B2(n_651), .C(n_656), .Y(n_636) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_639), .Y(n_646) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_640), .Y(n_659) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx2_ASAP7_75t_L g679 ( .A(n_649), .Y(n_679) );
INVx2_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B1(n_664), .B2(n_665), .Y(n_660) );
INVx6_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx4_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
BUFx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx8_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
CKINVDCx20_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OR2x6_ASAP7_75t_L g673 ( .A(n_674), .B(n_677), .Y(n_673) );
OR2x4_ASAP7_75t_L g697 ( .A(n_674), .B(n_678), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_675), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g704 ( .A(n_675), .Y(n_704) );
INVx1_ASAP7_75t_L g693 ( .A(n_676), .Y(n_693) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AOI31xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .A3(n_683), .B(n_685), .Y(n_678) );
INVxp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx6_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
BUFx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_698), .B1(n_701), .B2(n_702), .Y(n_694) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx8_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
CKINVDCx5p33_ASAP7_75t_R g700 ( .A(n_699), .Y(n_700) );
BUFx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
endmodule