module fake_netlist_5_1075_n_1222 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1222);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1222;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_977;
wire n_419;
wire n_653;
wire n_1194;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_1178;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_1161;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_1055;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_1191;
wire n_1198;
wire n_721;
wire n_998;
wire n_1157;
wire n_1099;
wire n_841;
wire n_1050;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_983;
wire n_725;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_629;
wire n_590;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_1110;
wire n_859;
wire n_1203;
wire n_951;
wire n_1121;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_1179;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1048;
wire n_932;
wire n_946;
wire n_417;
wire n_1008;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_212;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_1195;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_568;
wire n_509;
wire n_947;
wire n_373;
wire n_820;
wire n_936;
wire n_757;
wire n_1090;
wire n_1200;
wire n_307;
wire n_633;
wire n_1192;
wire n_530;
wire n_439;
wire n_1024;
wire n_1107;
wire n_1063;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1185;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_1143;
wire n_981;
wire n_804;
wire n_867;
wire n_186;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_1104;
wire n_792;
wire n_563;
wire n_1182;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_1163;
wire n_406;
wire n_519;
wire n_919;
wire n_908;
wire n_782;
wire n_470;
wire n_1108;
wire n_325;
wire n_449;
wire n_1100;
wire n_1207;
wire n_1214;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_1169;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_1221;
wire n_654;
wire n_370;
wire n_1172;
wire n_1095;
wire n_607;
wire n_976;
wire n_1096;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_1168;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1201;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_264;
wire n_669;
wire n_750;
wire n_742;
wire n_472;
wire n_454;
wire n_961;
wire n_1176;
wire n_955;
wire n_387;
wire n_771;
wire n_995;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_1149;
wire n_882;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_696;
wire n_1073;
wire n_255;
wire n_897;
wire n_798;
wire n_350;
wire n_196;
wire n_215;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_181;
wire n_436;
wire n_962;
wire n_1219;
wire n_1204;
wire n_1215;
wire n_1216;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_1171;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_1218;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1188;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_1165;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_681;
wire n_584;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_1177;
wire n_680;
wire n_974;
wire n_395;
wire n_553;
wire n_432;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_1159;
wire n_1210;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_328;
wire n_214;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_685;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_829;
wire n_928;
wire n_749;
wire n_1064;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_1173;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_1193;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_1197;
wire n_1211;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1187;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_1164;
wire n_420;
wire n_630;
wire n_1202;
wire n_489;
wire n_632;
wire n_699;
wire n_1174;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_846;
wire n_586;
wire n_1058;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_1101;
wire n_1053;
wire n_273;
wire n_1106;
wire n_585;
wire n_349;
wire n_1190;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_1116;
wire n_954;
wire n_627;
wire n_1212;
wire n_767;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_1175;
wire n_861;
wire n_534;
wire n_948;
wire n_1183;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_1217;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1131;
wire n_1059;
wire n_1084;
wire n_176;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_1005;
wire n_354;
wire n_647;
wire n_575;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_707;
wire n_795;
wire n_832;
wire n_695;
wire n_857;
wire n_180;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1220;
wire n_1044;
wire n_1205;
wire n_346;
wire n_937;
wire n_1209;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_1027;
wire n_490;
wire n_805;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_1037;
wire n_1160;
wire n_202;
wire n_1080;
wire n_266;
wire n_1162;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_1199;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_797;
wire n_409;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_1181;
wire n_1196;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_1213;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1186;
wire n_1004;
wire n_242;
wire n_817;
wire n_1032;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_200;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_1155;
wire n_438;
wire n_806;
wire n_522;
wire n_713;
wire n_1011;
wire n_1123;
wire n_1184;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_1189;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_1180;
wire n_1206;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_1170;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g175 ( 
.A(n_25),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_55),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_48),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_146),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_98),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_26),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_124),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_158),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_76),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_41),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_157),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_89),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_99),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_64),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_62),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_114),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_144),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_15),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_56),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_75),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_93),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

CKINVDCx11_ASAP7_75t_R g202 ( 
.A(n_19),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_108),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_100),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_101),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_148),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_14),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_133),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_70),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_136),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_20),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_9),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_32),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_115),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_2),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_130),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_147),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_156),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_107),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_19),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_8),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_110),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_6),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_73),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_85),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_90),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_202),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_176),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_177),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_183),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_178),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_183),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_184),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_185),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_187),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_188),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_189),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_193),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_190),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_182),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_194),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_195),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_196),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_200),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_197),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_203),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_204),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_206),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_231),
.Y(n_261)
);

BUFx8_ASAP7_75t_SL g262 ( 
.A(n_233),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_199),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_239),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_235),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_238),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_254),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_240),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_229),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_241),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_244),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_247),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_248),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_249),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_234),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_234),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_250),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_248),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_230),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_230),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_230),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_230),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_230),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_230),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_245),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_248),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_230),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_245),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_245),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_264),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_262),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_276),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_262),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_258),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_260),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_303),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_263),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_308),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_283),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_264),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g335 ( 
.A(n_265),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_299),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_302),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_267),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_259),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_291),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_292),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_299),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_293),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_281),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_280),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_265),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_261),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_339),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_320),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_316),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_351),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_339),
.Y(n_359)
);

INVxp33_ASAP7_75t_SL g360 ( 
.A(n_343),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_351),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_320),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_323),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_342),
.B(n_352),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_311),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_351),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_317),
.Y(n_368)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_319),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_343),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_309),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_311),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_342),
.B(n_266),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_321),
.B(n_266),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_314),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_314),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_310),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_309),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_333),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_312),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_313),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_315),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_333),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_335),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_335),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_349),
.Y(n_392)
);

INVxp33_ASAP7_75t_SL g393 ( 
.A(n_353),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_335),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_326),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_322),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_324),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_364),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_395),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_379),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_375),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_378),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_395),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_298),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_350),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_370),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_379),
.B(n_344),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_392),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_388),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_371),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_373),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_366),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_382),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_363),
.A2(n_326),
.B(n_341),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_397),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_385),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_356),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_396),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_345),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_387),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_358),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_361),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_390),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_369),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_390),
.B(n_325),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_356),
.B(n_338),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_393),
.A2(n_279),
.B1(n_329),
.B2(n_327),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_391),
.Y(n_437)
);

OA21x2_ASAP7_75t_L g438 ( 
.A1(n_391),
.A2(n_337),
.B(n_336),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_394),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_394),
.A2(n_346),
.B(n_340),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_362),
.B(n_331),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_362),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_389),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_360),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_376),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_360),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_365),
.B(n_354),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_355),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_359),
.A2(n_199),
.B1(n_228),
.B2(n_227),
.Y(n_450)
);

NOR2x1_ASAP7_75t_L g451 ( 
.A(n_365),
.B(n_279),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_378),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

AND2x6_ASAP7_75t_L g458 ( 
.A(n_379),
.B(n_347),
.Y(n_458)
);

OA21x2_ASAP7_75t_L g459 ( 
.A1(n_378),
.A2(n_332),
.B(n_330),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_357),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_357),
.B(n_269),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_364),
.A2(n_298),
.B1(n_271),
.B2(n_306),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_378),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_378),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_388),
.A2(n_227),
.B1(n_228),
.B2(n_300),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_395),
.B(n_273),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_357),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_379),
.B(n_179),
.Y(n_469)
);

OA21x2_ASAP7_75t_L g470 ( 
.A1(n_378),
.A2(n_191),
.B(n_186),
.Y(n_470)
);

CKINVDCx11_ASAP7_75t_R g471 ( 
.A(n_375),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_357),
.Y(n_472)
);

BUFx12f_ASAP7_75t_L g473 ( 
.A(n_374),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_392),
.B(n_323),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_374),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_364),
.B(n_278),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_364),
.B(n_285),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_364),
.B(n_294),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_403),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_403),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_407),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_414),
.B(n_295),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_414),
.B(n_296),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_415),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_407),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_398),
.B(n_297),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_401),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_404),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_323),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g490 ( 
.A(n_412),
.B(n_181),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_456),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_473),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_399),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_328),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_457),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_457),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_428),
.B(n_180),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_412),
.B(n_181),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_475),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_399),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_198),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_400),
.B(n_270),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_428),
.B(n_192),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_415),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_433),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_L g507 ( 
.A(n_458),
.B(n_208),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_463),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_411),
.B(n_201),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_463),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_464),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_464),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_465),
.Y(n_513)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_475),
.Y(n_514)
);

NAND2x1p5_ASAP7_75t_L g515 ( 
.A(n_408),
.B(n_205),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_465),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_459),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_478),
.B(n_209),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_459),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_406),
.B(n_210),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_408),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_408),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_492),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_508),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_500),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_508),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_498),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_500),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_488),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_514),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_510),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_492),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_R g533 ( 
.A(n_487),
.B(n_471),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_487),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_511),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_511),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_494),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_494),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_494),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_482),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_494),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_486),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_503),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_R g544 ( 
.A(n_484),
.B(n_473),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_503),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_482),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_512),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_493),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_483),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_506),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_483),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_484),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_497),
.B(n_476),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_484),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_479),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_505),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_505),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_505),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_502),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_502),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_502),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_R g563 ( 
.A(n_489),
.B(n_426),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_R g564 ( 
.A(n_533),
.B(n_438),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_554),
.B(n_476),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_524),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_549),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_526),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_542),
.B(n_518),
.C(n_520),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_549),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_552),
.B(n_450),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_530),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_553),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_531),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_549),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_540),
.A2(n_477),
.B1(n_462),
.B2(n_448),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_535),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_535),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_536),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_536),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_529),
.B(n_488),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_547),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_547),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_549),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_SL g585 ( 
.A(n_563),
.B(n_432),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_L g586 ( 
.A(n_551),
.B(n_477),
.C(n_466),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_548),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_548),
.B(n_461),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_543),
.B(n_435),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_556),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_538),
.B(n_422),
.Y(n_591)
);

AND3x2_ASAP7_75t_L g592 ( 
.A(n_527),
.B(n_426),
.C(n_448),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_545),
.B(n_504),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_556),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_534),
.B(n_449),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_529),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_529),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_538),
.B(n_422),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_557),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_555),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_546),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_558),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_559),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_560),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_525),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_561),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_562),
.B(n_422),
.Y(n_607)
);

INVxp33_ASAP7_75t_L g608 ( 
.A(n_544),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_537),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_550),
.B(n_416),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_539),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_528),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_541),
.Y(n_613)
);

OAI22x1_ASAP7_75t_L g614 ( 
.A1(n_532),
.A2(n_436),
.B1(n_453),
.B2(n_452),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_523),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_523),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_524),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_535),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_554),
.B(n_422),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_555),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_524),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_535),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_535),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_535),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_535),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_524),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_524),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_553),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_535),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_549),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_554),
.B(n_422),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_525),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_549),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_554),
.B(n_449),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_535),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_554),
.B(n_435),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_554),
.B(n_415),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_549),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_554),
.B(n_415),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_535),
.Y(n_640)
);

CKINVDCx6p67_ASAP7_75t_R g641 ( 
.A(n_523),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_535),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_554),
.B(n_425),
.Y(n_643)
);

BUFx8_ASAP7_75t_SL g644 ( 
.A(n_523),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_535),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_524),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_524),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_549),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_524),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_596),
.B(n_510),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_585),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_566),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_569),
.B(n_401),
.Y(n_654)
);

OR2x6_ASAP7_75t_L g655 ( 
.A(n_637),
.B(n_515),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_599),
.B(n_402),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_568),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_574),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_565),
.B(n_634),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_599),
.B(n_402),
.Y(n_660)
);

CKINVDCx16_ASAP7_75t_R g661 ( 
.A(n_573),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_634),
.B(n_513),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_578),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_617),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_579),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_586),
.A2(n_469),
.B1(n_458),
.B2(n_444),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_643),
.B(n_513),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_636),
.B(n_516),
.Y(n_668)
);

INVxp33_ASAP7_75t_L g669 ( 
.A(n_595),
.Y(n_669)
);

AO21x2_ASAP7_75t_L g670 ( 
.A1(n_637),
.A2(n_519),
.B(n_517),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_613),
.B(n_502),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_573),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_579),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_581),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_571),
.A2(n_469),
.B1(n_458),
.B2(n_421),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_639),
.B(n_621),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_596),
.B(n_516),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_587),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_626),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_639),
.B(n_517),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_613),
.B(n_589),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_610),
.B(n_421),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_587),
.Y(n_683)
);

INVx8_ASAP7_75t_L g684 ( 
.A(n_581),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_600),
.B(n_501),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_600),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_618),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_618),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_572),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_622),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_627),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_576),
.B(n_432),
.Y(n_692)
);

BUFx4f_ASAP7_75t_L g693 ( 
.A(n_641),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_603),
.B(n_628),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_571),
.A2(n_469),
.B1(n_458),
.B2(n_451),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_603),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_646),
.B(n_519),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_647),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_622),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_628),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_567),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_620),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_649),
.B(n_480),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_614),
.A2(n_469),
.B1(n_458),
.B2(n_434),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_623),
.B(n_480),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_623),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_616),
.B(n_509),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_624),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_624),
.B(n_481),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_593),
.B(n_443),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_632),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_585),
.B(n_602),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_625),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_616),
.B(n_615),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_644),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_620),
.Y(n_716)
);

AO21x2_ASAP7_75t_L g717 ( 
.A1(n_619),
.A2(n_423),
.B(n_507),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_625),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_629),
.Y(n_719)
);

INVx8_ASAP7_75t_L g720 ( 
.A(n_581),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_629),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_635),
.Y(n_722)
);

INVx1_ASAP7_75t_SL g723 ( 
.A(n_592),
.Y(n_723)
);

NOR2x1p5_ASAP7_75t_L g724 ( 
.A(n_605),
.B(n_410),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_567),
.Y(n_725)
);

NOR2x1p5_ASAP7_75t_L g726 ( 
.A(n_605),
.B(n_410),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_635),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_601),
.B(n_445),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_620),
.B(n_501),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_567),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_567),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_609),
.B(n_432),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_575),
.Y(n_733)
);

AND3x2_ASAP7_75t_L g734 ( 
.A(n_595),
.B(n_453),
.C(n_452),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_611),
.B(n_501),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_575),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_672),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_676),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_656),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_669),
.B(n_612),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_652),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_659),
.B(n_662),
.Y(n_742)
);

NAND2x1p5_ASAP7_75t_L g743 ( 
.A(n_674),
.B(n_696),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_657),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_659),
.B(n_619),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_658),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_661),
.B(n_612),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_664),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_679),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_682),
.B(n_710),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_662),
.B(n_714),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_691),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_698),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_689),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_653),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_663),
.Y(n_756)
);

NOR2x1p5_ASAP7_75t_L g757 ( 
.A(n_702),
.B(n_604),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_707),
.B(n_631),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_728),
.B(n_644),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_676),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_681),
.B(n_694),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_697),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_694),
.B(n_606),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_660),
.B(n_608),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_697),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_711),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_672),
.B(n_700),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_668),
.B(n_667),
.Y(n_768)
);

BUFx4_ASAP7_75t_L g769 ( 
.A(n_715),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_665),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_672),
.B(n_607),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_673),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_700),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_696),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_670),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_702),
.B(n_570),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_700),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_686),
.B(n_608),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_654),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_685),
.B(n_446),
.Y(n_780)
);

NAND3x1_ASAP7_75t_L g781 ( 
.A(n_668),
.B(n_454),
.C(n_447),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_716),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_667),
.B(n_631),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_680),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_713),
.B(n_588),
.Y(n_785)
);

OR2x6_ASAP7_75t_L g786 ( 
.A(n_684),
.B(n_607),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_680),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_685),
.B(n_446),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_692),
.B(n_588),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_678),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_683),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_701),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_687),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_688),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_690),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_699),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_706),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_L g798 ( 
.A(n_704),
.B(n_564),
.C(n_467),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_735),
.B(n_597),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_724),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_723),
.A2(n_671),
.B1(n_695),
.B2(n_675),
.Y(n_801)
);

OAI22xp33_ASAP7_75t_L g802 ( 
.A1(n_723),
.A2(n_564),
.B1(n_439),
.B2(n_432),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_716),
.B(n_570),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_666),
.A2(n_437),
.B1(n_439),
.B2(n_432),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_674),
.B(n_633),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_670),
.Y(n_806)
);

AO21x2_ASAP7_75t_L g807 ( 
.A1(n_717),
.A2(n_598),
.B(n_591),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_671),
.A2(n_469),
.B1(n_467),
.B2(n_458),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_674),
.B(n_729),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_729),
.B(n_633),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_735),
.B(n_455),
.Y(n_811)
);

INVx8_ASAP7_75t_L g812 ( 
.A(n_737),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_749),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_752),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_741),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_750),
.B(n_693),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_779),
.A2(n_732),
.B(n_712),
.C(n_225),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_781),
.A2(n_734),
.B1(n_197),
.B2(n_225),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_SL g819 ( 
.A1(n_747),
.A2(n_651),
.B1(n_455),
.B2(n_439),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_757),
.B(n_726),
.Y(n_820)
);

BUFx12f_ASAP7_75t_L g821 ( 
.A(n_754),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_742),
.B(n_651),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_740),
.B(n_778),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_751),
.B(n_708),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_739),
.B(n_718),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_768),
.B(n_719),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_800),
.B(n_693),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_760),
.B(n_721),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_744),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_746),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_748),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_745),
.B(n_722),
.Y(n_832)
);

AND3x2_ASAP7_75t_L g833 ( 
.A(n_759),
.B(n_441),
.C(n_727),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_761),
.B(n_763),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_738),
.B(n_650),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_753),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_737),
.B(n_439),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_764),
.B(n_655),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_738),
.B(n_650),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_784),
.B(n_787),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_798),
.A2(n_469),
.B1(n_655),
.B2(n_434),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_791),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_783),
.B(n_650),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_785),
.B(n_650),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_766),
.B(n_455),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_737),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_804),
.A2(n_655),
.B1(n_434),
.B2(n_439),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_773),
.B(n_455),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_758),
.B(n_789),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_794),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_780),
.B(n_455),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_801),
.A2(n_181),
.B1(n_222),
.B2(n_211),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_762),
.B(n_677),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_795),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_788),
.B(n_437),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_765),
.B(n_677),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_796),
.B(n_677),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_802),
.A2(n_720),
.B(n_684),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_773),
.B(n_437),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_773),
.B(n_736),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_797),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_769),
.Y(n_862)
);

NOR2xp67_ASAP7_75t_SL g863 ( 
.A(n_777),
.B(n_442),
.Y(n_863)
);

NAND3xp33_ASAP7_75t_L g864 ( 
.A(n_808),
.B(n_181),
.C(n_591),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_767),
.B(n_701),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_755),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_756),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_777),
.B(n_701),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_770),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_772),
.B(n_677),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_790),
.B(n_703),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_793),
.B(n_703),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_775),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_777),
.B(n_736),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_776),
.B(n_736),
.Y(n_875)
);

BUFx5_ASAP7_75t_L g876 ( 
.A(n_775),
.Y(n_876)
);

INVx8_ASAP7_75t_L g877 ( 
.A(n_776),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_771),
.B(n_705),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_811),
.B(n_725),
.Y(n_879)
);

OAI22xp33_ASAP7_75t_L g880 ( 
.A1(n_786),
.A2(n_720),
.B1(n_684),
.B2(n_598),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_799),
.B(n_705),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_810),
.B(n_725),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_774),
.B(n_709),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_803),
.B(n_733),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_782),
.B(n_709),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_810),
.B(n_725),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_792),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_803),
.B(n_733),
.Y(n_888)
);

NOR3xp33_ASAP7_75t_L g889 ( 
.A(n_809),
.B(n_509),
.C(n_638),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_806),
.B(n_597),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_849),
.B(n_806),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_880),
.A2(n_786),
.B1(n_805),
.B2(n_807),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_818),
.A2(n_805),
.B1(n_807),
.B2(n_720),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_820),
.B(n_743),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_817),
.A2(n_717),
.B(n_440),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_815),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_822),
.B(n_792),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_820),
.B(n_792),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_862),
.B(n_730),
.Y(n_899)
);

O2A1O1Ixp5_ASAP7_75t_L g900 ( 
.A1(n_816),
.A2(n_648),
.B(n_638),
.C(n_577),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_821),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_878),
.B(n_730),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_829),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_824),
.B(n_730),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_818),
.B(n_823),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_852),
.A2(n_582),
.B1(n_583),
.B2(n_580),
.Y(n_906)
);

BUFx8_ASAP7_75t_L g907 ( 
.A(n_846),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_830),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_840),
.B(n_731),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_881),
.B(n_731),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_836),
.B(n_731),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_883),
.B(n_733),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_838),
.A2(n_415),
.B1(n_581),
.B2(n_440),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_827),
.B(n_441),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_877),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_819),
.B(n_855),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_832),
.B(n_590),
.Y(n_917)
);

OAI22xp33_ASAP7_75t_L g918 ( 
.A1(n_864),
.A2(n_640),
.B1(n_645),
.B2(n_642),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_831),
.Y(n_919)
);

OAI21xp33_ASAP7_75t_L g920 ( 
.A1(n_843),
.A2(n_212),
.B(n_207),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_826),
.B(n_640),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_876),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_877),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_877),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_876),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_885),
.B(n_642),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_846),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_846),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_844),
.B(n_575),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_825),
.B(n_645),
.Y(n_930)
);

INVx5_ASAP7_75t_L g931 ( 
.A(n_812),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_889),
.B(n_575),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_851),
.B(n_584),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_834),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_845),
.B(n_584),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_865),
.B(n_648),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_812),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_859),
.A2(n_430),
.B(n_427),
.C(n_429),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_841),
.A2(n_581),
.B1(n_440),
.B2(n_438),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_833),
.B(n_216),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_873),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_858),
.A2(n_440),
.B(n_438),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_SL g943 ( 
.A1(n_847),
.A2(n_882),
.B1(n_886),
.B2(n_879),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_813),
.B(n_814),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_853),
.B(n_584),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_875),
.B(n_221),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_866),
.B(n_594),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_941),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_905),
.A2(n_848),
.B(n_835),
.C(n_839),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_L g950 ( 
.A1(n_893),
.A2(n_856),
.B(n_857),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_940),
.A2(n_863),
.B(n_888),
.C(n_884),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_895),
.A2(n_916),
.B(n_894),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_901),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_932),
.A2(n_837),
.B(n_870),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_909),
.B(n_891),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_900),
.A2(n_872),
.B(n_871),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_931),
.B(n_887),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_929),
.B(n_842),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_937),
.B(n_850),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_910),
.B(n_861),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_927),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_920),
.B(n_867),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_892),
.A2(n_828),
.B(n_854),
.Y(n_963)
);

NOR3xp33_ASAP7_75t_L g964 ( 
.A(n_946),
.B(n_874),
.C(n_860),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_944),
.Y(n_965)
);

AOI21x1_ASAP7_75t_L g966 ( 
.A1(n_899),
.A2(n_890),
.B(n_869),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_902),
.B(n_876),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_945),
.A2(n_868),
.B(n_515),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_896),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_908),
.B(n_876),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_927),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_898),
.A2(n_515),
.B(n_594),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_927),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_919),
.B(n_876),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_912),
.B(n_812),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_931),
.B(n_630),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_907),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_903),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_942),
.A2(n_438),
.B(n_584),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_918),
.A2(n_938),
.B(n_906),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_915),
.B(n_630),
.Y(n_981)
);

AO21x1_ASAP7_75t_L g982 ( 
.A1(n_897),
.A2(n_0),
.B(n_1),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_915),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_914),
.A2(n_470),
.B(n_215),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_947),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_906),
.A2(n_935),
.B(n_943),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_904),
.B(n_930),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_923),
.B(n_630),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_911),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_931),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_933),
.A2(n_427),
.B(n_429),
.C(n_424),
.Y(n_991)
);

BUFx4f_ASAP7_75t_L g992 ( 
.A(n_928),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_934),
.B(n_630),
.Y(n_993)
);

AOI21xp33_ASAP7_75t_L g994 ( 
.A1(n_926),
.A2(n_0),
.B(n_1),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_917),
.A2(n_470),
.B(n_217),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_913),
.A2(n_430),
.B1(n_424),
.B2(n_425),
.Y(n_996)
);

NOR2xp67_ASAP7_75t_L g997 ( 
.A(n_924),
.B(n_2),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_928),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_921),
.B(n_3),
.Y(n_999)
);

CKINVDCx10_ASAP7_75t_R g1000 ( 
.A(n_907),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_947),
.B(n_3),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_922),
.B(n_470),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_925),
.Y(n_1003)
);

OAI21xp33_ASAP7_75t_L g1004 ( 
.A1(n_939),
.A2(n_219),
.B(n_214),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_936),
.B(n_4),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_895),
.A2(n_470),
.B(n_409),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_893),
.A2(n_496),
.B1(n_481),
.B2(n_485),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_905),
.A2(n_472),
.B(n_468),
.C(n_460),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_909),
.B(n_4),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_909),
.B(n_5),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_893),
.A2(n_409),
.B1(n_499),
.B2(n_490),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_894),
.B(n_5),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_893),
.A2(n_485),
.B1(n_491),
.B2(n_495),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_1000),
.B(n_6),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_948),
.Y(n_1015)
);

NAND2x1p5_ASAP7_75t_L g1016 ( 
.A(n_957),
.B(n_493),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_952),
.A2(n_220),
.B(n_224),
.C(n_226),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_986),
.A2(n_431),
.B1(n_411),
.B2(n_418),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_1011),
.A2(n_951),
.B1(n_980),
.B2(n_1012),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_977),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_953),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_985),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_963),
.A2(n_994),
.B(n_982),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_984),
.A2(n_409),
.B(n_417),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_949),
.A2(n_418),
.B(n_417),
.Y(n_1025)
);

BUFx4f_ASAP7_75t_L g1026 ( 
.A(n_990),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_1012),
.A2(n_431),
.B1(n_405),
.B2(n_413),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_990),
.B(n_992),
.Y(n_1028)
);

CKINVDCx8_ASAP7_75t_R g1029 ( 
.A(n_990),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_998),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_965),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1020),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1015),
.Y(n_1033)
);

INVx4_ASAP7_75t_L g1034 ( 
.A(n_1026),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1023),
.B(n_950),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_1019),
.B(n_1029),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_1031),
.B(n_955),
.Y(n_1037)
);

OAI21xp33_ASAP7_75t_SL g1038 ( 
.A1(n_1028),
.A2(n_1030),
.B(n_1022),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1018),
.B(n_956),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1027),
.B(n_1001),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1017),
.B(n_989),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1026),
.B(n_1009),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_1014),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_1016),
.A2(n_1007),
.B1(n_1013),
.B2(n_964),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1025),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1024),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_SL g1047 ( 
.A1(n_1021),
.A2(n_1005),
.B1(n_962),
.B2(n_1006),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_1021),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1023),
.B(n_1010),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1023),
.A2(n_983),
.B1(n_997),
.B2(n_971),
.Y(n_1050)
);

O2A1O1Ixp5_ASAP7_75t_L g1051 ( 
.A1(n_1023),
.A2(n_976),
.B(n_954),
.C(n_966),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1015),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1023),
.B(n_999),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_1026),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1015),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_1029),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1056),
.B(n_998),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1043),
.B(n_959),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1033),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_1035),
.A2(n_1003),
.A3(n_969),
.B(n_978),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_1043),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_1043),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_SL g1063 ( 
.A1(n_1050),
.A2(n_1049),
.B(n_1053),
.C(n_1036),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1063),
.A2(n_1038),
.B(n_1039),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_1061),
.A2(n_1051),
.B(n_1047),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_1062),
.B(n_1032),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_1066),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1065),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_1064),
.A2(n_1057),
.B(n_1059),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1069),
.A2(n_1058),
.B(n_1055),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_1067),
.B(n_1034),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_1071),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1071),
.A2(n_1068),
.B1(n_1067),
.B2(n_1069),
.Y(n_1073)
);

AO31x2_ASAP7_75t_L g1074 ( 
.A1(n_1072),
.A2(n_1068),
.A3(n_1070),
.B(n_1067),
.Y(n_1074)
);

AO21x2_ASAP7_75t_L g1075 ( 
.A1(n_1073),
.A2(n_1070),
.B(n_1042),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_1075),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1075),
.B(n_1034),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1077),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1076),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1079),
.A2(n_1076),
.B(n_1074),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1078),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_SL g1082 ( 
.A1(n_1081),
.A2(n_1054),
.B1(n_1048),
.B2(n_1074),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1080),
.A2(n_1054),
.B1(n_1045),
.B2(n_1046),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1081),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_1084),
.B(n_1054),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_1082),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1083),
.B(n_1060),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_1085),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1085),
.Y(n_1089)
);

AOI221xp5_ASAP7_75t_L g1090 ( 
.A1(n_1088),
.A2(n_1086),
.B1(n_1087),
.B2(n_1052),
.C(n_1041),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_L g1091 ( 
.A(n_1089),
.B(n_1086),
.C(n_1040),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1091),
.A2(n_961),
.B1(n_973),
.B2(n_1037),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1090),
.Y(n_1093)
);

INVxp67_ASAP7_75t_SL g1094 ( 
.A(n_1093),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1092),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_1095),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_SL g1097 ( 
.A(n_1094),
.B(n_7),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1096),
.B(n_7),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1097),
.B(n_1060),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1098),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1099),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_1099),
.B(n_1060),
.Y(n_1102)
);

AOI222xp33_ASAP7_75t_L g1103 ( 
.A1(n_1101),
.A2(n_973),
.B1(n_961),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1102),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1100),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_1105),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1104),
.B(n_1044),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_1106),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_1107),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1108),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1109),
.B(n_1103),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1110),
.B(n_998),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1111),
.B(n_8),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1112),
.B(n_975),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_SL g1115 ( 
.A(n_1113),
.B(n_9),
.C(n_10),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1115),
.A2(n_11),
.B(n_12),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1114),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1116),
.B(n_13),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1117),
.B(n_16),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1116),
.B(n_16),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1120),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_17),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1118),
.Y(n_1123)
);

AOI221xp5_ASAP7_75t_L g1124 ( 
.A1(n_1123),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.C(n_21),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1121),
.B(n_18),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1124),
.A2(n_1122),
.B1(n_22),
.B2(n_23),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1125),
.Y(n_1127)
);

AOI221xp5_ASAP7_75t_L g1128 ( 
.A1(n_1127),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.C(n_24),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_SL g1129 ( 
.A(n_1126),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_1129),
.B(n_24),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1128),
.A2(n_25),
.B(n_26),
.Y(n_1131)
);

OAI31xp33_ASAP7_75t_L g1132 ( 
.A1(n_1131),
.A2(n_27),
.A3(n_28),
.B(n_29),
.Y(n_1132)
);

AOI221xp5_ASAP7_75t_L g1133 ( 
.A1(n_1130),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.C(n_30),
.Y(n_1133)
);

NOR3xp33_ASAP7_75t_SL g1134 ( 
.A(n_1132),
.B(n_30),
.C(n_31),
.Y(n_1134)
);

OAI221xp5_ASAP7_75t_L g1135 ( 
.A1(n_1133),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.C(n_36),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1134),
.B(n_37),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_1135),
.B(n_38),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_L g1138 ( 
.A(n_1134),
.B(n_1008),
.C(n_39),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1136),
.Y(n_1139)
);

NAND4xp75_ASAP7_75t_L g1140 ( 
.A(n_1137),
.B(n_1138),
.C(n_42),
.D(n_43),
.Y(n_1140)
);

NOR2x1_ASAP7_75t_L g1141 ( 
.A(n_1137),
.B(n_40),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1139),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1141),
.B(n_1140),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1142),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1143),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1144),
.B(n_44),
.Y(n_1146)
);

NAND4xp75_ASAP7_75t_L g1147 ( 
.A(n_1145),
.B(n_45),
.C(n_46),
.D(n_47),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1147),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_1148)
);

NOR4xp75_ASAP7_75t_L g1149 ( 
.A(n_1146),
.B(n_52),
.C(n_53),
.D(n_54),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_SL g1150 ( 
.A1(n_1148),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1150)
);

OAI221xp5_ASAP7_75t_L g1151 ( 
.A1(n_1149),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.C(n_65),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_SL g1152 ( 
.A(n_1151),
.B(n_66),
.C(n_67),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1150),
.Y(n_1153)
);

OAI211xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1153),
.A2(n_68),
.B(n_69),
.C(n_71),
.Y(n_1154)
);

XNOR2x1_ASAP7_75t_L g1155 ( 
.A(n_1152),
.B(n_72),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1153),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1156),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1155),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_1154),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1157),
.B(n_74),
.Y(n_1160)
);

XNOR2x1_ASAP7_75t_L g1161 ( 
.A(n_1158),
.B(n_1159),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1161),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1160),
.Y(n_1163)
);

AOI22x1_ASAP7_75t_L g1164 ( 
.A1(n_1162),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1163),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1164),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1165),
.Y(n_1167)
);

NAND4xp25_ASAP7_75t_L g1168 ( 
.A(n_1167),
.B(n_83),
.C(n_84),
.D(n_86),
.Y(n_1168)
);

OAI31xp33_ASAP7_75t_L g1169 ( 
.A1(n_1166),
.A2(n_87),
.A3(n_88),
.B(n_91),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1169),
.Y(n_1170)
);

OAI22x1_ASAP7_75t_L g1171 ( 
.A1(n_1168),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1170),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1171),
.Y(n_1173)
);

XNOR2xp5_ASAP7_75t_L g1174 ( 
.A(n_1170),
.B(n_96),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1170),
.B(n_97),
.Y(n_1175)
);

OAI22x1_ASAP7_75t_L g1176 ( 
.A1(n_1172),
.A2(n_489),
.B1(n_981),
.B2(n_105),
.Y(n_1176)
);

NAND3xp33_ASAP7_75t_SL g1177 ( 
.A(n_1173),
.B(n_103),
.C(n_104),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1175),
.Y(n_1178)
);

OAI22x1_ASAP7_75t_L g1179 ( 
.A1(n_1174),
.A2(n_489),
.B1(n_981),
.B2(n_111),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_1178),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_SL g1181 ( 
.A1(n_1179),
.A2(n_1176),
.B1(n_1177),
.B2(n_489),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1178),
.A2(n_106),
.B(n_109),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1180),
.A2(n_988),
.B1(n_419),
.B2(n_412),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1181),
.A2(n_112),
.B(n_113),
.Y(n_1184)
);

AOI21xp33_ASAP7_75t_SL g1185 ( 
.A1(n_1182),
.A2(n_116),
.B(n_117),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1180),
.A2(n_118),
.B(n_119),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1180),
.B(n_120),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1180),
.B(n_121),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1180),
.A2(n_122),
.B(n_123),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1180),
.A2(n_988),
.B1(n_126),
.B2(n_127),
.Y(n_1190)
);

AOI222xp33_ASAP7_75t_L g1191 ( 
.A1(n_1180),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.C1(n_132),
.C2(n_134),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1180),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_1192)
);

AOI222xp33_ASAP7_75t_L g1193 ( 
.A1(n_1180),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.C1(n_143),
.C2(n_145),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1180),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1194),
.B(n_150),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1185),
.A2(n_1187),
.B(n_1184),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1187),
.A2(n_1190),
.B(n_1189),
.Y(n_1197)
);

AOI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1188),
.A2(n_151),
.B(n_152),
.Y(n_1198)
);

NOR2x1_ASAP7_75t_L g1199 ( 
.A(n_1186),
.B(n_153),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1191),
.B(n_154),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1193),
.Y(n_1201)
);

XNOR2xp5_ASAP7_75t_L g1202 ( 
.A(n_1192),
.B(n_155),
.Y(n_1202)
);

NOR2x1_ASAP7_75t_L g1203 ( 
.A(n_1183),
.B(n_159),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1201),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1196),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_1205)
);

INVxp67_ASAP7_75t_SL g1206 ( 
.A(n_1197),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1200),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1202),
.Y(n_1208)
);

XNOR2xp5_ASAP7_75t_L g1209 ( 
.A(n_1199),
.B(n_165),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1203),
.B(n_166),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1204),
.A2(n_1206),
.B1(n_1208),
.B2(n_1207),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1210),
.B(n_1198),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1209),
.A2(n_1195),
.B(n_168),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1211),
.A2(n_1205),
.B(n_170),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1214),
.A2(n_1212),
.B1(n_1213),
.B2(n_173),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1215),
.A2(n_167),
.B1(n_172),
.B2(n_174),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1216),
.B(n_968),
.Y(n_1217)
);

OAI221xp5_ASAP7_75t_R g1218 ( 
.A1(n_1217),
.A2(n_993),
.B1(n_972),
.B2(n_974),
.C(n_970),
.Y(n_1218)
);

AOI221xp5_ASAP7_75t_L g1219 ( 
.A1(n_1218),
.A2(n_958),
.B1(n_967),
.B2(n_960),
.C(n_987),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1219),
.A2(n_1004),
.B1(n_1002),
.B2(n_996),
.Y(n_1220)
);

OAI31xp33_ASAP7_75t_L g1221 ( 
.A1(n_1220),
.A2(n_979),
.A3(n_991),
.B(n_995),
.Y(n_1221)
);

AOI211xp5_ASAP7_75t_L g1222 ( 
.A1(n_1221),
.A2(n_522),
.B(n_493),
.C(n_521),
.Y(n_1222)
);


endmodule