module fake_jpeg_12598_n_263 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_263);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_49),
.Y(n_88)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_63),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_58),
.Y(n_101)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_62),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_65),
.B(n_73),
.Y(n_119)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_16),
.B(n_14),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_72),
.Y(n_85)
);

CKINVDCx9p33_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_68),
.Y(n_100)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_75),
.Y(n_99)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_2),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_77),
.Y(n_117)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_79),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_82),
.Y(n_122)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

CKINVDCx11_ASAP7_75t_R g111 ( 
.A(n_81),
.Y(n_111)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_12),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_48),
.A2(n_43),
.B1(n_19),
.B2(n_26),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_94),
.A2(n_96),
.B1(n_112),
.B2(n_118),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_46),
.A2(n_18),
.B1(n_33),
.B2(n_28),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_40),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_71),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_18),
.B1(n_40),
.B2(n_39),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_114),
.B1(n_115),
.B2(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_50),
.A2(n_70),
.B1(n_75),
.B2(n_74),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_62),
.A2(n_39),
.B1(n_43),
.B2(n_38),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_60),
.A2(n_19),
.B1(n_36),
.B2(n_33),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_38),
.B1(n_36),
.B2(n_28),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_45),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_69),
.A2(n_23),
.B1(n_21),
.B2(n_5),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_66),
.B1(n_58),
.B2(n_47),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_95),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_2),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_127),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_56),
.A2(n_61),
.B1(n_51),
.B2(n_52),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_54),
.B(n_4),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_99),
.Y(n_160)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_132),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_131),
.B(n_137),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_88),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_91),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_135),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_117),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx2_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_6),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_142),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_158),
.B1(n_162),
.B2(n_101),
.Y(n_164)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_7),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_7),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_143),
.B(n_146),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_100),
.A2(n_81),
.B1(n_55),
.B2(n_58),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_151),
.B1(n_161),
.B2(n_106),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_8),
.Y(n_146)
);

INVx6_ASAP7_75t_SL g147 ( 
.A(n_111),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_147),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_8),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_153),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_87),
.B(n_103),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_155),
.Y(n_185)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_11),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_157),
.C(n_159),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_99),
.B(n_11),
.C(n_102),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_99),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_156),
.C(n_138),
.Y(n_175)
);

BUFx4f_ASAP7_75t_SL g161 ( 
.A(n_93),
.Y(n_161)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_159),
.A2(n_144),
.B1(n_129),
.B2(n_135),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_167),
.B1(n_177),
.B2(n_184),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_164),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_112),
.B1(n_92),
.B2(n_97),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_92),
.B1(n_89),
.B2(n_97),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_181),
.B1(n_147),
.B2(n_162),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_172),
.A2(n_171),
.B1(n_184),
.B2(n_167),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_152),
.C(n_141),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_149),
.A2(n_89),
.B1(n_126),
.B2(n_93),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_126),
.B1(n_113),
.B2(n_101),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_142),
.A2(n_113),
.B1(n_106),
.B2(n_98),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_154),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_191),
.B(n_193),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_137),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_196),
.C(n_175),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_180),
.B(n_108),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_197),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_98),
.C(n_108),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_84),
.B(n_140),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_179),
.B(n_140),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_202),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_199),
.A2(n_192),
.B1(n_181),
.B2(n_168),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_140),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_177),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_161),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_136),
.B1(n_155),
.B2(n_86),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_204),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_170),
.A2(n_86),
.B1(n_123),
.B2(n_116),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_201),
.B1(n_198),
.B2(n_203),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_215),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_186),
.B(n_171),
.C(n_173),
.Y(n_213)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_194),
.C(n_190),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_176),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_178),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_217),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_189),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_192),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_227),
.C(n_230),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_221),
.A2(n_219),
.B1(n_217),
.B2(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_225),
.B(n_231),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_178),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_229),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_187),
.C(n_204),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_183),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_201),
.C(n_174),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_174),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_205),
.B(n_206),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_219),
.B1(n_210),
.B2(n_218),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_238),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_211),
.C(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_228),
.B(n_211),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_223),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_191),
.B1(n_166),
.B2(n_182),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_220),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_246),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_230),
.C(n_231),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_241),
.C(n_237),
.Y(n_248)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_243),
.B(n_244),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_248),
.B(n_249),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_235),
.C(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_234),
.C(n_232),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_169),
.C(n_166),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_252),
.A2(n_247),
.B1(n_245),
.B2(n_240),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_250),
.C(n_169),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_252),
.B(n_183),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_253),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);

NOR3xp33_ASAP7_75t_SL g259 ( 
.A(n_258),
.B(n_84),
.C(n_161),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_165),
.C(n_133),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_260),
.B(n_116),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_95),
.Y(n_263)
);


endmodule