module fake_jpeg_9661_n_102 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_SL g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_64),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_68),
.Y(n_77)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_7),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_8),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_9),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_62),
.B1(n_59),
.B2(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_11),
.B1(n_14),
.B2(n_18),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_58),
.B1(n_61),
.B2(n_52),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_49),
.B1(n_54),
.B2(n_16),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_79),
.B(n_81),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_86),
.B(n_87),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_88),
.B1(n_83),
.B2(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_91),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_77),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_78),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_90),
.C(n_23),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_41),
.Y(n_96)
);

OAI221xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_19),
.B1(n_25),
.B2(n_27),
.C(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_29),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_30),
.B(n_31),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_32),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_33),
.B(n_36),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_37),
.Y(n_102)
);


endmodule