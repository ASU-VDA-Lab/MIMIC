module fake_jpeg_28133_n_294 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.Y(n_45)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_54),
.A2(n_60),
.B1(n_41),
.B2(n_37),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_26),
.B1(n_18),
.B2(n_32),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_55),
.A2(n_63),
.B1(n_25),
.B2(n_30),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_32),
.B1(n_26),
.B2(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_41),
.B1(n_40),
.B2(n_43),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_66),
.A2(n_36),
.B1(n_28),
.B2(n_25),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_69),
.B(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_72),
.B(n_74),
.Y(n_111)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_42),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_22),
.B1(n_41),
.B2(n_44),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_75),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_80),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_44),
.B(n_43),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_79),
.A2(n_89),
.B(n_36),
.C(n_28),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_33),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx2_ASAP7_75t_SL g105 ( 
.A(n_81),
.Y(n_105)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_35),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_88),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_43),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_56),
.B(n_21),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_0),
.B(n_33),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_91),
.Y(n_108)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

NAND2x1_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_41),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_31),
.C(n_23),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_97),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_49),
.A2(n_21),
.B(n_31),
.C(n_17),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_10),
.C(n_1),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_35),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_17),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_36),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_30),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_45),
.B(n_30),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_24),
.Y(n_129)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_79),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_94),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_117),
.B1(n_123),
.B2(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_115),
.B(n_119),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_81),
.B1(n_1),
.B2(n_2),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_127),
.A2(n_75),
.B1(n_80),
.B2(n_102),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_144),
.B1(n_154),
.B2(n_110),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_120),
.B(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_73),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_93),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_76),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_129),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_99),
.C(n_95),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_151),
.C(n_125),
.Y(n_162)
);

AO21x2_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_97),
.B(n_100),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_153),
.B1(n_124),
.B2(n_117),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_101),
.B1(n_97),
.B2(n_84),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_156),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_91),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_71),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_71),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_149),
.B(n_152),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_67),
.C(n_82),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_84),
.B1(n_68),
.B2(n_86),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_68),
.B1(n_86),
.B2(n_23),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_83),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_23),
.Y(n_157)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_112),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_125),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_21),
.B(n_31),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_162),
.B(n_165),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_163),
.A2(n_166),
.B1(n_176),
.B2(n_181),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_151),
.C(n_156),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_171),
.C(n_183),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_143),
.B1(n_134),
.B2(n_149),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_180),
.B1(n_155),
.B2(n_139),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_173),
.B(n_182),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_129),
.B1(n_120),
.B2(n_121),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_184),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_104),
.B1(n_121),
.B2(n_131),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_131),
.B1(n_24),
.B2(n_31),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_112),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_143),
.A2(n_36),
.B1(n_0),
.B2(n_2),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_150),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_153),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_137),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_139),
.A2(n_3),
.B(n_4),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_145),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_199),
.B(n_204),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_141),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_203),
.B1(n_207),
.B2(n_213),
.Y(n_221)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_174),
.Y(n_202)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_133),
.Y(n_205)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_190),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_206),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_169),
.A2(n_144),
.B1(n_152),
.B2(n_135),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_142),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_211),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_178),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_170),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_163),
.A2(n_132),
.B1(n_6),
.B2(n_7),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_16),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_188),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_215),
.B(n_213),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_171),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_230),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_209),
.B(n_162),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_224),
.B(n_231),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_176),
.C(n_166),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_229),
.C(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

AOI22x1_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_186),
.B1(n_177),
.B2(n_172),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_197),
.B1(n_207),
.B2(n_193),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_168),
.C(n_170),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_5),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_5),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_6),
.B(n_7),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_203),
.B(n_9),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_225),
.A2(n_198),
.B1(n_194),
.B2(n_205),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_239),
.B1(n_230),
.B2(n_191),
.Y(n_260)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_237),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_218),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_228),
.A2(n_198),
.B1(n_202),
.B2(n_210),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_240),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_233),
.B1(n_220),
.B2(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_215),
.Y(n_258)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_246),
.A2(n_247),
.B(n_248),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_249),
.A2(n_191),
.B(n_195),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_216),
.B(n_222),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_260),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_222),
.B(n_212),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_255),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_257),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_224),
.C(n_236),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_234),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_263),
.B(n_264),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_236),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_247),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_268),
.Y(n_279)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_238),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_270),
.B(n_267),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_238),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_219),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_261),
.Y(n_273)
);

FAx1_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_231),
.CI(n_232),
.CON(n_282),
.SN(n_282)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_266),
.A2(n_253),
.B(n_248),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_276),
.B(n_265),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_254),
.C(n_250),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_256),
.B1(n_246),
.B2(n_251),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_232),
.B1(n_201),
.B2(n_196),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_278),
.A2(n_271),
.B(n_252),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_282),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_281),
.B(n_283),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_214),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_277),
.B1(n_196),
.B2(n_201),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_276),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

OAI311xp33_ASAP7_75t_L g290 ( 
.A1(n_288),
.A2(n_289),
.A3(n_285),
.B1(n_273),
.C1(n_274),
.Y(n_290)
);

OAI321xp33_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_196),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C(n_14),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_8),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_10),
.B(n_11),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_15),
.Y(n_294)
);


endmodule