module fake_aes_3336_n_30 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
OA21x2_ASAP7_75t_L g12 ( .A1(n_4), .A2(n_2), .B(n_5), .Y(n_12) );
BUFx3_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
OAI22xp5_ASAP7_75t_L g14 ( .A1(n_9), .A2(n_3), .B1(n_6), .B2(n_0), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_10), .B(n_0), .Y(n_16) );
AND2x2_ASAP7_75t_SL g17 ( .A(n_16), .B(n_11), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_15), .B(n_1), .Y(n_18) );
OAI21x1_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_12), .B(n_14), .Y(n_19) );
OA21x2_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_16), .B(n_15), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_19), .B(n_18), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_17), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_17), .Y(n_23) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_23), .Y(n_24) );
AOI21xp5_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_20), .B(n_18), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_12), .Y(n_26) );
NOR2x1_ASAP7_75t_L g27 ( .A(n_25), .B(n_12), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_27), .B1(n_13), .B2(n_20), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_13), .B1(n_2), .B2(n_7), .Y(n_30) );
endmodule