module fake_jpeg_22858_n_124 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_124);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_28),
.B1(n_17),
.B2(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_30),
.B(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_32),
.B(n_37),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_22),
.B(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g39 ( 
.A1(n_22),
.A2(n_4),
.B(n_5),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_15),
.B1(n_20),
.B2(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_7),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_50),
.B1(n_58),
.B2(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_49),
.B(n_52),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_19),
.B1(n_20),
.B2(n_15),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_17),
.Y(n_57)
);

AND2x4_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_21),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_57),
.B(n_44),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_21),
.B1(n_27),
.B2(n_11),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_7),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_63),
.B(n_10),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_35),
.B1(n_40),
.B2(n_13),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_71),
.C(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_59),
.B1(n_47),
.B2(n_62),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_76),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_62),
.C(n_44),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_49),
.B1(n_48),
.B2(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_85),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_68),
.C(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_53),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_43),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_68),
.C(n_73),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_102),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_91),
.A2(n_69),
.B1(n_70),
.B2(n_43),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_101),
.B1(n_92),
.B2(n_99),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_72),
.B1(n_69),
.B2(n_54),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_87),
.B1(n_85),
.B2(n_90),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_79),
.B(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_65),
.B(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_95),
.B1(n_98),
.B2(n_108),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_93),
.B1(n_99),
.B2(n_101),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

AO221x1_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_96),
.B1(n_103),
.B2(n_83),
.C(n_21),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_89),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_107),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_113),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_95),
.B1(n_97),
.B2(n_100),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_103),
.C(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_110),
.B(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_114),
.B(n_115),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_120),
.C(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_106),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_122),
.Y(n_124)
);


endmodule