module real_jpeg_13903_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_3),
.A2(n_18),
.B1(n_20),
.B2(n_28),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_3),
.A2(n_5),
.B(n_22),
.C(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_3),
.B(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_3),
.B(n_34),
.C(n_36),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_3),
.B(n_17),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

AO22x1_ASAP7_75t_L g17 ( 
.A1(n_5),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_17)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_7),
.A2(n_18),
.B1(n_20),
.B2(n_25),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_7),
.A2(n_25),
.B1(n_35),
.B2(n_36),
.Y(n_72)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_84),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_83),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_57),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_13),
.B(n_57),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_31),
.C(n_46),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_14),
.A2(n_15),
.B1(n_31),
.B2(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_21),
.B(n_26),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_16),
.A2(n_21),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_19),
.B(n_23),
.C(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_18),
.A2(n_20),
.B1(n_34),
.B2(n_39),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_18),
.A2(n_19),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_20),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_22),
.A2(n_23),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_28),
.B(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_28),
.B(n_32),
.Y(n_107)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_31),
.B(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_31),
.A2(n_88),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_31),
.Y(n_101)
);

OA21x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_40),
.B(n_42),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2x1_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_45),
.Y(n_44)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_33),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_80)
);

AO22x1_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_33)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_35),
.B(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_46),
.A2(n_47),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_55),
.B1(n_56),
.B2(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_72),
.B(n_73),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_77),
.B2(n_78),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_75),
.B2(n_76),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_70),
.B2(n_71),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_70),
.B(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_71),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_82),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_93),
.C(n_95),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_111),
.B(n_116),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_97),
.B(n_110),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_90),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_90)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_92),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_107),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B(n_109),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B(n_108),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_112),
.B(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);


endmodule