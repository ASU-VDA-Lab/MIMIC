module fake_jpeg_26435_n_102 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_0),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_25),
.Y(n_30)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_28),
.Y(n_32)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_38),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_18),
.B1(n_20),
.B2(n_12),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_25),
.B1(n_17),
.B2(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_11),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_18),
.C(n_15),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_22),
.A2(n_21),
.B1(n_15),
.B2(n_13),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_13),
.B1(n_23),
.B2(n_26),
.Y(n_42)
);

NOR3xp33_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_11),
.C(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_37),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_44),
.Y(n_53)
);

AOI32xp33_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_27),
.A3(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_48),
.B(n_34),
.C(n_29),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_47),
.B1(n_32),
.B2(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_49),
.Y(n_58)
);

NAND2x1_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_55),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_46),
.B(n_43),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_60),
.B1(n_48),
.B2(n_35),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_34),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_36),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_53),
.Y(n_76)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_55),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_35),
.B1(n_36),
.B2(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_58),
.B(n_53),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_75),
.B(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_63),
.C(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_1),
.B(n_2),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_65),
.C(n_63),
.Y(n_81)
);

AOI221xp5_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_70),
.B1(n_7),
.B2(n_5),
.C(n_8),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_74),
.B(n_79),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_4),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_2),
.Y(n_92)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_9),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_93),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_8),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_89),
.C(n_88),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_95),
.B(n_9),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_10),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_94),
.C(n_88),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_99),
.A2(n_100),
.B(n_96),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_4),
.Y(n_102)
);


endmodule