module real_aes_7812_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_0), .A2(n_212), .B(n_216), .C(n_253), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_1), .A2(n_207), .B(n_276), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_3), .B(n_230), .Y(n_283) );
INVx1_ASAP7_75t_L g190 ( .A(n_4), .Y(n_190) );
AND2x6_ASAP7_75t_L g212 ( .A(n_4), .B(n_188), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_4), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g240 ( .A(n_5), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_6), .B(n_221), .Y(n_257) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_7), .A2(n_24), .B1(n_89), .B2(n_90), .Y(n_88) );
INVx1_ASAP7_75t_L g205 ( .A(n_8), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_9), .A2(n_241), .B(n_266), .C(n_268), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_10), .B(n_230), .Y(n_269) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_11), .A2(n_26), .B1(n_89), .B2(n_93), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_12), .B(n_325), .Y(n_324) );
OAI22xp5_ASAP7_75t_SL g169 ( .A1(n_13), .A2(n_170), .B1(n_171), .B2(n_177), .Y(n_169) );
INVx1_ASAP7_75t_L g177 ( .A(n_13), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_14), .A2(n_220), .B(n_222), .C(n_226), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_15), .B(n_221), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_16), .B(n_221), .Y(n_301) );
CKINVDCx16_ASAP7_75t_R g286 ( .A(n_17), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_18), .A2(n_80), .B1(n_167), .B2(n_168), .Y(n_79) );
INVx1_ASAP7_75t_L g167 ( .A(n_18), .Y(n_167) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_19), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_20), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_21), .Y(n_122) );
INVx1_ASAP7_75t_L g322 ( .A(n_22), .Y(n_322) );
INVx2_ASAP7_75t_L g210 ( .A(n_23), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_25), .Y(n_260) );
OAI221xp5_ASAP7_75t_L g181 ( .A1(n_26), .A2(n_40), .B1(n_51), .B2(n_182), .C(n_183), .Y(n_181) );
INVxp67_ASAP7_75t_L g184 ( .A(n_26), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_27), .A2(n_220), .B(n_279), .C(n_281), .Y(n_278) );
AOI22xp5_ASAP7_75t_SL g500 ( .A1(n_27), .A2(n_80), .B1(n_168), .B2(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_27), .Y(n_501) );
INVxp67_ASAP7_75t_L g323 ( .A(n_28), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_29), .A2(n_54), .B1(n_112), .B2(n_118), .Y(n_111) );
CKINVDCx14_ASAP7_75t_R g277 ( .A(n_30), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_31), .A2(n_216), .B(n_299), .C(n_304), .Y(n_298) );
AOI22xp33_ASAP7_75t_SL g159 ( .A1(n_32), .A2(n_70), .B1(n_160), .B2(n_163), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_33), .A2(n_238), .B(n_239), .C(n_242), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_34), .A2(n_62), .B1(n_146), .B2(n_150), .Y(n_145) );
AOI22xp33_ASAP7_75t_SL g154 ( .A1(n_35), .A2(n_69), .B1(n_155), .B2(n_157), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_36), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_37), .Y(n_319) );
AOI22xp33_ASAP7_75t_SL g135 ( .A1(n_38), .A2(n_42), .B1(n_136), .B2(n_141), .Y(n_135) );
INVx1_ASAP7_75t_L g214 ( .A(n_39), .Y(n_214) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_40), .A2(n_66), .B1(n_89), .B2(n_93), .Y(n_98) );
INVxp67_ASAP7_75t_L g185 ( .A(n_40), .Y(n_185) );
CKINVDCx14_ASAP7_75t_R g236 ( .A(n_41), .Y(n_236) );
INVx1_ASAP7_75t_L g188 ( .A(n_43), .Y(n_188) );
INVx1_ASAP7_75t_L g204 ( .A(n_44), .Y(n_204) );
INVx1_ASAP7_75t_SL g280 ( .A(n_45), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_46), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_47), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_48), .B(n_230), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_49), .A2(n_80), .B1(n_168), .B2(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_49), .Y(n_511) );
INVx1_ASAP7_75t_L g289 ( .A(n_50), .Y(n_289) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_51), .A2(n_72), .B1(n_89), .B2(n_90), .Y(n_96) );
OAI22xp5_ASAP7_75t_SL g174 ( .A1(n_52), .A2(n_63), .B1(n_175), .B2(n_176), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_52), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_53), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_55), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_56), .A2(n_207), .B(n_235), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_57), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_58), .A2(n_207), .B(n_263), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_59), .A2(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g264 ( .A(n_60), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g297 ( .A(n_61), .Y(n_297) );
INVx1_ASAP7_75t_L g176 ( .A(n_63), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_64), .A2(n_207), .B(n_213), .Y(n_206) );
INVx1_ASAP7_75t_L g267 ( .A(n_65), .Y(n_267) );
INVx2_ASAP7_75t_L g202 ( .A(n_67), .Y(n_202) );
INVx1_ASAP7_75t_L g254 ( .A(n_68), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g287 ( .A1(n_71), .A2(n_216), .B(n_288), .C(n_291), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_73), .B(n_200), .Y(n_244) );
INVx1_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_75), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_75), .Y(n_172) );
INVx2_ASAP7_75t_L g223 ( .A(n_76), .Y(n_223) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_178), .B1(n_191), .B2(n_496), .C(n_499), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_169), .Y(n_78) );
INVx2_ASAP7_75t_L g168 ( .A(n_80), .Y(n_168) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_133), .Y(n_80) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_104), .C(n_121), .Y(n_81) );
OAI22xp5_ASAP7_75t_L g82 ( .A1(n_83), .A2(n_84), .B1(n_99), .B2(n_100), .Y(n_82) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
OR2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_94), .Y(n_85) );
INVx2_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
OR2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
AND2x2_ASAP7_75t_L g103 ( .A(n_87), .B(n_92), .Y(n_103) );
AND2x2_ASAP7_75t_L g140 ( .A(n_87), .B(n_116), .Y(n_140) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g107 ( .A(n_88), .B(n_92), .Y(n_107) );
AND2x2_ASAP7_75t_L g117 ( .A(n_88), .B(n_98), .Y(n_117) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g93 ( .A(n_91), .Y(n_93) );
INVx2_ASAP7_75t_L g116 ( .A(n_92), .Y(n_116) );
INVx1_ASAP7_75t_L g166 ( .A(n_92), .Y(n_166) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NAND2x1p5_ASAP7_75t_L g102 ( .A(n_95), .B(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g158 ( .A(n_95), .B(n_140), .Y(n_158) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_97), .Y(n_95) );
INVx1_ASAP7_75t_L g109 ( .A(n_96), .Y(n_109) );
INVx1_ASAP7_75t_L g115 ( .A(n_96), .Y(n_115) );
INVx1_ASAP7_75t_L g132 ( .A(n_96), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_96), .B(n_98), .Y(n_144) );
AND2x2_ASAP7_75t_L g108 ( .A(n_97), .B(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g139 ( .A(n_98), .B(n_132), .Y(n_139) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x4_ASAP7_75t_L g152 ( .A(n_103), .B(n_108), .Y(n_152) );
AND2x2_ASAP7_75t_L g162 ( .A(n_103), .B(n_139), .Y(n_162) );
OAI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_110), .B(n_111), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AND2x6_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g129 ( .A(n_107), .Y(n_129) );
AND2x6_ASAP7_75t_L g148 ( .A(n_108), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g156 ( .A(n_108), .B(n_140), .Y(n_156) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx1_ASAP7_75t_L g120 ( .A(n_115), .Y(n_120) );
INVx1_ASAP7_75t_L g126 ( .A(n_116), .Y(n_126) );
AND2x4_ASAP7_75t_L g119 ( .A(n_117), .B(n_120), .Y(n_119) );
NAND2x1p5_ASAP7_75t_L g125 ( .A(n_117), .B(n_126), .Y(n_125) );
BUFx12f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_127), .B2(n_128), .Y(n_121) );
INVx3_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_153), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_145), .Y(n_134) );
BUFx4f_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x4_ASAP7_75t_L g142 ( .A(n_140), .B(n_143), .Y(n_142) );
BUFx2_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OR2x6_ASAP7_75t_L g165 ( .A(n_144), .B(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx11_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx6_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_159), .Y(n_153) );
BUFx2_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx8_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx6_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_167), .A2(n_300), .B(n_301), .C(n_302), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g178 ( .A(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
AND3x1_ASAP7_75t_SL g180 ( .A(n_181), .B(n_186), .C(n_189), .Y(n_180) );
INVxp67_ASAP7_75t_L g505 ( .A(n_181), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
INVx1_ASAP7_75t_SL g506 ( .A(n_186), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_186), .A2(n_216), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g515 ( .A(n_186), .Y(n_515) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_187), .B(n_190), .Y(n_509) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_SL g514 ( .A(n_189), .B(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_422), .Y(n_193) );
NOR4xp25_ASAP7_75t_L g194 ( .A(n_195), .B(n_364), .C(n_394), .D(n_404), .Y(n_194) );
OAI211xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_270), .B(n_327), .C(n_354), .Y(n_195) );
OAI222xp33_ASAP7_75t_L g449 ( .A1(n_196), .A2(n_369), .B1(n_450), .B2(n_451), .C1(n_452), .C2(n_453), .Y(n_449) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_245), .Y(n_196) );
AOI33xp33_ASAP7_75t_L g375 ( .A1(n_197), .A2(n_362), .A3(n_363), .B1(n_376), .B2(n_381), .B3(n_383), .Y(n_375) );
OAI211xp5_ASAP7_75t_SL g432 ( .A1(n_197), .A2(n_433), .B(n_435), .C(n_437), .Y(n_432) );
OR2x2_ASAP7_75t_L g448 ( .A(n_197), .B(n_434), .Y(n_448) );
INVx1_ASAP7_75t_L g481 ( .A(n_197), .Y(n_481) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_232), .Y(n_197) );
INVx2_ASAP7_75t_L g358 ( .A(n_198), .Y(n_358) );
AND2x2_ASAP7_75t_L g374 ( .A(n_198), .B(n_261), .Y(n_374) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_198), .Y(n_409) );
AND2x2_ASAP7_75t_L g438 ( .A(n_198), .B(n_232), .Y(n_438) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_206), .B(n_229), .Y(n_198) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_199), .A2(n_262), .B(n_269), .Y(n_261) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_199), .A2(n_275), .B(n_283), .Y(n_274) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx4_ASAP7_75t_L g231 ( .A(n_200), .Y(n_231) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g315 ( .A(n_201), .Y(n_315) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
AND2x2_ASAP7_75t_SL g233 ( .A(n_202), .B(n_203), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
BUFx2_ASAP7_75t_L g317 ( .A(n_207), .Y(n_317) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_212), .Y(n_207) );
NAND2x1p5_ASAP7_75t_L g251 ( .A(n_208), .B(n_212), .Y(n_251) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_211), .Y(n_208) );
INVx1_ASAP7_75t_L g303 ( .A(n_209), .Y(n_303) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g217 ( .A(n_210), .Y(n_217) );
INVx1_ASAP7_75t_L g227 ( .A(n_210), .Y(n_227) );
INVx1_ASAP7_75t_L g218 ( .A(n_211), .Y(n_218) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_211), .Y(n_221) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_211), .Y(n_225) );
INVx3_ASAP7_75t_L g241 ( .A(n_211), .Y(n_241) );
INVx4_ASAP7_75t_SL g228 ( .A(n_212), .Y(n_228) );
BUFx3_ASAP7_75t_L g304 ( .A(n_212), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_SL g213 ( .A1(n_214), .A2(n_215), .B(n_219), .C(n_228), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_SL g235 ( .A1(n_215), .A2(n_228), .B(n_236), .C(n_237), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_SL g263 ( .A1(n_215), .A2(n_228), .B(n_264), .C(n_265), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g276 ( .A1(n_215), .A2(n_228), .B(n_277), .C(n_278), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_SL g318 ( .A1(n_215), .A2(n_228), .B(n_319), .C(n_320), .Y(n_318) );
INVx5_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g498 ( .A(n_216), .B(n_304), .Y(n_498) );
AND2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
BUFx3_ASAP7_75t_L g243 ( .A(n_217), .Y(n_243) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_217), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_220), .B(n_280), .Y(n_279) );
INVx4_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g238 ( .A(n_221), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_224), .B(n_267), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g321 ( .A1(n_224), .A2(n_300), .B1(n_322), .B2(n_323), .Y(n_321) );
INVx4_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g256 ( .A(n_225), .Y(n_256) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g291 ( .A(n_228), .Y(n_291) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_231), .B(n_260), .Y(n_259) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_231), .A2(n_285), .B(n_292), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_231), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g338 ( .A(n_232), .Y(n_338) );
BUFx3_ASAP7_75t_L g346 ( .A(n_232), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_232), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g357 ( .A(n_232), .B(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_232), .B(n_246), .Y(n_386) );
AND2x2_ASAP7_75t_L g455 ( .A(n_232), .B(n_389), .Y(n_455) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_244), .Y(n_232) );
INVx1_ASAP7_75t_L g248 ( .A(n_233), .Y(n_248) );
INVx2_ASAP7_75t_L g294 ( .A(n_233), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g296 ( .A1(n_233), .A2(n_251), .B(n_297), .C(n_298), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx5_ASAP7_75t_L g300 ( .A(n_241), .Y(n_300) );
INVx2_ASAP7_75t_L g258 ( .A(n_242), .Y(n_258) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g268 ( .A(n_243), .Y(n_268) );
INVx2_ASAP7_75t_SL g349 ( .A(n_245), .Y(n_349) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_261), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_246), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g391 ( .A(n_246), .Y(n_391) );
AND2x2_ASAP7_75t_L g402 ( .A(n_246), .B(n_358), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_246), .B(n_387), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_246), .B(n_389), .Y(n_434) );
AND2x2_ASAP7_75t_L g493 ( .A(n_246), .B(n_438), .Y(n_493) );
INVx4_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g363 ( .A(n_247), .B(n_261), .Y(n_363) );
AND2x2_ASAP7_75t_L g373 ( .A(n_247), .B(n_374), .Y(n_373) );
BUFx3_ASAP7_75t_L g395 ( .A(n_247), .Y(n_395) );
AND3x2_ASAP7_75t_L g454 ( .A(n_247), .B(n_455), .C(n_456), .Y(n_454) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_259), .Y(n_247) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_252), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g285 ( .A1(n_251), .A2(n_286), .B(n_287), .Y(n_285) );
O2A1O1Ixp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_257), .C(n_258), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g288 ( .A1(n_255), .A2(n_258), .B(n_289), .C(n_290), .Y(n_288) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_261), .Y(n_345) );
INVx1_ASAP7_75t_SL g389 ( .A(n_261), .Y(n_389) );
NAND3xp33_ASAP7_75t_L g401 ( .A(n_261), .B(n_338), .C(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_307), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g424 ( .A1(n_271), .A2(n_373), .B(n_425), .C(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_273), .B(n_295), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_273), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_SL g441 ( .A(n_273), .Y(n_441) );
AND2x2_ASAP7_75t_L g462 ( .A(n_273), .B(n_309), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_273), .B(n_371), .Y(n_490) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_284), .Y(n_273) );
AND2x2_ASAP7_75t_L g335 ( .A(n_274), .B(n_326), .Y(n_335) );
INVx2_ASAP7_75t_L g342 ( .A(n_274), .Y(n_342) );
AND2x2_ASAP7_75t_L g362 ( .A(n_274), .B(n_309), .Y(n_362) );
AND2x2_ASAP7_75t_L g412 ( .A(n_274), .B(n_295), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_274), .Y(n_416) );
OAI322xp33_ASAP7_75t_L g499 ( .A1(n_277), .A2(n_500), .A3(n_502), .B1(n_506), .B2(n_507), .C1(n_510), .C2(n_512), .Y(n_499) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_SL g326 ( .A(n_284), .Y(n_326) );
BUFx2_ASAP7_75t_L g352 ( .A(n_284), .Y(n_352) );
AND2x2_ASAP7_75t_L g479 ( .A(n_284), .B(n_295), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g325 ( .A(n_294), .Y(n_325) );
INVx3_ASAP7_75t_SL g309 ( .A(n_295), .Y(n_309) );
AND2x2_ASAP7_75t_L g334 ( .A(n_295), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g341 ( .A(n_295), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g371 ( .A(n_295), .B(n_331), .Y(n_371) );
OR2x2_ASAP7_75t_L g380 ( .A(n_295), .B(n_326), .Y(n_380) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_295), .Y(n_398) );
AND2x2_ASAP7_75t_L g403 ( .A(n_295), .B(n_356), .Y(n_403) );
AND2x2_ASAP7_75t_L g431 ( .A(n_295), .B(n_311), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_295), .B(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g469 ( .A(n_295), .B(n_310), .Y(n_469) );
OR2x6_ASAP7_75t_L g295 ( .A(n_296), .B(n_305), .Y(n_295) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_303), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x2_ASAP7_75t_L g393 ( .A(n_309), .B(n_342), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_309), .B(n_335), .Y(n_421) );
AND2x2_ASAP7_75t_L g439 ( .A(n_309), .B(n_356), .Y(n_439) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_326), .Y(n_310) );
AND2x2_ASAP7_75t_L g340 ( .A(n_311), .B(n_326), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_311), .B(n_369), .Y(n_368) );
BUFx3_ASAP7_75t_L g378 ( .A(n_311), .Y(n_378) );
OR2x2_ASAP7_75t_L g426 ( .A(n_311), .B(n_346), .Y(n_426) );
OA21x2_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_316), .B(n_324), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AO21x2_ASAP7_75t_L g331 ( .A1(n_313), .A2(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g332 ( .A(n_316), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_324), .Y(n_333) );
AND2x2_ASAP7_75t_L g361 ( .A(n_326), .B(n_331), .Y(n_361) );
INVx1_ASAP7_75t_L g369 ( .A(n_326), .Y(n_369) );
AND2x2_ASAP7_75t_L g464 ( .A(n_326), .B(n_342), .Y(n_464) );
AOI222xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_336), .B1(n_339), .B2(n_343), .C1(n_347), .C2(n_350), .Y(n_327) );
INVx1_ASAP7_75t_L g459 ( .A(n_328), .Y(n_459) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_334), .Y(n_328) );
AND2x2_ASAP7_75t_L g355 ( .A(n_329), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g366 ( .A(n_329), .B(n_335), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_329), .B(n_357), .Y(n_382) );
OAI222xp33_ASAP7_75t_L g404 ( .A1(n_329), .A2(n_405), .B1(n_410), .B2(n_411), .C1(n_419), .C2(n_421), .Y(n_404) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g392 ( .A(n_331), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_331), .B(n_412), .Y(n_452) );
AND2x2_ASAP7_75t_L g463 ( .A(n_331), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g471 ( .A(n_334), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_336), .B(n_387), .Y(n_450) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_338), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g408 ( .A(n_338), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx3_ASAP7_75t_L g353 ( .A(n_341), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g443 ( .A1(n_341), .A2(n_444), .B(n_447), .C(n_449), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_341), .B(n_378), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_341), .B(n_361), .Y(n_483) );
AND2x2_ASAP7_75t_L g356 ( .A(n_342), .B(n_352), .Y(n_356) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g383 ( .A(n_345), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_346), .B(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g435 ( .A(n_346), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g474 ( .A(n_346), .B(n_374), .Y(n_474) );
INVx1_ASAP7_75t_L g486 ( .A(n_346), .Y(n_486) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_349), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g467 ( .A(n_352), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_357), .B(n_359), .C(n_363), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_355), .A2(n_385), .B1(n_400), .B2(n_403), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_356), .B(n_370), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_356), .B(n_378), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_357), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g420 ( .A(n_357), .Y(n_420) );
AND2x2_ASAP7_75t_L g427 ( .A(n_357), .B(n_407), .Y(n_427) );
INVx2_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
NOR4xp25_ASAP7_75t_L g365 ( .A(n_362), .B(n_366), .C(n_367), .D(n_370), .Y(n_365) );
INVx1_ASAP7_75t_SL g436 ( .A(n_363), .Y(n_436) );
AND2x2_ASAP7_75t_L g480 ( .A(n_363), .B(n_481), .Y(n_480) );
OAI211xp5_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_372), .B(n_375), .C(n_384), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_371), .B(n_441), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_373), .A2(n_492), .B1(n_493), .B2(n_494), .Y(n_491) );
INVx1_ASAP7_75t_SL g446 ( .A(n_374), .Y(n_446) );
AND2x2_ASAP7_75t_L g485 ( .A(n_374), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_378), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_382), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_383), .B(n_408), .Y(n_468) );
OAI21xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_390), .B(n_392), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g460 ( .A(n_387), .Y(n_460) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx2_ASAP7_75t_L g488 ( .A(n_388), .Y(n_488) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_389), .Y(n_415) );
OAI21xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B(n_399), .Y(n_394) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_395), .Y(n_407) );
OR2x2_ASAP7_75t_L g445 ( .A(n_395), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI21xp33_ASAP7_75t_SL g440 ( .A1(n_398), .A2(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_402), .A2(n_429), .B1(n_432), .B2(n_439), .C(n_440), .Y(n_428) );
INVx1_ASAP7_75t_SL g472 ( .A(n_403), .Y(n_472) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
OR2x2_ASAP7_75t_L g419 ( .A(n_407), .B(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g456 ( .A(n_409), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_416), .B2(n_417), .Y(n_411) );
INVx1_ASAP7_75t_L g451 ( .A(n_412), .Y(n_451) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_415), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NOR4xp25_ASAP7_75t_L g422 ( .A(n_423), .B(n_457), .C(n_470), .D(n_482), .Y(n_422) );
NAND3xp33_ASAP7_75t_SL g423 ( .A(n_424), .B(n_428), .C(n_443), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_426), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_433), .B(n_438), .Y(n_442) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI221xp5_ASAP7_75t_SL g470 ( .A1(n_445), .A2(n_471), .B1(n_472), .B2(n_473), .C(n_475), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_447), .A2(n_462), .B(n_463), .C(n_465), .Y(n_461) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_448), .A2(n_466), .B1(n_468), .B2(n_469), .Y(n_465) );
INVx2_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_460), .C(n_461), .Y(n_457) );
INVx1_ASAP7_75t_L g476 ( .A(n_469), .Y(n_476) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OAI21xp5_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_477), .B(n_480), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI221xp5_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_484), .B1(n_487), .B2(n_489), .C(n_491), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVxp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
CKINVDCx14_ASAP7_75t_R g502 ( .A(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
endmodule