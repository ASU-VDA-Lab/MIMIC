module fake_jpeg_22976_n_75 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_75);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_38;
wire n_74;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_69;
wire n_40;
wire n_71;
wire n_48;
wire n_35;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_70;
wire n_66;

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_2),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_42),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_45),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_48),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_40),
.B1(n_35),
.B2(n_37),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_1),
.B1(n_3),
.B2(n_38),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_36),
.B1(n_1),
.B2(n_3),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_39),
.B1(n_34),
.B2(n_6),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_4),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

OAI22x1_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_49),
.B1(n_5),
.B2(n_9),
.Y(n_58)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_19),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_16),
.C(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_64),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_66),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_60),
.B(n_67),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_64),
.B(n_21),
.Y(n_71)
);

OAI31xp33_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_20),
.A3(n_22),
.B(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_25),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_27),
.C(n_28),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_29),
.Y(n_75)
);


endmodule