module fake_jpeg_18638_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_22),
.B1(n_32),
.B2(n_27),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_46),
.B1(n_56),
.B2(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_22),
.B1(n_32),
.B2(n_27),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_47),
.B1(n_35),
.B2(n_41),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_22),
.B1(n_27),
.B2(n_31),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_30),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_16),
.B1(n_29),
.B2(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_57),
.B(n_60),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_35),
.B1(n_55),
.B2(n_30),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_59),
.B(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_45),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_33),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_37),
.C(n_41),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_33),
.B1(n_39),
.B2(n_35),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_67),
.Y(n_88)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_33),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_24),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_25),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_77),
.B1(n_78),
.B2(n_81),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_16),
.B1(n_29),
.B2(n_17),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_21),
.B1(n_34),
.B2(n_37),
.Y(n_107)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_76),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_35),
.B1(n_26),
.B2(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_30),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_83),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_85),
.B1(n_81),
.B2(n_100),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_41),
.B1(n_28),
.B2(n_37),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_72),
.B1(n_71),
.B2(n_60),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_SL g97 ( 
.A(n_83),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_34),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_65),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_34),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_100),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_66),
.A3(n_59),
.B1(n_67),
.B2(n_57),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_20),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

BUFx16f_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_64),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_115),
.B1(n_127),
.B2(n_130),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_99),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_121),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_91),
.B(n_63),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_78),
.C(n_84),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_128),
.C(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_133),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_74),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_126),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_80),
.B(n_73),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_101),
.B(n_86),
.Y(n_153)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_82),
.B1(n_76),
.B2(n_20),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_37),
.C(n_20),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_89),
.A2(n_21),
.B1(n_64),
.B2(n_2),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_15),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_87),
.B1(n_94),
.B2(n_90),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_88),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_142),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_114),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_151),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_105),
.C(n_101),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_146),
.C(n_147),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_105),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_90),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_110),
.C(n_128),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_153),
.A2(n_132),
.B(n_131),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_113),
.A2(n_104),
.B1(n_103),
.B2(n_93),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_155),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_113),
.A2(n_104),
.B1(n_103),
.B2(n_108),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_134),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_169),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_166),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_114),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_125),
.B1(n_130),
.B2(n_123),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_114),
.B(n_123),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_145),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_108),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_12),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g179 ( 
.A(n_172),
.Y(n_179)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_146),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_178),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_147),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_163),
.B(n_151),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_186),
.C(n_169),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_162),
.A2(n_150),
.B1(n_142),
.B2(n_143),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_190),
.B1(n_161),
.B2(n_170),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_150),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_162),
.A2(n_161),
.B1(n_168),
.B2(n_165),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_201),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_186),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_164),
.C(n_152),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_177),
.C(n_178),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_158),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

HB1xp67_ASAP7_75t_SL g195 ( 
.A(n_184),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_195),
.A2(n_200),
.B(n_187),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_185),
.A2(n_174),
.B1(n_154),
.B2(n_155),
.Y(n_197)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_190),
.A2(n_140),
.B1(n_14),
.B2(n_12),
.Y(n_198)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_1),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_189),
.B(n_182),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_189),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_196),
.C(n_192),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_198),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_196),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_215),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_206),
.A2(n_201),
.B(n_199),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_212),
.A2(n_213),
.B(n_193),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_217),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_202),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_179),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_197),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_220),
.B(n_221),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_210),
.C(n_208),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_224),
.A3(n_218),
.B1(n_4),
.B2(n_5),
.C1(n_7),
.C2(n_3),
.Y(n_227)
);

AO21x1_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_2),
.B(n_3),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_225),
.A2(n_218),
.B(n_4),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_226),
.Y(n_228)
);

AOI321xp33_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_227),
.A3(n_5),
.B1(n_7),
.B2(n_8),
.C(n_4),
.Y(n_229)
);

OAI321xp33_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_11),
.Y(n_231)
);


endmodule