module fake_jpeg_30209_n_116 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_116);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_1),
.B(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_54),
.Y(n_63)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_17),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_47),
.C(n_48),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_62),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_38),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_49),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_68),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_39),
.B(n_38),
.C(n_3),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_54),
.B1(n_44),
.B2(n_39),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_87),
.B(n_6),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_61),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_79),
.Y(n_96)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_85),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_88),
.B1(n_6),
.B2(n_7),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_2),
.B(n_5),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_20),
.B1(n_35),
.B2(n_34),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_95),
.B1(n_8),
.B2(n_9),
.Y(n_103)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_97),
.B1(n_18),
.B2(n_19),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_99),
.B(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_80),
.C(n_86),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_23),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_90),
.B(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_8),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_104),
.Y(n_111)
);

AOI221xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_107),
.B1(n_108),
.B2(n_101),
.C(n_27),
.Y(n_110)
);

OAI22x1_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_109),
.B(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_111),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_99),
.C(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_94),
.Y(n_115)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_105),
.A3(n_98),
.B1(n_29),
.B2(n_30),
.C1(n_24),
.C2(n_33),
.Y(n_116)
);


endmodule