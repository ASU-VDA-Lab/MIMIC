module fake_jpeg_31305_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

HB1xp67_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx16f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx12_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_SL g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_SL g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_22),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_23),
.Y(n_26)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_17),
.A2(n_14),
.B1(n_15),
.B2(n_12),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_20),
.B1(n_18),
.B2(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_14),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_34),
.C(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_19),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_35),
.B1(n_22),
.B2(n_23),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_9),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_39),
.C(n_41),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_29),
.B(n_2),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_43),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_26),
.C(n_29),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_13),
.B(n_1),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_50),
.C(n_45),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_49),
.B(n_50),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.C(n_13),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_13),
.C(n_10),
.Y(n_54)
);

NOR3xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_6),
.C(n_1),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_6),
.B1(n_10),
.B2(n_16),
.Y(n_57)
);


endmodule