module fake_ibex_1983_n_913 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_913);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_913;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_732;
wire n_673;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_807;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g166 ( 
.A(n_47),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_25),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_43),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_62),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_93),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_108),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_5),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_71),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_9),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_12),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_48),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_30),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_18),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_5),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_34),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_11),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_9),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_130),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_4),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_58),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_88),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_135),
.B(n_36),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_46),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_111),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_131),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_76),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_95),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_35),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_52),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_114),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_63),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_56),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_96),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_98),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_57),
.B(n_104),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_25),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_69),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_38),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_55),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_30),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_94),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_31),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_20),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_128),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_15),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_89),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_156),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_129),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_155),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_82),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_26),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_160),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_21),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_138),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_64),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_99),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_67),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_110),
.Y(n_243)
);

BUFx4f_ASAP7_75t_SL g244 ( 
.A(n_12),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_18),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_20),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_42),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_92),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_97),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_78),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_L g251 ( 
.A(n_42),
.B(n_31),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_84),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_112),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_75),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_85),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_86),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_117),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_74),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_40),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_147),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_72),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_8),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_120),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_101),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_113),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_87),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_106),
.B(n_150),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_125),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_39),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_35),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_23),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_45),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_24),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_21),
.Y(n_274)
);

INVx4_ASAP7_75t_SL g275 ( 
.A(n_222),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_187),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_223),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_278)
);

INVxp33_ASAP7_75t_SL g279 ( 
.A(n_212),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_221),
.B(n_0),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_199),
.Y(n_283)
);

AND2x4_ASAP7_75t_L g284 ( 
.A(n_187),
.B(n_1),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_210),
.Y(n_286)
);

AOI22x1_ASAP7_75t_SL g287 ( 
.A1(n_223),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_287)
);

BUFx8_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_187),
.B(n_3),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_199),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_207),
.Y(n_292)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_222),
.B(n_44),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_207),
.A2(n_91),
.B(n_164),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_214),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_214),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_258),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_255),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_192),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_188),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_237),
.B(n_6),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_208),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_208),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_192),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_237),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_181),
.B(n_7),
.Y(n_309)
);

AOI22x1_ASAP7_75t_SL g310 ( 
.A1(n_181),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_179),
.B(n_10),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_197),
.B(n_225),
.Y(n_312)
);

BUFx12f_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_190),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_190),
.B(n_11),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_194),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_245),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_227),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_245),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_166),
.B(n_13),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_230),
.B(n_14),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_247),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_323)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_258),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_262),
.B(n_271),
.Y(n_327)
);

AND2x2_ASAP7_75t_SL g328 ( 
.A(n_203),
.B(n_167),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_259),
.B(n_17),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_249),
.B(n_19),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_228),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_244),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_249),
.B(n_22),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_274),
.B(n_170),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_236),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_169),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_172),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_173),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_174),
.B(n_27),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_236),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_246),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_177),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g343 ( 
.A(n_266),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_168),
.B(n_29),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_246),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_169),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_184),
.B(n_32),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_286),
.B(n_180),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

OAI21xp33_ASAP7_75t_SL g350 ( 
.A1(n_328),
.A2(n_251),
.B(n_186),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_280),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

BUFx8_ASAP7_75t_SL g354 ( 
.A(n_313),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_308),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_284),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

BUFx6f_ASAP7_75t_SL g358 ( 
.A(n_328),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_346),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_314),
.B(n_168),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_304),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_289),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_276),
.B(n_168),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_279),
.B(n_261),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_289),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_289),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_304),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_277),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_277),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_276),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_279),
.B(n_261),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_290),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_290),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_276),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_343),
.B(n_263),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_281),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_300),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_281),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_293),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_315),
.A2(n_269),
.B1(n_273),
.B2(n_270),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_330),
.B(n_171),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_315),
.A2(n_189),
.B1(n_183),
.B2(n_220),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_300),
.Y(n_385)
);

NAND3xp33_ASAP7_75t_L g386 ( 
.A(n_322),
.B(n_193),
.C(n_191),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_337),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_299),
.B(n_195),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_337),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_299),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_293),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_311),
.A2(n_233),
.B1(n_231),
.B2(n_235),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_305),
.B(n_175),
.Y(n_394)
);

AO21x2_ASAP7_75t_L g395 ( 
.A1(n_294),
.A2(n_219),
.B(n_201),
.Y(n_395)
);

AND2x6_ASAP7_75t_L g396 ( 
.A(n_329),
.B(n_198),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_297),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_288),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_330),
.B(n_182),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_297),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_333),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_303),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_334),
.B(n_202),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_305),
.B(n_176),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_283),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_306),
.B(n_204),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_333),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_321),
.B(n_209),
.C(n_205),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_R g410 ( 
.A(n_288),
.B(n_206),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_324),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_306),
.B(n_178),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_283),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_319),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_324),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_324),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_291),
.Y(n_418)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_319),
.Y(n_419)
);

INVx6_ASAP7_75t_L g420 ( 
.A(n_275),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_291),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_320),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_320),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_326),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_292),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_326),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_292),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_295),
.Y(n_428)
);

AND3x2_ASAP7_75t_L g429 ( 
.A(n_344),
.B(n_215),
.C(n_213),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_275),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_295),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_296),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_317),
.B(n_185),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_346),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_296),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_298),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_325),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_298),
.Y(n_438)
);

AOI21x1_ASAP7_75t_L g439 ( 
.A1(n_294),
.A2(n_218),
.B(n_217),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_360),
.B(n_344),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_348),
.B(n_288),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_363),
.B(n_311),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_366),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_354),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_363),
.B(n_282),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_361),
.B(n_338),
.Y(n_447)
);

OAI22xp33_ASAP7_75t_L g448 ( 
.A1(n_361),
.A2(n_336),
.B1(n_318),
.B2(n_323),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_368),
.B(n_401),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_SL g450 ( 
.A(n_382),
.B(n_309),
.C(n_231),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_364),
.B(n_312),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_358),
.A2(n_252),
.B1(n_264),
.B2(n_235),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_353),
.B(n_339),
.Y(n_454)
);

O2A1O1Ixp5_ASAP7_75t_L g455 ( 
.A1(n_439),
.A2(n_347),
.B(n_342),
.C(n_301),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_395),
.A2(n_367),
.B(n_366),
.Y(n_456)
);

O2A1O1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_350),
.A2(n_327),
.B(n_331),
.C(n_345),
.Y(n_457)
);

NAND3xp33_ASAP7_75t_L g458 ( 
.A(n_384),
.B(n_310),
.C(n_287),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_401),
.B(n_341),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_376),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_353),
.B(n_196),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_408),
.B(n_388),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_373),
.B(n_340),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_360),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_358),
.A2(n_233),
.B1(n_252),
.B2(n_232),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_372),
.B(n_200),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_429),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_383),
.B(n_341),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_396),
.A2(n_352),
.B1(n_357),
.B2(n_356),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_381),
.B(n_211),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_381),
.B(n_216),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_358),
.A2(n_232),
.B1(n_206),
.B2(n_264),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_395),
.A2(n_229),
.B(n_224),
.Y(n_473)
);

A2O1A1Ixp33_ASAP7_75t_L g474 ( 
.A1(n_403),
.A2(n_397),
.B(n_400),
.C(n_350),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_R g475 ( 
.A(n_355),
.B(n_272),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_399),
.B(n_302),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_388),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_396),
.A2(n_272),
.B1(n_278),
.B2(n_332),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_396),
.A2(n_310),
.B1(n_287),
.B2(n_257),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_388),
.B(n_335),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_388),
.B(n_335),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_376),
.B(n_307),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_393),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_390),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_390),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_351),
.B(n_316),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_391),
.B(n_226),
.Y(n_488)
);

OR2x6_ASAP7_75t_L g489 ( 
.A(n_398),
.B(n_316),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_395),
.A2(n_256),
.B(n_239),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_396),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_397),
.Y(n_492)
);

AOI221xp5_ASAP7_75t_L g493 ( 
.A1(n_386),
.A2(n_260),
.B1(n_268),
.B2(n_250),
.C(n_248),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_402),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_391),
.B(n_234),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_414),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_396),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_437),
.B(n_241),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_377),
.B(n_267),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_414),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_352),
.B(n_275),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_356),
.B(n_275),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_357),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_410),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_359),
.B(n_37),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_362),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_362),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_392),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_464),
.B(n_355),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_456),
.A2(n_392),
.B(n_433),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_451),
.B(n_409),
.Y(n_511)
);

AOI21x1_ASAP7_75t_L g512 ( 
.A1(n_456),
.A2(n_439),
.B(n_370),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_443),
.B(n_409),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_473),
.A2(n_404),
.B(n_394),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_475),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_473),
.A2(n_412),
.B(n_407),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_487),
.Y(n_517)
);

OAI21xp33_ASAP7_75t_L g518 ( 
.A1(n_446),
.A2(n_370),
.B(n_369),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_440),
.B(n_463),
.Y(n_519)
);

AOI221xp5_ASAP7_75t_L g520 ( 
.A1(n_483),
.A2(n_428),
.B1(n_436),
.B2(n_418),
.C(n_406),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_504),
.B(n_434),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_489),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_489),
.B(n_427),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_453),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_469),
.B(n_365),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_489),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_508),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_508),
.Y(n_528)
);

NOR2x1_ASAP7_75t_L g529 ( 
.A(n_450),
.B(n_378),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_459),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_444),
.B(n_413),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_444),
.B(n_413),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_483),
.A2(n_380),
.B1(n_436),
.B2(n_428),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_447),
.B(n_418),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_465),
.Y(n_535)
);

NOR2x1_ASAP7_75t_L g536 ( 
.A(n_450),
.B(n_421),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_455),
.A2(n_422),
.B(n_423),
.Y(n_537)
);

A2O1A1Ixp33_ASAP7_75t_L g538 ( 
.A1(n_457),
.A2(n_426),
.B(n_424),
.C(n_432),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_448),
.A2(n_421),
.B1(n_425),
.B2(n_432),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_449),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_492),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_477),
.A2(n_425),
.B1(n_435),
.B2(n_431),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_454),
.A2(n_430),
.B(n_426),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_490),
.A2(n_424),
.B(n_430),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_462),
.A2(n_438),
.B1(n_419),
.B2(n_405),
.Y(n_545)
);

AO22x1_ASAP7_75t_L g546 ( 
.A1(n_445),
.A2(n_419),
.B1(n_41),
.B2(n_417),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_467),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_493),
.A2(n_419),
.B1(n_415),
.B2(n_417),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_472),
.B(n_419),
.Y(n_549)
);

AOI21x1_ASAP7_75t_L g550 ( 
.A1(n_501),
.A2(n_416),
.B(n_415),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_494),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_502),
.A2(n_387),
.B(n_389),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_455),
.A2(n_387),
.B(n_389),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_507),
.Y(n_554)
);

A2O1A1Ixp33_ASAP7_75t_L g555 ( 
.A1(n_457),
.A2(n_405),
.B(n_411),
.C(n_374),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_468),
.B(n_420),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_478),
.B(n_411),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_494),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_476),
.B(n_420),
.Y(n_559)
);

O2A1O1Ixp33_ASAP7_75t_L g560 ( 
.A1(n_448),
.A2(n_385),
.B(n_379),
.C(n_375),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_480),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_481),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_498),
.B(n_49),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_491),
.B(n_482),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_497),
.A2(n_506),
.B1(n_503),
.B2(n_486),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_497),
.A2(n_506),
.B1(n_503),
.B2(n_479),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_499),
.B(n_50),
.Y(n_567)
);

INVx4_ASAP7_75t_SL g568 ( 
.A(n_442),
.Y(n_568)
);

O2A1O1Ixp33_ASAP7_75t_SL g569 ( 
.A1(n_461),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_499),
.B(n_59),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_496),
.A2(n_349),
.B(n_61),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_458),
.A2(n_349),
.B1(n_65),
.B2(n_66),
.Y(n_572)
);

O2A1O1Ixp33_ASAP7_75t_SL g573 ( 
.A1(n_466),
.A2(n_60),
.B(n_68),
.C(n_70),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_452),
.A2(n_77),
.B(n_79),
.Y(n_574)
);

AO21x1_ASAP7_75t_L g575 ( 
.A1(n_460),
.A2(n_80),
.B(n_81),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_505),
.B(n_83),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_484),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_485),
.Y(n_578)
);

O2A1O1Ixp33_ASAP7_75t_SL g579 ( 
.A1(n_470),
.A2(n_495),
.B(n_471),
.C(n_488),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_500),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_517),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_531),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_535),
.B(n_103),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_517),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_544),
.A2(n_107),
.B(n_109),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_540),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_530),
.Y(n_587)
);

BUFx4f_ASAP7_75t_L g588 ( 
.A(n_515),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_532),
.A2(n_539),
.B1(n_534),
.B2(n_520),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_541),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_526),
.Y(n_591)
);

A2O1A1Ixp33_ASAP7_75t_L g592 ( 
.A1(n_511),
.A2(n_115),
.B(n_116),
.C(n_118),
.Y(n_592)
);

O2A1O1Ixp33_ASAP7_75t_SL g593 ( 
.A1(n_563),
.A2(n_121),
.B(n_124),
.C(n_127),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_520),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g595 ( 
.A1(n_514),
.A2(n_137),
.B(n_140),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_524),
.B(n_141),
.Y(n_596)
);

A2O1A1Ixp33_ASAP7_75t_L g597 ( 
.A1(n_516),
.A2(n_143),
.B(n_144),
.C(n_146),
.Y(n_597)
);

OAI22x1_ASAP7_75t_L g598 ( 
.A1(n_536),
.A2(n_148),
.B1(n_149),
.B2(n_151),
.Y(n_598)
);

OAI22x1_ASAP7_75t_L g599 ( 
.A1(n_529),
.A2(n_152),
.B1(n_153),
.B2(n_157),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_523),
.Y(n_600)
);

INVxp67_ASAP7_75t_SL g601 ( 
.A(n_517),
.Y(n_601)
);

O2A1O1Ixp33_ASAP7_75t_L g602 ( 
.A1(n_513),
.A2(n_533),
.B(n_565),
.C(n_564),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_554),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_557),
.B(n_561),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_562),
.B(n_523),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_577),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_578),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_567),
.A2(n_570),
.B(n_576),
.Y(n_608)
);

AO31x2_ASAP7_75t_L g609 ( 
.A1(n_555),
.A2(n_516),
.A3(n_538),
.B(n_571),
.Y(n_609)
);

AOI211x1_ASAP7_75t_L g610 ( 
.A1(n_518),
.A2(n_546),
.B(n_542),
.C(n_572),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_580),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_549),
.B(n_509),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_547),
.B(n_568),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_527),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_521),
.B(n_528),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_551),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_568),
.B(n_558),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_548),
.B(n_545),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_525),
.A2(n_552),
.B(n_543),
.Y(n_619)
);

AOI221x1_ASAP7_75t_L g620 ( 
.A1(n_556),
.A2(n_559),
.B1(n_569),
.B2(n_573),
.C(n_579),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_522),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_524),
.B(n_483),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_522),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_519),
.B(n_451),
.Y(n_624)
);

AOI21xp33_ASAP7_75t_L g625 ( 
.A1(n_509),
.A2(n_441),
.B(n_483),
.Y(n_625)
);

AOI221xp5_ASAP7_75t_L g626 ( 
.A1(n_519),
.A2(n_448),
.B1(n_483),
.B2(n_451),
.C(n_350),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_540),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_519),
.B(n_451),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_512),
.A2(n_553),
.B(n_550),
.Y(n_629)
);

AND2x2_ASAP7_75t_SL g630 ( 
.A(n_515),
.B(n_453),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_517),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_515),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_515),
.B(n_393),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_519),
.B(n_451),
.Y(n_634)
);

OA21x2_ASAP7_75t_L g635 ( 
.A1(n_537),
.A2(n_490),
.B(n_473),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_519),
.B(n_451),
.Y(n_636)
);

AO31x2_ASAP7_75t_L g637 ( 
.A1(n_575),
.A2(n_490),
.A3(n_473),
.B(n_456),
.Y(n_637)
);

NAND2x1p5_ASAP7_75t_L g638 ( 
.A(n_522),
.B(n_526),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_540),
.Y(n_639)
);

O2A1O1Ixp5_ASAP7_75t_L g640 ( 
.A1(n_514),
.A2(n_510),
.B(n_516),
.C(n_490),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_531),
.A2(n_532),
.B1(n_539),
.B2(n_566),
.Y(n_641)
);

OAI21x1_ASAP7_75t_SL g642 ( 
.A1(n_566),
.A2(n_487),
.B(n_574),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_512),
.A2(n_553),
.B(n_550),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_515),
.Y(n_644)
);

INVxp33_ASAP7_75t_SL g645 ( 
.A(n_521),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_519),
.B(n_451),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_540),
.Y(n_647)
);

NAND2x1p5_ASAP7_75t_L g648 ( 
.A(n_522),
.B(n_526),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_540),
.Y(n_649)
);

AO21x2_ASAP7_75t_L g650 ( 
.A1(n_544),
.A2(n_490),
.B(n_473),
.Y(n_650)
);

NOR4xp25_ASAP7_75t_L g651 ( 
.A(n_560),
.B(n_457),
.C(n_350),
.D(n_474),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_519),
.B(n_451),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_540),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_540),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_512),
.A2(n_553),
.B(n_550),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_515),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_522),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_SL g658 ( 
.A1(n_582),
.A2(n_641),
.B(n_589),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_586),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_640),
.A2(n_602),
.B(n_641),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_627),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_581),
.Y(n_662)
);

OA21x2_ASAP7_75t_L g663 ( 
.A1(n_629),
.A2(n_643),
.B(n_655),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_639),
.Y(n_664)
);

NAND2x1p5_ASAP7_75t_L g665 ( 
.A(n_600),
.B(n_613),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_647),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_624),
.B(n_628),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_649),
.B(n_653),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_654),
.B(n_587),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_603),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_634),
.B(n_636),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_588),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_591),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_606),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_646),
.B(n_652),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_590),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_584),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_607),
.Y(n_678)
);

AO31x2_ASAP7_75t_L g679 ( 
.A1(n_620),
.A2(n_598),
.A3(n_599),
.B(n_594),
.Y(n_679)
);

NAND2x1p5_ASAP7_75t_L g680 ( 
.A(n_584),
.B(n_588),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_611),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_635),
.A2(n_650),
.B(n_619),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_632),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_644),
.Y(n_684)
);

NOR2x1_ASAP7_75t_R g685 ( 
.A(n_656),
.B(n_645),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_614),
.Y(n_686)
);

INVxp67_ASAP7_75t_SL g687 ( 
.A(n_604),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_638),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_626),
.B(n_622),
.Y(n_689)
);

AO31x2_ASAP7_75t_L g690 ( 
.A1(n_594),
.A2(n_597),
.A3(n_592),
.B(n_585),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_621),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_616),
.Y(n_692)
);

NAND2x1p5_ASAP7_75t_L g693 ( 
.A(n_631),
.B(n_617),
.Y(n_693)
);

INVx6_ASAP7_75t_L g694 ( 
.A(n_633),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_623),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_648),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_633),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_630),
.B(n_657),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_583),
.Y(n_699)
);

NOR2x1_ASAP7_75t_R g700 ( 
.A(n_612),
.B(n_601),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_625),
.A2(n_618),
.B(n_651),
.C(n_608),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_615),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_650),
.A2(n_651),
.B(n_593),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_608),
.B(n_596),
.Y(n_704)
);

BUFx12f_ASAP7_75t_L g705 ( 
.A(n_610),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_609),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_609),
.B(n_637),
.Y(n_707)
);

AO21x2_ASAP7_75t_L g708 ( 
.A1(n_610),
.A2(n_637),
.B(n_609),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_637),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_586),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_586),
.B(n_627),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_605),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_626),
.B(n_604),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_587),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_586),
.B(n_627),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_582),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_L g717 ( 
.A1(n_640),
.A2(n_602),
.B(n_456),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_624),
.B(n_628),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_586),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_586),
.B(n_627),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_587),
.Y(n_721)
);

NAND2x1p5_ASAP7_75t_L g722 ( 
.A(n_600),
.B(n_522),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_624),
.B(n_628),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_640),
.A2(n_602),
.B(n_456),
.Y(n_724)
);

OAI21x1_ASAP7_75t_SL g725 ( 
.A1(n_594),
.A2(n_595),
.B(n_642),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_667),
.B(n_718),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_716),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_716),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_680),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_663),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_691),
.Y(n_731)
);

BUFx10_ASAP7_75t_L g732 ( 
.A(n_675),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_670),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_680),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_SL g735 ( 
.A1(n_697),
.A2(n_698),
.B1(n_688),
.B2(n_684),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_677),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_674),
.Y(n_737)
);

AO21x2_ASAP7_75t_L g738 ( 
.A1(n_703),
.A2(n_660),
.B(n_724),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_723),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_678),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_675),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_687),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_659),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_661),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_672),
.Y(n_745)
);

OA21x2_ASAP7_75t_L g746 ( 
.A1(n_717),
.A2(n_724),
.B(n_682),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_671),
.B(n_676),
.Y(n_747)
);

BUFx2_ASAP7_75t_R g748 ( 
.A(n_696),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_664),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_666),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_700),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_709),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_710),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_719),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_707),
.Y(n_755)
);

CKINVDCx16_ASAP7_75t_R g756 ( 
.A(n_697),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_691),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_662),
.Y(n_758)
);

BUFx12f_ASAP7_75t_L g759 ( 
.A(n_683),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_714),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_668),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_712),
.B(n_704),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_689),
.B(n_713),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_721),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_701),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_689),
.B(n_713),
.Y(n_766)
);

NAND2x1_ASAP7_75t_L g767 ( 
.A(n_658),
.B(n_725),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_701),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_686),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_712),
.B(n_720),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_704),
.A2(n_702),
.B(n_699),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_681),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_668),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_706),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_665),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_669),
.B(n_720),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_730),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_742),
.Y(n_778)
);

BUFx2_ASAP7_75t_SL g779 ( 
.A(n_732),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_755),
.B(n_708),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_751),
.B(n_696),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_755),
.B(n_708),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_765),
.B(n_705),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_765),
.B(n_669),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_768),
.B(n_715),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_768),
.B(n_715),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_763),
.B(n_679),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_766),
.B(n_679),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_747),
.B(n_711),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_727),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_731),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_747),
.B(n_711),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_728),
.B(n_692),
.Y(n_793)
);

NAND2x1p5_ASAP7_75t_L g794 ( 
.A(n_736),
.B(n_775),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_728),
.B(n_733),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_771),
.B(n_679),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_733),
.B(n_679),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_757),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_737),
.B(n_694),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_762),
.B(n_695),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_770),
.B(n_695),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_740),
.B(n_694),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_767),
.A2(n_693),
.B(n_690),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_758),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_743),
.B(n_673),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_SL g806 ( 
.A(n_751),
.B(n_685),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_743),
.B(n_673),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_752),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_726),
.A2(n_722),
.B1(n_665),
.B2(n_693),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_758),
.B(n_722),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_744),
.B(n_690),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_774),
.B(n_752),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_797),
.B(n_746),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_777),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_805),
.B(n_750),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_800),
.B(n_746),
.Y(n_816)
);

AND2x4_ASAP7_75t_SL g817 ( 
.A(n_789),
.B(n_732),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_778),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_805),
.B(n_750),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_807),
.B(n_753),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_807),
.B(n_753),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_795),
.B(n_754),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_795),
.B(n_754),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_797),
.B(n_746),
.Y(n_824)
);

NAND2x1_ASAP7_75t_SL g825 ( 
.A(n_808),
.B(n_736),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_806),
.B(n_739),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_800),
.B(n_746),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_793),
.B(n_749),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_793),
.B(n_749),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_780),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_811),
.B(n_782),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_811),
.B(n_738),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_782),
.B(n_738),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_818),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_818),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_815),
.B(n_790),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_814),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_819),
.B(n_791),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_820),
.B(n_798),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_821),
.B(n_784),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_816),
.B(n_780),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_826),
.B(n_783),
.Y(n_842)
);

AO22x1_ASAP7_75t_L g843 ( 
.A1(n_828),
.A2(n_804),
.B1(n_812),
.B2(n_808),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_829),
.B(n_822),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_816),
.B(n_787),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_825),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_823),
.B(n_784),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_830),
.B(n_785),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_830),
.B(n_785),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_827),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_845),
.B(n_827),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_850),
.B(n_831),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_842),
.A2(n_783),
.B1(n_789),
.B2(n_792),
.Y(n_853)
);

XNOR2x1_ASAP7_75t_L g854 ( 
.A(n_843),
.B(n_741),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_842),
.A2(n_741),
.B1(n_806),
.B2(n_832),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_836),
.B(n_831),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_837),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_838),
.Y(n_858)
);

NAND4xp25_ASAP7_75t_L g859 ( 
.A(n_839),
.B(n_735),
.C(n_809),
.D(n_787),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_845),
.A2(n_792),
.B1(n_786),
.B2(n_802),
.Y(n_860)
);

NAND3xp33_ASAP7_75t_L g861 ( 
.A(n_843),
.B(n_788),
.C(n_796),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_848),
.A2(n_832),
.B1(n_786),
.B2(n_824),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_834),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_841),
.B(n_813),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_851),
.B(n_841),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_854),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_861),
.A2(n_846),
.B(n_825),
.Y(n_867)
);

NOR2x1_ASAP7_75t_R g868 ( 
.A(n_855),
.B(n_759),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_SL g869 ( 
.A1(n_858),
.A2(n_756),
.B1(n_864),
.B2(n_862),
.Y(n_869)
);

NAND3xp33_ASAP7_75t_L g870 ( 
.A(n_859),
.B(n_788),
.C(n_796),
.Y(n_870)
);

AOI222xp33_ASAP7_75t_L g871 ( 
.A1(n_853),
.A2(n_844),
.B1(n_847),
.B2(n_840),
.C1(n_849),
.C2(n_781),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_864),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_852),
.B(n_813),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_856),
.B(n_857),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_853),
.A2(n_817),
.B(n_767),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_863),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_876),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_865),
.Y(n_878)
);

OAI22xp33_ASAP7_75t_L g879 ( 
.A1(n_870),
.A2(n_810),
.B1(n_804),
.B2(n_801),
.Y(n_879)
);

AOI31xp33_ASAP7_75t_L g880 ( 
.A1(n_868),
.A2(n_860),
.A3(n_794),
.B(n_810),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_872),
.B(n_833),
.Y(n_881)
);

OAI22xp33_ASAP7_75t_SL g882 ( 
.A1(n_866),
.A2(n_867),
.B1(n_875),
.B2(n_869),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_880),
.A2(n_873),
.B1(n_874),
.B2(n_860),
.Y(n_883)
);

NAND4xp25_ASAP7_75t_L g884 ( 
.A(n_882),
.B(n_871),
.C(n_803),
.D(n_868),
.Y(n_884)
);

AOI21xp33_ASAP7_75t_L g885 ( 
.A1(n_879),
.A2(n_745),
.B(n_801),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_884),
.B(n_878),
.Y(n_886)
);

NAND4xp25_ASAP7_75t_SL g887 ( 
.A(n_885),
.B(n_883),
.C(n_877),
.D(n_881),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_L g888 ( 
.A(n_886),
.B(n_877),
.C(n_879),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_887),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_889),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_888),
.B(n_745),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_890),
.B(n_835),
.Y(n_892)
);

NAND3xp33_ASAP7_75t_L g893 ( 
.A(n_891),
.B(n_772),
.C(n_764),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_892),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_SL g895 ( 
.A1(n_893),
.A2(n_891),
.B(n_748),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_892),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_894),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_SL g898 ( 
.A1(n_896),
.A2(n_759),
.B1(n_779),
.B2(n_773),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_SL g899 ( 
.A1(n_895),
.A2(n_729),
.B(n_734),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_894),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_894),
.Y(n_901)
);

AO22x2_ASAP7_75t_L g902 ( 
.A1(n_897),
.A2(n_776),
.B1(n_729),
.B2(n_734),
.Y(n_902)
);

OAI21x1_ASAP7_75t_SL g903 ( 
.A1(n_900),
.A2(n_803),
.B(n_736),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_901),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_899),
.A2(n_769),
.B(n_760),
.Y(n_905)
);

OAI21xp33_ASAP7_75t_L g906 ( 
.A1(n_898),
.A2(n_776),
.B(n_775),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_897),
.Y(n_907)
);

XNOR2xp5_ASAP7_75t_L g908 ( 
.A(n_904),
.B(n_761),
.Y(n_908)
);

AOI31xp33_ASAP7_75t_L g909 ( 
.A1(n_906),
.A2(n_794),
.A3(n_799),
.B(n_802),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_907),
.A2(n_772),
.B(n_764),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_908),
.B(n_903),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_911),
.A2(n_910),
.B(n_902),
.Y(n_912)
);

AOI211xp5_ASAP7_75t_L g913 ( 
.A1(n_912),
.A2(n_905),
.B(n_909),
.C(n_799),
.Y(n_913)
);


endmodule