module fake_jpeg_1198_n_451 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_451);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_451;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_55),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_56),
.B(n_57),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_16),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_60),
.B(n_62),
.Y(n_167)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_13),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_63),
.Y(n_158)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_64),
.Y(n_179)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_65),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_33),
.B(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_66),
.B(n_82),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_74),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_33),
.B(n_13),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_75),
.B(n_84),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_79),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_22),
.A2(n_11),
.B(n_2),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_80),
.B(n_6),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_18),
.B(n_0),
.C(n_2),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_34),
.B(n_0),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_87),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_34),
.B(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_88),
.B(n_89),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_3),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_47),
.B(n_6),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_94),
.B(n_109),
.Y(n_183)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_47),
.B(n_53),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_103),
.B(n_106),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_6),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_37),
.B(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_25),
.B(n_10),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_110),
.B(n_91),
.Y(n_190)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_28),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_114),
.Y(n_142)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_116),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_74),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_117),
.B(n_191),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_64),
.B(n_37),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_122),
.B(n_135),
.Y(n_215)
);

NAND4xp25_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_42),
.C(n_45),
.D(n_54),
.Y(n_126)
);

NAND4xp25_ASAP7_75t_L g249 ( 
.A(n_126),
.B(n_110),
.C(n_184),
.D(n_189),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_52),
.B1(n_42),
.B2(n_23),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_128),
.A2(n_140),
.B1(n_181),
.B2(n_187),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_27),
.B1(n_23),
.B2(n_52),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g209 ( 
.A1(n_133),
.A2(n_134),
.B1(n_147),
.B2(n_149),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_87),
.A2(n_27),
.B1(n_69),
.B2(n_58),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_93),
.B(n_21),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_67),
.A2(n_27),
.B1(n_45),
.B2(n_54),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_96),
.B(n_21),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_144),
.B(n_146),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_97),
.B(n_19),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_55),
.A2(n_19),
.B1(n_28),
.B2(n_44),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_55),
.A2(n_28),
.B1(n_44),
.B2(n_40),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_71),
.A2(n_25),
.B1(n_36),
.B2(n_32),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_150),
.A2(n_170),
.B1(n_155),
.B2(n_171),
.Y(n_226)
);

AO22x1_ASAP7_75t_L g155 ( 
.A1(n_61),
.A2(n_40),
.B1(n_36),
.B2(n_32),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_150),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_157),
.B(n_190),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_58),
.A2(n_30),
.B1(n_8),
.B2(n_9),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g229 ( 
.A1(n_166),
.A2(n_185),
.B1(n_125),
.B2(n_162),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_73),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_112),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_69),
.A2(n_65),
.B1(n_92),
.B2(n_86),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_98),
.A2(n_7),
.B1(n_10),
.B2(n_108),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_101),
.A2(n_10),
.B1(n_104),
.B2(n_102),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_188),
.A2(n_174),
.B1(n_186),
.B2(n_193),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_76),
.B(n_83),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_79),
.B(n_81),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_142),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_139),
.Y(n_196)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_196),
.Y(n_298)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_198),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_199),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_200),
.Y(n_272)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_123),
.B(n_163),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_206),
.Y(n_268)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

BUFx2_ASAP7_75t_SL g204 ( 
.A(n_153),
.Y(n_204)
);

BUFx8_ASAP7_75t_L g280 ( 
.A(n_204),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_151),
.B1(n_121),
.B2(n_143),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_205),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_207),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_154),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_208),
.B(n_213),
.Y(n_269)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_210),
.Y(n_293)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_211),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_192),
.A2(n_140),
.B1(n_133),
.B2(n_185),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_212),
.A2(n_219),
.B1(n_226),
.B2(n_237),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_124),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_216),
.B(n_217),
.Y(n_271)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_167),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_218),
.B(n_220),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_136),
.A2(n_161),
.B1(n_149),
.B2(n_147),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_175),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_221),
.B(n_223),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_180),
.A2(n_166),
.B(n_134),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_222),
.A2(n_209),
.B(n_229),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_137),
.B(n_178),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_224),
.B(n_225),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_148),
.B(n_160),
.Y(n_225)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_129),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_227),
.A2(n_229),
.B1(n_233),
.B2(n_234),
.Y(n_285)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_138),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_228),
.B(n_230),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_124),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_170),
.B(n_145),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_238),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_156),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_232),
.B(n_235),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_131),
.A2(n_158),
.B1(n_118),
.B2(n_182),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_138),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_119),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_176),
.B(n_174),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_130),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_119),
.B(n_130),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_244),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g243 ( 
.A1(n_152),
.A2(n_171),
.B1(n_164),
.B2(n_186),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_243),
.A2(n_245),
.B1(n_236),
.B2(n_212),
.Y(n_273)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_152),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_164),
.A2(n_190),
.B1(n_192),
.B2(n_163),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_127),
.B(n_168),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_247),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_127),
.B(n_168),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_128),
.A2(n_114),
.B1(n_48),
.B2(n_27),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_248),
.A2(n_254),
.B1(n_195),
.B2(n_207),
.Y(n_300)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_250),
.B(n_200),
.C(n_194),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_252),
.Y(n_292)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_156),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_156),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_256),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_122),
.B(n_184),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_120),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_255),
.B(n_257),
.Y(n_294)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_139),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_124),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_226),
.A2(n_200),
.B1(n_231),
.B2(n_245),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_258),
.A2(n_273),
.B1(n_275),
.B2(n_282),
.Y(n_307)
);

AND2x2_ASAP7_75t_SL g263 ( 
.A(n_242),
.B(n_215),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_263),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_267),
.B(n_276),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_239),
.A2(n_254),
.B1(n_209),
.B2(n_219),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_210),
.B(n_223),
.C(n_222),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_301),
.C(n_281),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_209),
.A2(n_225),
.B1(n_229),
.B2(n_221),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_284),
.A2(n_303),
.B(n_285),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_209),
.A2(n_229),
.B1(n_224),
.B2(n_211),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_287),
.A2(n_296),
.B1(n_302),
.B2(n_304),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_243),
.A2(n_256),
.B1(n_196),
.B2(n_214),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_299),
.B1(n_286),
.B2(n_260),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_198),
.A2(n_203),
.B1(n_216),
.B2(n_228),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_244),
.A2(n_234),
.B1(n_227),
.B2(n_201),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_238),
.B(n_253),
.C(n_252),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_217),
.A2(n_249),
.B1(n_197),
.B2(n_255),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_L g303 ( 
.A(n_251),
.B(n_235),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_226),
.A2(n_200),
.B1(n_231),
.B2(n_245),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_270),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_308),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_270),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g309 ( 
.A1(n_284),
.A2(n_273),
.B(n_272),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_309),
.B(n_319),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_262),
.A2(n_272),
.B1(n_275),
.B2(n_304),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_310),
.A2(n_332),
.B1(n_336),
.B2(n_340),
.Y(n_345)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_268),
.B(n_274),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_312),
.B(n_322),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_313),
.A2(n_320),
.B(n_331),
.Y(n_347)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_261),
.B(n_305),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_316),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_298),
.C(n_264),
.Y(n_346)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

O2A1O1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_287),
.A2(n_278),
.B(n_282),
.C(n_261),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_258),
.B(n_279),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_321),
.B(n_328),
.Y(n_362)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_293),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_323),
.Y(n_360)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_260),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_324),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_269),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_325),
.B(n_326),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_279),
.B(n_267),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_263),
.B(n_290),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_259),
.B(n_294),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_263),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_259),
.B(n_263),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_333),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_303),
.A2(n_295),
.B(n_283),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_262),
.A2(n_289),
.B1(n_295),
.B2(n_291),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_301),
.Y(n_333)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_302),
.B(n_292),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_337),
.A2(n_338),
.B(n_341),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_265),
.B(n_281),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_265),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_339),
.A2(n_286),
.B(n_297),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_266),
.A2(n_271),
.B1(n_299),
.B2(n_277),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_280),
.A2(n_264),
.B(n_297),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_277),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_342),
.B(n_343),
.C(n_346),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_280),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_344),
.Y(n_369)
);

AOI322xp5_ASAP7_75t_L g348 ( 
.A1(n_322),
.A2(n_266),
.A3(n_280),
.B1(n_296),
.B2(n_298),
.C1(n_326),
.C2(n_309),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_348),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_307),
.A2(n_321),
.B1(n_334),
.B2(n_314),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_352),
.A2(n_316),
.B1(n_336),
.B2(n_323),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_317),
.C(n_333),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_354),
.B(n_361),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_320),
.A2(n_310),
.B(n_307),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_357),
.A2(n_335),
.B(n_347),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_332),
.A2(n_334),
.B1(n_315),
.B2(n_337),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_358),
.A2(n_311),
.B1(n_335),
.B2(n_345),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_317),
.B(n_306),
.C(n_308),
.Y(n_361)
);

OAI22x1_ASAP7_75t_L g364 ( 
.A1(n_320),
.A2(n_316),
.B1(n_325),
.B2(n_327),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_364),
.A2(n_338),
.B1(n_324),
.B2(n_319),
.Y(n_372)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_355),
.Y(n_366)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_352),
.A2(n_340),
.B1(n_316),
.B2(n_328),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_367),
.A2(n_368),
.B1(n_353),
.B2(n_362),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_355),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_371),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g371 ( 
.A1(n_356),
.A2(n_341),
.B(n_339),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_372),
.A2(n_380),
.B(n_347),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_351),
.B(n_312),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_373),
.B(n_384),
.Y(n_392)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_375),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_349),
.Y(n_376)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_376),
.Y(n_393)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_344),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_381),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_379),
.A2(n_368),
.B1(n_383),
.B2(n_381),
.Y(n_400)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_365),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_365),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_383),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_350),
.B(n_362),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_349),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_385),
.B(n_351),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_354),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_388),
.B(n_398),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_374),
.B(n_346),
.C(n_382),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_389),
.B(n_399),
.C(n_402),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_390),
.A2(n_401),
.B(n_376),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_368),
.A2(n_358),
.B1(n_345),
.B2(n_357),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_394),
.A2(n_400),
.B1(n_367),
.B2(n_372),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_356),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_364),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_363),
.C(n_342),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_363),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_404),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_401),
.A2(n_380),
.B(n_385),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_410),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_394),
.A2(n_400),
.B1(n_397),
.B2(n_379),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_406),
.A2(n_372),
.B1(n_393),
.B2(n_387),
.Y(n_422)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_396),
.Y(n_407)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_407),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_359),
.Y(n_408)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_408),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_409),
.A2(n_395),
.B1(n_369),
.B2(n_378),
.Y(n_419)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_391),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_412),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_375),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_402),
.B(n_359),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_414),
.A2(n_415),
.B1(n_416),
.B2(n_389),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_SL g415 ( 
.A(n_395),
.B(n_356),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_373),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_419),
.A2(n_421),
.B1(n_422),
.B2(n_405),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_424),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_406),
.A2(n_369),
.B1(n_377),
.B2(n_387),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_388),
.C(n_398),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_350),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_428),
.Y(n_438)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_417),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_412),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_431),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_424),
.B(n_413),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_432),
.Y(n_436)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_426),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_404),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_434),
.A2(n_429),
.B(n_423),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_433),
.B(n_403),
.C(n_421),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_439),
.Y(n_442)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_432),
.A2(n_415),
.B(n_425),
.C(n_423),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_440),
.A2(n_419),
.B(n_411),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_430),
.C(n_440),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_441),
.B(n_444),
.C(n_391),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_443),
.A2(n_437),
.B(n_393),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_437),
.B(n_438),
.C(n_422),
.Y(n_444)
);

INVxp33_ASAP7_75t_L g448 ( 
.A(n_445),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_446),
.B(n_447),
.C(n_407),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_442),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_449),
.B(n_386),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_448),
.Y(n_451)
);


endmodule