module real_aes_335_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_498;
wire n_481;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
wire n_237;
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_0), .A2(n_204), .B1(n_281), .B2(n_282), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_1), .A2(n_164), .B1(n_266), .B2(n_350), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_2), .A2(n_115), .B1(n_281), .B2(n_282), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_3), .A2(n_131), .B1(n_538), .B2(n_621), .Y(n_620) );
AO22x2_ASAP7_75t_L g255 ( .A1(n_4), .A2(n_150), .B1(n_245), .B2(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g634 ( .A(n_4), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_5), .A2(n_151), .B1(n_304), .B2(n_350), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_6), .A2(n_92), .B1(n_342), .B2(n_345), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_7), .A2(n_208), .B1(n_266), .B2(n_269), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_8), .A2(n_173), .B1(n_333), .B2(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_9), .B(n_605), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_10), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_11), .Y(n_560) );
AO22x2_ASAP7_75t_L g252 ( .A1(n_12), .A2(n_47), .B1(n_245), .B2(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_12), .B(n_633), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_13), .A2(n_184), .B1(n_330), .B2(n_333), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_14), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g646 ( .A1(n_15), .A2(n_66), .B1(n_272), .B2(n_275), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_16), .A2(n_180), .B1(n_294), .B2(n_446), .Y(n_569) );
AO222x2_ASAP7_75t_SL g301 ( .A1(n_17), .A2(n_35), .B1(n_123), .B2(n_241), .C1(n_257), .C2(n_261), .Y(n_301) );
AO22x2_ASAP7_75t_L g510 ( .A1(n_18), .A2(n_511), .B1(n_540), .B2(n_541), .Y(n_510) );
INVx1_ASAP7_75t_L g541 ( .A(n_18), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_19), .A2(n_65), .B1(n_287), .B2(n_345), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_20), .A2(n_46), .B1(n_338), .B2(n_676), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_21), .A2(n_126), .B1(n_285), .B2(n_291), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_22), .A2(n_119), .B1(n_269), .B2(n_304), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_23), .A2(n_161), .B1(n_534), .B2(n_535), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_24), .A2(n_199), .B1(n_272), .B2(n_306), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_25), .A2(n_167), .B1(n_377), .B2(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_26), .A2(n_203), .B1(n_376), .B2(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_27), .A2(n_120), .B1(n_287), .B2(n_290), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_28), .A2(n_175), .B1(n_418), .B2(n_421), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_29), .A2(n_136), .B1(n_668), .B2(n_669), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_30), .A2(n_105), .B1(n_281), .B2(n_282), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_31), .A2(n_146), .B1(n_557), .B2(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_32), .A2(n_129), .B1(n_338), .B2(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_33), .A2(n_109), .B1(n_294), .B2(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_34), .A2(n_95), .B1(n_352), .B2(n_415), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_36), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_37), .A2(n_207), .B1(n_496), .B2(n_498), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_38), .A2(n_148), .B1(n_505), .B2(n_598), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_39), .A2(n_211), .B1(n_579), .B2(n_617), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_40), .A2(n_73), .B1(n_330), .B2(n_678), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_41), .A2(n_93), .B1(n_404), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_42), .A2(n_69), .B1(n_272), .B2(n_306), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_43), .A2(n_210), .B1(n_344), .B2(n_345), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_44), .A2(n_141), .B1(n_527), .B2(n_528), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_45), .A2(n_118), .B1(n_257), .B2(n_261), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_48), .A2(n_162), .B1(n_257), .B2(n_261), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g265 ( .A1(n_49), .A2(n_84), .B1(n_266), .B2(n_269), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_50), .Y(n_406) );
AO222x2_ASAP7_75t_SL g240 ( .A1(n_51), .A2(n_144), .B1(n_160), .B2(n_241), .C1(n_257), .C2(n_261), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_52), .A2(n_181), .B1(n_538), .B2(n_539), .Y(n_537) );
AND2x2_ASAP7_75t_L g477 ( .A(n_53), .B(n_478), .Y(n_477) );
OA22x2_ASAP7_75t_L g547 ( .A1(n_54), .A2(n_548), .B1(n_549), .B2(n_571), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_54), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_55), .A2(n_86), .B1(n_415), .B2(n_671), .Y(n_670) );
INVx3_ASAP7_75t_L g245 ( .A(n_56), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_57), .A2(n_113), .B1(n_293), .B2(n_294), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_58), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_59), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_60), .A2(n_156), .B1(n_285), .B2(n_287), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_61), .A2(n_212), .B1(n_257), .B2(n_261), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_62), .A2(n_174), .B1(n_390), .B2(n_523), .Y(n_522) );
AOI222xp33_ASAP7_75t_L g357 ( .A1(n_63), .A2(n_75), .B1(n_152), .B2(n_358), .C1(n_359), .C2(n_361), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_64), .A2(n_638), .B1(n_655), .B2(n_656), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_64), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_67), .A2(n_202), .B1(n_281), .B2(n_282), .Y(n_570) );
INVx1_ASAP7_75t_SL g246 ( .A(n_68), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_68), .B(n_103), .Y(n_635) );
AO22x1_ASAP7_75t_L g480 ( .A1(n_70), .A2(n_127), .B1(n_383), .B2(n_481), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_71), .A2(n_209), .B1(n_523), .B2(n_593), .Y(n_592) );
AOI22xp5_ASAP7_75t_SL g614 ( .A1(n_72), .A2(n_171), .B1(n_598), .B2(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g228 ( .A(n_74), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_76), .B(n_438), .Y(n_437) );
XOR2x2_ASAP7_75t_L g574 ( .A(n_77), .B(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_78), .A2(n_172), .B1(n_272), .B2(n_275), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_79), .Y(n_369) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_80), .A2(n_223), .B(n_232), .C(n_636), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_81), .A2(n_107), .B1(n_257), .B2(n_361), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_82), .A2(n_117), .B1(n_293), .B2(n_294), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_83), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_85), .A2(n_112), .B1(n_505), .B2(n_506), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_87), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_88), .A2(n_98), .B1(n_404), .B2(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_89), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_90), .A2(n_143), .B1(n_281), .B2(n_282), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_91), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_94), .A2(n_200), .B1(n_352), .B2(n_355), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_96), .A2(n_153), .B1(n_287), .B2(n_290), .Y(n_443) );
INVx1_ASAP7_75t_L g472 ( .A(n_97), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_99), .A2(n_215), .B1(n_508), .B2(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_100), .A2(n_216), .B1(n_583), .B2(n_585), .Y(n_582) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_101), .A2(n_138), .B1(n_281), .B2(n_282), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_102), .A2(n_154), .B1(n_506), .B2(n_596), .Y(n_595) );
AO22x2_ASAP7_75t_L g248 ( .A1(n_103), .A2(n_163), .B1(n_245), .B2(n_249), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_104), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_106), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_108), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_110), .A2(n_195), .B1(n_530), .B2(n_531), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_111), .A2(n_178), .B1(n_287), .B2(n_290), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_114), .A2(n_125), .B1(n_266), .B2(n_269), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_116), .A2(n_221), .B1(n_323), .B2(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g247 ( .A(n_121), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_122), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_124), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_128), .A2(n_145), .B1(n_282), .B2(n_674), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_130), .A2(n_179), .B1(n_338), .B2(n_340), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_132), .A2(n_183), .B1(n_578), .B2(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g601 ( .A(n_133), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_134), .A2(n_137), .B1(n_293), .B2(n_294), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_135), .A2(n_149), .B1(n_611), .B2(n_612), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_139), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_140), .A2(n_193), .B1(n_287), .B2(n_290), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_142), .A2(n_168), .B1(n_345), .B2(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_147), .A2(n_198), .B1(n_285), .B2(n_291), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_155), .A2(n_158), .B1(n_290), .B2(n_291), .Y(n_289) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_157), .A2(n_165), .B1(n_272), .B2(n_275), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_159), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_166), .A2(n_190), .B1(n_418), .B2(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_169), .B(n_453), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_170), .B(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_L g230 ( .A(n_176), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g630 ( .A(n_176), .Y(n_630) );
AO21x1_ASAP7_75t_L g684 ( .A1(n_176), .A2(n_226), .B(n_685), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g643 ( .A(n_177), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_182), .A2(n_188), .B1(n_345), .B2(n_412), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_185), .A2(n_213), .B1(n_377), .B2(n_586), .Y(n_666) );
INVx1_ASAP7_75t_L g231 ( .A(n_186), .Y(n_231) );
AND2x2_ASAP7_75t_R g658 ( .A(n_186), .B(n_630), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_187), .B(n_358), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_189), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_191), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_192), .B(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_194), .A2(n_219), .B1(n_290), .B2(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_L g227 ( .A(n_196), .Y(n_227) );
XNOR2x1_ASAP7_75t_L g662 ( .A(n_197), .B(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_L g686 ( .A(n_197), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_201), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_205), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_206), .A2(n_218), .B1(n_293), .B2(n_294), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_214), .B(n_453), .Y(n_452) );
OA22x2_ASAP7_75t_L g318 ( .A1(n_217), .A2(n_319), .B1(n_320), .B2(n_362), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_217), .Y(n_319) );
AO21x2_ASAP7_75t_L g426 ( .A1(n_217), .A2(n_320), .B(n_427), .Y(n_426) );
AOI22x1_ASAP7_75t_L g237 ( .A1(n_220), .A2(n_238), .B1(n_295), .B2(n_296), .Y(n_237) );
INVx1_ASAP7_75t_L g296 ( .A(n_220), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_229), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVxp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_231), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g685 ( .A(n_231), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_543), .B1(n_625), .B2(n_626), .C(n_627), .Y(n_232) );
INVx1_ASAP7_75t_L g625 ( .A(n_233), .Y(n_625) );
XOR2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_430), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_316), .B1(n_317), .B2(n_429), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g429 ( .A(n_236), .Y(n_429) );
AO22x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_297), .B1(n_298), .B2(n_315), .Y(n_236) );
INVx1_ASAP7_75t_L g315 ( .A(n_237), .Y(n_315) );
INVx1_ASAP7_75t_L g295 ( .A(n_238), .Y(n_295) );
NAND2x1_ASAP7_75t_SL g238 ( .A(n_239), .B(n_278), .Y(n_238) );
NOR2xp67_ASAP7_75t_L g239 ( .A(n_240), .B(n_264), .Y(n_239) );
BUFx2_ASAP7_75t_L g358 ( .A(n_241), .Y(n_358) );
INVx2_ASAP7_75t_SL g642 ( .A(n_241), .Y(n_642) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_250), .Y(n_241) );
AND2x2_ASAP7_75t_L g269 ( .A(n_242), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g275 ( .A(n_242), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g306 ( .A(n_242), .B(n_276), .Y(n_306) );
AND2x2_ASAP7_75t_L g350 ( .A(n_242), .B(n_270), .Y(n_350) );
AND2x4_ASAP7_75t_L g356 ( .A(n_242), .B(n_276), .Y(n_356) );
AND2x2_ASAP7_75t_L g374 ( .A(n_242), .B(n_250), .Y(n_374) );
AND2x4_ASAP7_75t_L g423 ( .A(n_242), .B(n_270), .Y(n_423) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_248), .Y(n_242) );
AND2x2_ASAP7_75t_L g259 ( .A(n_243), .B(n_260), .Y(n_259) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_243), .Y(n_262) );
INVx2_ASAP7_75t_L g268 ( .A(n_243), .Y(n_268) );
OAI22x1_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B1(n_246), .B2(n_247), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g249 ( .A(n_245), .Y(n_249) );
INVx2_ASAP7_75t_L g253 ( .A(n_245), .Y(n_253) );
INVx1_ASAP7_75t_L g256 ( .A(n_245), .Y(n_256) );
INVx2_ASAP7_75t_L g260 ( .A(n_248), .Y(n_260) );
AND2x2_ASAP7_75t_L g267 ( .A(n_248), .B(n_268), .Y(n_267) );
BUFx2_ASAP7_75t_L g283 ( .A(n_248), .Y(n_283) );
AND2x2_ASAP7_75t_L g285 ( .A(n_250), .B(n_286), .Y(n_285) );
AND2x6_ASAP7_75t_L g290 ( .A(n_250), .B(n_267), .Y(n_290) );
AND2x2_ASAP7_75t_L g293 ( .A(n_250), .B(n_259), .Y(n_293) );
AND2x2_ASAP7_75t_L g332 ( .A(n_250), .B(n_267), .Y(n_332) );
AND2x4_ASAP7_75t_L g339 ( .A(n_250), .B(n_259), .Y(n_339) );
AND2x4_ASAP7_75t_L g347 ( .A(n_250), .B(n_286), .Y(n_347) );
AND2x2_ASAP7_75t_L g446 ( .A(n_250), .B(n_259), .Y(n_446) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_254), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g258 ( .A(n_252), .B(n_254), .Y(n_258) );
AND2x2_ASAP7_75t_L g263 ( .A(n_252), .B(n_255), .Y(n_263) );
INVx1_ASAP7_75t_L g274 ( .A(n_252), .Y(n_274) );
INVxp67_ASAP7_75t_L g270 ( .A(n_254), .Y(n_270) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g273 ( .A(n_255), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_SL g360 ( .A(n_257), .Y(n_360) );
AND2x4_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_L g266 ( .A(n_258), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g291 ( .A(n_258), .B(n_286), .Y(n_291) );
AND2x2_ASAP7_75t_L g304 ( .A(n_258), .B(n_267), .Y(n_304) );
AND2x4_ASAP7_75t_L g342 ( .A(n_258), .B(n_286), .Y(n_342) );
AND2x2_ASAP7_75t_L g378 ( .A(n_258), .B(n_259), .Y(n_378) );
AND2x4_ASAP7_75t_L g420 ( .A(n_258), .B(n_267), .Y(n_420) );
AND2x4_ASAP7_75t_L g272 ( .A(n_259), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g354 ( .A(n_259), .B(n_273), .Y(n_354) );
AND2x4_ASAP7_75t_L g286 ( .A(n_260), .B(n_268), .Y(n_286) );
AND2x2_ASAP7_75t_SL g261 ( .A(n_262), .B(n_263), .Y(n_261) );
AND2x2_ASAP7_75t_SL g361 ( .A(n_262), .B(n_263), .Y(n_361) );
AND2x2_ASAP7_75t_L g384 ( .A(n_262), .B(n_263), .Y(n_384) );
AND2x4_ASAP7_75t_L g282 ( .A(n_263), .B(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g294 ( .A(n_263), .B(n_286), .Y(n_294) );
AND2x4_ASAP7_75t_L g328 ( .A(n_263), .B(n_283), .Y(n_328) );
AND2x4_ASAP7_75t_L g344 ( .A(n_263), .B(n_286), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_271), .Y(n_264) );
AND2x2_ASAP7_75t_SL g281 ( .A(n_267), .B(n_273), .Y(n_281) );
AND2x2_ASAP7_75t_L g325 ( .A(n_267), .B(n_273), .Y(n_325) );
AND2x2_ASAP7_75t_L g674 ( .A(n_267), .B(n_273), .Y(n_674) );
INVxp67_ASAP7_75t_L g563 ( .A(n_269), .Y(n_563) );
AND2x6_ASAP7_75t_L g287 ( .A(n_273), .B(n_286), .Y(n_287) );
AND2x4_ASAP7_75t_L g335 ( .A(n_273), .B(n_286), .Y(n_335) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_274), .Y(n_277) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2x1_ASAP7_75t_L g278 ( .A(n_279), .B(n_288), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_284), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
XOR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_314), .Y(n_298) );
NAND2x1_ASAP7_75t_L g299 ( .A(n_300), .B(n_307), .Y(n_299) );
NOR2x1_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVxp67_ASAP7_75t_L g561 ( .A(n_304), .Y(n_561) );
NOR2x1_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_363), .B1(n_364), .B2(n_425), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_319), .Y(n_428) );
INVx1_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
NOR2x1_ASAP7_75t_SL g427 ( .A(n_320), .B(n_428), .Y(n_427) );
NAND4xp75_ASAP7_75t_L g320 ( .A(n_321), .B(n_336), .C(n_348), .D(n_357), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_329), .Y(n_321) );
INVx1_ASAP7_75t_L g497 ( .A(n_323), .Y(n_497) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g594 ( .A(n_324), .Y(n_594) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_325), .Y(n_390) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_327), .A2(n_387), .B1(n_388), .B2(n_391), .Y(n_386) );
INVx2_ASAP7_75t_L g498 ( .A(n_327), .Y(n_498) );
INVx5_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g523 ( .A(n_328), .Y(n_523) );
BUFx3_ASAP7_75t_L g612 ( .A(n_328), .Y(n_612) );
INVx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g396 ( .A(n_331), .Y(n_396) );
INVx2_ASAP7_75t_SL g505 ( .A(n_331), .Y(n_505) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx2_ASAP7_75t_L g538 ( .A(n_332), .Y(n_538) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_334), .A2(n_393), .B1(n_394), .B2(n_397), .Y(n_392) );
INVx2_ASAP7_75t_L g539 ( .A(n_334), .Y(n_539) );
INVx2_ASAP7_75t_L g598 ( .A(n_334), .Y(n_598) );
INVx2_ASAP7_75t_L g680 ( .A(n_334), .Y(n_680) );
INVx8_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_343), .Y(n_336) );
BUFx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx6_ASAP7_75t_L g401 ( .A(n_339), .Y(n_401) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_340), .Y(n_621) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g465 ( .A(n_341), .Y(n_465) );
INVx1_ASAP7_75t_L g678 ( .A(n_341), .Y(n_678) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_342), .Y(n_412) );
BUFx3_ASAP7_75t_L g521 ( .A(n_342), .Y(n_521) );
BUFx2_ASAP7_75t_SL g404 ( .A(n_344), .Y(n_404) );
INVx2_ASAP7_75t_L g536 ( .A(n_344), .Y(n_536) );
BUFx2_ASAP7_75t_SL g591 ( .A(n_344), .Y(n_591) );
BUFx3_ASAP7_75t_L g676 ( .A(n_344), .Y(n_676) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_SL g409 ( .A(n_346), .Y(n_409) );
INVx4_ASAP7_75t_L g502 ( .A(n_346), .Y(n_502) );
INVx2_ASAP7_75t_SL g534 ( .A(n_346), .Y(n_534) );
INVx2_ASAP7_75t_L g615 ( .A(n_346), .Y(n_615) );
INVx8_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx2_ASAP7_75t_SL g485 ( .A(n_352), .Y(n_485) );
INVx4_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g531 ( .A(n_353), .Y(n_531) );
INVx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_354), .Y(n_557) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_354), .Y(n_671) );
BUFx6f_ASAP7_75t_SL g607 ( .A(n_355), .Y(n_607) );
BUFx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g416 ( .A(n_356), .Y(n_416) );
INVx2_ASAP7_75t_L g488 ( .A(n_356), .Y(n_488) );
BUFx6f_ASAP7_75t_SL g530 ( .A(n_356), .Y(n_530) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
XNOR2x1_ASAP7_75t_L g365 ( .A(n_366), .B(n_424), .Y(n_365) );
NAND4xp75_ASAP7_75t_L g366 ( .A(n_367), .B(n_385), .C(n_398), .D(n_413), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_375), .B2(n_379), .C(n_380), .Y(n_368) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g514 ( .A(n_372), .Y(n_514) );
INVx3_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx4_ASAP7_75t_SL g438 ( .A(n_373), .Y(n_438) );
INVx4_ASAP7_75t_SL g453 ( .A(n_373), .Y(n_453) );
BUFx2_ASAP7_75t_L g479 ( .A(n_373), .Y(n_479) );
INVx3_ASAP7_75t_L g605 ( .A(n_373), .Y(n_605) );
INVx6_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g482 ( .A(n_378), .Y(n_482) );
BUFx3_ASAP7_75t_L g584 ( .A(n_378), .Y(n_584) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g619 ( .A(n_383), .Y(n_619) );
BUFx12f_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx3_ASAP7_75t_L g518 ( .A(n_384), .Y(n_518) );
NOR2x1_ASAP7_75t_L g385 ( .A(n_386), .B(n_392), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_405), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_399) );
INVx2_ASAP7_75t_L g508 ( .A(n_401), .Y(n_508) );
INVx2_ASAP7_75t_L g609 ( .A(n_401), .Y(n_609) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B1(n_410), .B2(n_411), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_412), .Y(n_506) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_417), .Y(n_413) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_416), .A2(n_555), .B1(n_556), .B2(n_558), .Y(n_554) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g491 ( .A(n_419), .Y(n_491) );
BUFx2_ASAP7_75t_L g578 ( .A(n_419), .Y(n_578) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx3_ASAP7_75t_L g527 ( .A(n_420), .Y(n_527) );
BUFx2_ASAP7_75t_L g668 ( .A(n_420), .Y(n_668) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_422), .A2(n_490), .B1(n_491), .B2(n_492), .Y(n_489) );
INVx2_ASAP7_75t_SL g528 ( .A(n_422), .Y(n_528) );
INVx2_ASAP7_75t_L g579 ( .A(n_422), .Y(n_579) );
INVx2_ASAP7_75t_SL g669 ( .A(n_422), .Y(n_669) );
INVx6_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_467), .B1(n_468), .B2(n_542), .Y(n_430) );
INVx1_ASAP7_75t_L g542 ( .A(n_431), .Y(n_542) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
XNOR2x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_448), .Y(n_432) );
XNOR2x1_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
NOR2x1_ASAP7_75t_L g435 ( .A(n_436), .B(n_442), .Y(n_435) );
NAND4xp25_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .C(n_440), .D(n_441), .Y(n_436) );
NAND4xp25_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .C(n_445), .D(n_447), .Y(n_442) );
XOR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_466), .Y(n_448) );
NAND2x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_458), .Y(n_449) );
NOR2x1_ASAP7_75t_L g450 ( .A(n_451), .B(n_455), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
BUFx2_ASAP7_75t_L g581 ( .A(n_453), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
NOR2x1_ASAP7_75t_L g458 ( .A(n_459), .B(n_462), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
XNOR2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_510), .Y(n_470) );
OAI21x1_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_509), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_472), .B(n_475), .Y(n_509) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_493), .Y(n_475) );
NOR4xp75_ASAP7_75t_L g476 ( .A(n_477), .B(n_480), .C(n_483), .D(n_489), .Y(n_476) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_486), .B2(n_487), .Y(n_483) );
INVx3_ASAP7_75t_L g588 ( .A(n_487), .Y(n_588) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_499), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g611 ( .A(n_497), .Y(n_611) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_502), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
INVx2_ASAP7_75t_SL g540 ( .A(n_511), .Y(n_540) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_524), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_519), .Y(n_512) );
OAI21xp33_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_515), .B(n_516), .Y(n_513) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g586 ( .A(n_518), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_532), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_529), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_537), .Y(n_532) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g626 ( .A(n_543), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_572), .B1(n_623), .B2(n_624), .Y(n_543) );
INVx1_ASAP7_75t_L g623 ( .A(n_544), .Y(n_623) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g571 ( .A(n_549), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_564), .Y(n_549) );
NOR3xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .C(n_559), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx6f_ASAP7_75t_SL g617 ( .A(n_557), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_562), .B2(n_563), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_568), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g624 ( .A(n_572), .Y(n_624) );
OAI22xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_599), .B1(n_600), .B2(n_622), .Y(n_572) );
INVx3_ASAP7_75t_L g622 ( .A(n_573), .Y(n_622) );
INVx5_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2x1_ASAP7_75t_L g575 ( .A(n_576), .B(n_589), .Y(n_575) );
NAND4xp25_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .C(n_582), .D(n_587), .Y(n_576) );
BUFx6f_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND4xp25_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .C(n_595), .D(n_597), .Y(n_589) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
XNOR2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_603), .B(n_613), .Y(n_602) );
NAND4xp25_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .C(n_608), .D(n_610), .Y(n_603) );
NAND4xp25_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .C(n_618), .D(n_620), .Y(n_613) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_629), .B(n_632), .Y(n_683) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
OAI222xp33_ASAP7_75t_R g636 ( .A1(n_637), .A2(n_657), .B1(n_659), .B2(n_681), .C1(n_684), .C2(n_686), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_638), .Y(n_656) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_640), .B(n_648), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_645), .Y(n_640) );
OAI21xp5_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_643), .B(n_644), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_652), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx3_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_672), .Y(n_663) );
NAND4xp25_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .C(n_667), .D(n_670), .Y(n_664) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .C(n_677), .D(n_679), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_682), .Y(n_681) );
CKINVDCx6p67_ASAP7_75t_R g682 ( .A(n_683), .Y(n_682) );
endmodule