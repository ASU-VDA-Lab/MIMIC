module real_jpeg_16248_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_8),
.B1(n_20),
.B2(n_22),
.Y(n_19)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_1),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_1),
.A2(n_3),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_1),
.Y(n_191)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_2),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_3),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_3),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_3),
.B(n_152),
.Y(n_151)
);

AOI31xp33_ASAP7_75t_SL g187 ( 
.A1(n_3),
.A2(n_124),
.A3(n_188),
.B(n_190),
.Y(n_187)
);

NAND2x1_ASAP7_75t_SL g233 ( 
.A(n_3),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_3),
.B(n_64),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_3),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_3),
.B(n_309),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_4),
.Y(n_173)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_4),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_5),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_6),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_6),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_6),
.B(n_106),
.Y(n_105)
);

NAND2x1_ASAP7_75t_SL g116 ( 
.A(n_6),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_6),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_6),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_6),
.B(n_274),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_7),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_7),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_7),
.B(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g197 ( 
.A(n_9),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_9),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_10),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_10),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_10),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_10),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_10),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_10),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_10),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_11),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_13),
.B(n_55),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_13),
.B(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_14),
.Y(n_87)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_14),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_14),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_15),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_15),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_15),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_15),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_15),
.B(n_93),
.Y(n_283)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_16),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_16),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_16),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_16),
.B(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_17),
.Y(n_139)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g117 ( 
.A(n_18),
.Y(n_117)
);

BUFx12f_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_216),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_180),
.B(n_213),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_25),
.B(n_181),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_112),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_69),
.C(n_96),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_27),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_49),
.C(n_58),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2x1_ASAP7_75t_SL g240 ( 
.A(n_29),
.B(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_30),
.B(n_41),
.C(n_48),
.Y(n_130)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_34),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_48),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_49),
.B(n_58),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_50),
.B(n_54),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_52),
.Y(n_320)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_53),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_57),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_65),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_59),
.A2(n_63),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_59),
.Y(n_225)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_63),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_63),
.B(n_296),
.C(n_298),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_63),
.A2(n_226),
.B1(n_298),
.B2(n_299),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_65),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_67),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_69),
.B(n_96),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_84),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_76),
.B1(n_82),
.B2(n_83),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_71),
.B(n_82),
.C(n_84),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_74),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.C(n_92),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_85),
.B(n_92),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_85),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_85),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_88),
.B(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_100),
.C(n_110),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_105),
.B1(n_110),
.B2(n_111),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_105),
.A2(n_110),
.B1(n_229),
.B2(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_110),
.B(n_229),
.C(n_233),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_147),
.B1(n_178),
.B2(n_179),
.Y(n_112)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_131),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_123),
.C(n_130),
.Y(n_114)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_115),
.B(n_211),
.Y(n_210)
);

XNOR2x2_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_119),
.C(n_122),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_123),
.A2(n_124),
.B1(n_130),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_126),
.B(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_131)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.Y(n_134)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_135),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_331)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_141),
.Y(n_315)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_163),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_158),
.B1(n_159),
.B2(n_162),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_155),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_157),
.Y(n_275)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_210),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_184),
.B(n_210),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_192),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_187),
.Y(n_221)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_202),
.C(n_204),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_193),
.B(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_194),
.B(n_198),
.Y(n_282)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_194),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_194),
.A2(n_307),
.B1(n_308),
.B2(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_244),
.B(n_344),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_242),
.Y(n_218)
);

NOR2x1_ASAP7_75t_L g345 ( 
.A(n_219),
.B(n_242),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.C(n_240),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_220),
.B(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_222),
.B(n_240),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.C(n_238),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_223),
.B(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_228),
.B(n_239),
.Y(n_336)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2x2_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_339),
.B(n_343),
.Y(n_246)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_325),
.B(n_338),
.Y(n_247)
);

OAI21x1_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_290),
.B(n_324),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_278),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_250),
.B(n_278),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_258),
.C(n_267),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_257),
.C(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_258),
.A2(n_259),
.B1(n_267),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_260),
.B(n_264),
.Y(n_297)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_263),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

AO22x1_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_273),
.B1(n_276),
.B2(n_277),
.Y(n_267)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_273),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_276),
.Y(n_280)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_274),
.Y(n_310)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_284),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_279),
.B(n_285),
.C(n_287),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_280),
.B(n_282),
.C(n_283),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

AOI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_301),
.B(n_323),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_295),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_297),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_311),
.B(n_322),
.Y(n_301)
);

NOR2xp67_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_306),
.Y(n_322)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_318),
.B(n_321),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_316),
.Y(n_321)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_337),
.Y(n_325)
);

NOR2x1p5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_337),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_334),
.B2(n_335),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_332),
.B2(n_333),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_333),
.C(n_334),
.Y(n_340)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_340),
.B(n_341),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);


endmodule