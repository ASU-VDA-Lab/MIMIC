module fake_jpeg_29270_n_198 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_1),
.Y(n_73)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_1),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_51),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_29),
.B1(n_22),
.B2(n_21),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_60),
.B1(n_68),
.B2(n_51),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_23),
.B1(n_21),
.B2(n_34),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_67),
.B1(n_71),
.B2(n_72),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_23),
.B1(n_21),
.B2(n_34),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_48),
.B1(n_37),
.B2(n_43),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_22),
.B1(n_23),
.B2(n_34),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_28),
.C(n_32),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_73),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_16),
.B1(n_32),
.B2(n_28),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_37),
.A2(n_16),
.B1(n_26),
.B2(n_30),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_16),
.B1(n_30),
.B2(n_18),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_18),
.B1(n_26),
.B2(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_42),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_86),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_39),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_84),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_88),
.Y(n_102)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_51),
.B1(n_50),
.B2(n_44),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_93),
.B1(n_99),
.B2(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_83),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_39),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_45),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_101),
.B1(n_2),
.B2(n_5),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_24),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_90),
.Y(n_104)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_1),
.Y(n_112)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_33),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_95),
.Y(n_116)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_33),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_97),
.C(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_31),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_31),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_48),
.B1(n_43),
.B2(n_46),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_57),
.A2(n_49),
.B1(n_46),
.B2(n_3),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_70),
.C(n_49),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_107),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_62),
.B(n_55),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_62),
.C(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_112),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_120),
.B1(n_81),
.B2(n_101),
.Y(n_124)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_83),
.B1(n_86),
.B2(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_93),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_123),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_120),
.A2(n_74),
.B1(n_76),
.B2(n_84),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_113),
.B(n_107),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_128),
.B1(n_133),
.B2(n_136),
.Y(n_148)
);

BUFx24_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_76),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_132),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_82),
.B1(n_99),
.B2(n_84),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_80),
.B1(n_78),
.B2(n_77),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_119),
.B1(n_118),
.B2(n_105),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_100),
.B1(n_92),
.B2(n_90),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_115),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_95),
.B1(n_98),
.B2(n_7),
.Y(n_136)
);

AOI322xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_109),
.A3(n_105),
.B1(n_116),
.B2(n_106),
.C1(n_103),
.C2(n_112),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_11),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_127),
.B(n_125),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_132),
.B(n_136),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_147),
.B(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_103),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_150),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_113),
.B1(n_108),
.B2(n_105),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_146),
.A2(n_130),
.B1(n_134),
.B2(n_109),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_113),
.C(n_119),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_129),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_152),
.C(n_153),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_124),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_128),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_159),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_147),
.B1(n_153),
.B2(n_138),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_163),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_5),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_149),
.C(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_164),
.B(n_172),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_169),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_173),
.B(n_162),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_157),
.A2(n_148),
.B1(n_139),
.B2(n_140),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_142),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_152),
.A2(n_148),
.B(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_6),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_167),
.B1(n_159),
.B2(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_177),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_168),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_151),
.B1(n_155),
.B2(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_182),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_170),
.B1(n_164),
.B2(n_171),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_171),
.C(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_187),
.B(n_170),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_189),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_178),
.C(n_179),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_179),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_190),
.A2(n_176),
.B(n_184),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_191),
.A2(n_185),
.B(n_187),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_193),
.A2(n_194),
.B(n_15),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_14),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_14),
.C(n_10),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_10),
.Y(n_198)
);


endmodule