module fake_jpeg_15212_n_382 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_382);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_382;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_40),
.B(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_41),
.B(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_43),
.B(n_18),
.Y(n_80)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_63),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_30),
.B(n_17),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_17),
.B1(n_14),
.B2(n_21),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_67),
.A2(n_71),
.B1(n_115),
.B2(n_101),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_28),
.B1(n_21),
.B2(n_33),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_36),
.B1(n_18),
.B2(n_15),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_74),
.A2(n_84),
.B1(n_95),
.B2(n_99),
.Y(n_125)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_77),
.B(n_85),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_18),
.B1(n_36),
.B2(n_15),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_86),
.B1(n_97),
.B2(n_91),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_91),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_39),
.A2(n_36),
.B1(n_35),
.B2(n_34),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_14),
.B1(n_33),
.B2(n_29),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_43),
.B(n_35),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_65),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_93),
.B(n_77),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_32),
.B1(n_26),
.B2(n_25),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_44),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_45),
.A2(n_32),
.B1(n_26),
.B2(n_25),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_43),
.B(n_31),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_6),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_57),
.A2(n_12),
.B1(n_2),
.B2(n_4),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_111),
.B1(n_114),
.B2(n_73),
.Y(n_133)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_12),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_107),
.B(n_112),
.Y(n_150)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx2_ASAP7_75t_SL g141 ( 
.A(n_108),
.Y(n_141)
);

BUFx8_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_62),
.B(n_31),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_12),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_113),
.B(n_9),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_42),
.A2(n_52),
.B1(n_51),
.B2(n_31),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_110),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_116),
.B(n_118),
.Y(n_174)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_121),
.B(n_165),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_78),
.A2(n_59),
.B1(n_46),
.B2(n_31),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_123),
.A2(n_135),
.B1(n_161),
.B2(n_159),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_131),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_31),
.B(n_20),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_127),
.A2(n_146),
.B(n_159),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_78),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_138),
.Y(n_185)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_88),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_134),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_139),
.B1(n_166),
.B2(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_46),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_76),
.B(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_136),
.B(n_156),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_70),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_46),
.B1(n_7),
.B2(n_8),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

BUFx2_ASAP7_75t_SL g170 ( 
.A(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_109),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_87),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_144),
.B(n_154),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_70),
.A2(n_6),
.B(n_9),
.Y(n_146)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_153),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_87),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_73),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_158),
.A2(n_162),
.B1(n_117),
.B2(n_120),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_75),
.A2(n_10),
.B(n_11),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_101),
.A2(n_10),
.B1(n_11),
.B2(n_93),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_162),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_68),
.A2(n_90),
.B(n_96),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_164),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_125),
.A2(n_109),
.B1(n_81),
.B2(n_83),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_169),
.B(n_182),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_92),
.C(n_106),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_171),
.B(n_186),
.C(n_194),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_172),
.A2(n_188),
.B1(n_207),
.B2(n_209),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_176),
.A2(n_201),
.B(n_185),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_137),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_121),
.B(n_68),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_132),
.A2(n_81),
.B1(n_83),
.B2(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_128),
.B(n_146),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_128),
.B(n_134),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_155),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_128),
.C(n_150),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_201),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_152),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_211),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_129),
.A2(n_138),
.B1(n_158),
.B2(n_141),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_137),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_202),
.B(n_210),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_149),
.A2(n_153),
.B1(n_151),
.B2(n_160),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_208),
.A2(n_180),
.B1(n_173),
.B2(n_195),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_147),
.A2(n_130),
.B1(n_148),
.B2(n_140),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_119),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_164),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_119),
.B(n_145),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_202),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_213),
.B(n_220),
.Y(n_261)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_124),
.B1(n_118),
.B2(n_126),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_215),
.A2(n_244),
.B1(n_253),
.B2(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_168),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_217),
.A2(n_218),
.B(n_229),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_124),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_175),
.Y(n_220)
);

BUFx12_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_231),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_190),
.B(n_186),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_225),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_211),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_226),
.B(n_227),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_204),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_178),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_233),
.A2(n_242),
.B(n_250),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_195),
.B1(n_209),
.B2(n_179),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_189),
.B(n_200),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_235),
.B(n_245),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_177),
.C(n_176),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_232),
.C(n_239),
.Y(n_256)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_181),
.A2(n_172),
.B1(n_177),
.B2(n_171),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_239),
.A2(n_232),
.B1(n_229),
.B2(n_224),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_178),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_176),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_249),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_185),
.A2(n_208),
.B1(n_192),
.B2(n_184),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_196),
.B(n_210),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_184),
.Y(n_247)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_193),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_182),
.B(n_192),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_183),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_183),
.A2(n_191),
.B(n_206),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_251),
.B(n_252),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_207),
.A2(n_191),
.B(n_206),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_252),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_254),
.A2(n_274),
.B(n_273),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_255),
.B(n_256),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_257),
.A2(n_274),
.B1(n_286),
.B2(n_280),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_243),
.A2(n_244),
.B1(n_221),
.B2(n_219),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_258),
.A2(n_264),
.B1(n_266),
.B2(n_273),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_221),
.A2(n_236),
.B1(n_216),
.B2(n_237),
.Y(n_264)
);

XOR2x2_ASAP7_75t_L g265 ( 
.A(n_217),
.B(n_235),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_269),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_236),
.B1(n_240),
.B2(n_217),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_222),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_270),
.B(n_277),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_241),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_272),
.B(n_213),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_234),
.A2(n_228),
.B1(n_218),
.B2(n_238),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_215),
.B(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_218),
.B(n_251),
.C(n_250),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_249),
.C(n_220),
.Y(n_288)
);

AND2x6_ASAP7_75t_L g281 ( 
.A(n_231),
.B(n_245),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_281),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_225),
.A2(n_247),
.B1(n_230),
.B2(n_233),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_282),
.A2(n_242),
.B1(n_246),
.B2(n_223),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_301),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_289),
.B(n_294),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_279),
.Y(n_291)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_261),
.Y(n_292)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_223),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_295),
.B(n_296),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_263),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_297),
.Y(n_330)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_263),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_299),
.A2(n_302),
.B(n_307),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_223),
.C(n_256),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_259),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_306),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_274),
.B1(n_276),
.B2(n_265),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_258),
.B1(n_260),
.B2(n_254),
.Y(n_318)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_268),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_267),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_313),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_310),
.A2(n_292),
.B1(n_307),
.B2(n_306),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_311),
.A2(n_314),
.B(n_271),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_284),
.B(n_259),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_260),
.B(n_284),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_267),
.B(n_269),
.C(n_266),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_271),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_318),
.A2(n_326),
.B1(n_333),
.B2(n_287),
.Y(n_340)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_320),
.Y(n_339)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_305),
.A2(n_285),
.B1(n_278),
.B2(n_283),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_311),
.A2(n_285),
.B(n_283),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_327),
.A2(n_329),
.B(n_304),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_291),
.A2(n_305),
.B(n_313),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_301),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_325),
.C(n_322),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_298),
.A2(n_302),
.B1(n_288),
.B2(n_297),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_335),
.A2(n_290),
.B(n_308),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_336),
.A2(n_343),
.B(n_320),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_317),
.A2(n_287),
.B1(n_303),
.B2(n_310),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_SL g359 ( 
.A1(n_337),
.A2(n_342),
.B(n_341),
.C(n_340),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_309),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_344),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_340),
.B(n_345),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_341),
.A2(n_347),
.B(n_348),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_330),
.A2(n_300),
.B1(n_308),
.B2(n_321),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_315),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_331),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_350),
.Y(n_362)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_334),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_329),
.B(n_333),
.C(n_316),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_352),
.C(n_328),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_326),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_335),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_351),
.B(n_324),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_316),
.B(n_327),
.C(n_332),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_353),
.B(n_355),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_339),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_354),
.A2(n_359),
.B1(n_352),
.B2(n_349),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_356),
.A2(n_358),
.B(n_359),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_328),
.C(n_346),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_358),
.B(n_363),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_342),
.Y(n_363)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_364),
.Y(n_372)
);

AOI221xp5_ASAP7_75t_L g365 ( 
.A1(n_361),
.A2(n_337),
.B1(n_350),
.B2(n_359),
.C(n_354),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_365),
.A2(n_356),
.B1(n_359),
.B2(n_362),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_357),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_362),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_360),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_370),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_371),
.B(n_373),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_375),
.B(n_371),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_376),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_374),
.B(n_372),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_368),
.C(n_369),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_370),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_377),
.C(n_360),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_365),
.Y(n_382)
);


endmodule