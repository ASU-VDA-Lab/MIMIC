module fake_jpeg_20049_n_154 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_10),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_9),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_22),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_16),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_79),
.Y(n_85)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_82),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_83),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_73),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_76),
.B1(n_49),
.B2(n_59),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_94),
.B1(n_95),
.B2(n_61),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_66),
.C(n_67),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_91),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_65),
.B1(n_68),
.B2(n_63),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_63),
.B1(n_57),
.B2(n_72),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_75),
.B1(n_48),
.B2(n_50),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_75),
.B1(n_48),
.B2(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_103),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_101),
.B1(n_105),
.B2(n_55),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_1),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_85),
.B1(n_88),
.B2(n_93),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_107),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_73),
.B1(n_71),
.B2(n_70),
.Y(n_105)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_0),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_58),
.C(n_53),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_120),
.C(n_2),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_51),
.B1(n_64),
.B2(n_52),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_116),
.B1(n_122),
.B2(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_121),
.Y(n_126)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_14),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_124),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_18),
.C(n_43),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_0),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_13),
.B1(n_42),
.B2(n_40),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_12),
.B1(n_39),
.B2(n_34),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_128),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_44),
.B(n_32),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_129),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_112),
.B(n_2),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_3),
.B(n_4),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_131),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_23),
.C(n_21),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_122),
.C(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_139),
.Y(n_142)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_143),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_142),
.B1(n_128),
.B2(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_138),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_126),
.B1(n_136),
.B2(n_140),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_147),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_148),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_149),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_137),
.A3(n_20),
.B1(n_19),
.B2(n_131),
.C1(n_119),
.C2(n_4),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_151),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_5),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_5),
.Y(n_154)
);


endmodule