module fake_jpeg_23966_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_17),
.Y(n_66)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_42),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_9),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_29),
.Y(n_65)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_33),
.B1(n_16),
.B2(n_28),
.Y(n_67)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_59),
.B(n_75),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_21),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_61),
.B(n_32),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_17),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_77),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_28),
.B1(n_16),
.B2(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_71),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_22),
.B1(n_28),
.B2(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_78),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_81),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_22),
.B1(n_20),
.B2(n_30),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_25),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_42),
.B1(n_39),
.B2(n_32),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_70),
.B1(n_56),
.B2(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_49),
.B(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_47),
.B1(n_32),
.B2(n_20),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_85),
.A2(n_53),
.B1(n_44),
.B2(n_51),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_96),
.Y(n_124)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_95),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_14),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_22),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_105),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_32),
.B1(n_19),
.B2(n_36),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_106),
.B1(n_99),
.B2(n_93),
.Y(n_136)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_55),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_103),
.Y(n_150)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_101),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_57),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_21),
.C(n_44),
.Y(n_132)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_21),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_56),
.A2(n_32),
.B1(n_45),
.B2(n_31),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_21),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_121),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_35),
.B1(n_34),
.B2(n_23),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_109),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_47),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_35),
.B1(n_27),
.B2(n_34),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_53),
.A2(n_80),
.B1(n_71),
.B2(n_75),
.Y(n_119)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_0),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_76),
.B(n_21),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_123),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_90),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_126),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_127),
.B(n_144),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_151),
.C(n_142),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_21),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_85),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_91),
.B(n_14),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_96),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_149),
.B1(n_151),
.B2(n_115),
.Y(n_153)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_50),
.B1(n_51),
.B2(n_27),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_102),
.A2(n_50),
.B1(n_27),
.B2(n_34),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_153),
.A2(n_159),
.B1(n_160),
.B2(n_166),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_92),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_163),
.C(n_171),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_155),
.B(n_143),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_158),
.A2(n_0),
.B(n_1),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_119),
.B1(n_102),
.B2(n_118),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_105),
.B1(n_108),
.B2(n_111),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_161),
.B(n_167),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_101),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_168),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_141),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_164),
.A2(n_165),
.B(n_147),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_104),
.B(n_98),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_95),
.B1(n_89),
.B2(n_113),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_133),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_113),
.B1(n_88),
.B2(n_120),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_87),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_87),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_173),
.B(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_54),
.B1(n_52),
.B2(n_23),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_178),
.B(n_182),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_54),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_54),
.B1(n_31),
.B2(n_23),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_31),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_185),
.C(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_129),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_112),
.C(n_1),
.Y(n_185)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_129),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_190),
.B(n_196),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_168),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_191),
.Y(n_222)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_202),
.Y(n_221)
);

AO22x1_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_152),
.B1(n_146),
.B2(n_129),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_176),
.B1(n_179),
.B2(n_2),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_128),
.Y(n_196)
);

AOI22x1_ASAP7_75t_SL g197 ( 
.A1(n_164),
.A2(n_152),
.B1(n_144),
.B2(n_12),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_197),
.A2(n_213),
.B1(n_156),
.B2(n_186),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_158),
.A2(n_128),
.B1(n_130),
.B2(n_125),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_215),
.B1(n_219),
.B2(n_195),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_211),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_210),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_212),
.A2(n_4),
.B(n_6),
.Y(n_235)
);

NAND2x1_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_1),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_1),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g226 ( 
.A(n_214),
.B(n_185),
.Y(n_226)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_163),
.A2(n_125),
.B(n_4),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_2),
.C(n_4),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_181),
.C(n_156),
.Y(n_230)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_164),
.B(n_160),
.C(n_183),
.D(n_153),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_223),
.B(n_218),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_180),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_226),
.C(n_228),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_236),
.B1(n_245),
.B2(n_213),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_227),
.A2(n_233),
.B1(n_200),
.B2(n_194),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_187),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_220),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_232),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_244),
.B(n_247),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_202),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_204),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_243),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_6),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_242),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_214),
.C(n_217),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_195),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_203),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_189),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_192),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_242),
.Y(n_272)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_259),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_221),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_219),
.B1(n_189),
.B2(n_198),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_257),
.B1(n_262),
.B2(n_230),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_267),
.B1(n_271),
.B2(n_227),
.Y(n_277)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_260),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_233),
.A2(n_215),
.B1(n_194),
.B2(n_192),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_203),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_268),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_238),
.A2(n_197),
.B1(n_200),
.B2(n_206),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_224),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_218),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_223),
.C(n_228),
.Y(n_285)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_285),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_252),
.Y(n_274)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_239),
.B1(n_201),
.B2(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_280),
.A2(n_255),
.B1(n_267),
.B2(n_261),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_254),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_283),
.B(n_250),
.Y(n_301)
);

INVx3_ASAP7_75t_SL g284 ( 
.A(n_251),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_211),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_SL g288 ( 
.A(n_253),
.B(n_226),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_249),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_260),
.A2(n_212),
.B(n_235),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_289),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_226),
.C(n_193),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_258),
.C(n_270),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_295),
.Y(n_318)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_258),
.Y(n_295)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_285),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_305),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_299),
.B1(n_303),
.B2(n_304),
.Y(n_307)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_280),
.B(n_249),
.Y(n_302)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_263),
.C(n_209),
.Y(n_305)
);

AOI21x1_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_274),
.B(n_287),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_292),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_316),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_273),
.B1(n_278),
.B2(n_284),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_313),
.C(n_314),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_312),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_275),
.B1(n_282),
.B2(n_286),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_293),
.A2(n_289),
.B(n_281),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_302),
.A2(n_276),
.B1(n_295),
.B2(n_297),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_276),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_292),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_323),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_321),
.A2(n_326),
.B1(n_317),
.B2(n_306),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_310),
.B(n_9),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_10),
.C(n_11),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_308),
.C(n_313),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_315),
.B(n_10),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_318),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_331),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_330),
.B(n_333),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_307),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_327),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_336),
.B(n_337),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_13),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_329),
.B(n_330),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_339),
.A2(n_338),
.B(n_332),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_331),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_342),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_340),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_13),
.Y(n_345)
);


endmodule