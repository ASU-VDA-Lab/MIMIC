module fake_netlist_5_398_n_188 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_188);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_188;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_176;
wire n_140;
wire n_136;
wire n_86;
wire n_146;
wire n_124;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_53;
wire n_160;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_183;
wire n_185;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_181;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_77;
wire n_102;
wire n_64;
wire n_106;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_134;
wire n_187;
wire n_32;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_141;
wire n_97;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVxp67_ASAP7_75t_SL g53 ( 
.A(n_31),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVxp33_ASAP7_75t_SL g55 ( 
.A(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_1),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_47),
.B1(n_39),
.B2(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_6),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

AND3x2_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_44),
.C(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_SL g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_7),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_33),
.B(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_32),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_55),
.B1(n_54),
.B2(n_38),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_33),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_42),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_41),
.B1(n_43),
.B2(n_51),
.Y(n_93)
);

OAI21x1_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_76),
.B(n_63),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_R g95 ( 
.A(n_80),
.B(n_43),
.Y(n_95)
);

AO21x1_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_76),
.B(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_33),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_72),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_88),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_81),
.B(n_78),
.C(n_79),
.Y(n_101)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_71),
.B(n_59),
.Y(n_102)
);

NOR2x1_ASAP7_75t_R g103 ( 
.A(n_86),
.B(n_33),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

AOI21x1_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_75),
.B(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_83),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_89),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_57),
.B1(n_100),
.B2(n_96),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_83),
.Y(n_111)
);

O2A1O1Ixp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_84),
.B(n_73),
.C(n_75),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_80),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_102),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_110),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_95),
.B1(n_86),
.B2(n_33),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_64),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_64),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_112),
.B(n_111),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_111),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

OR2x6_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_116),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_114),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_122),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_114),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_114),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_119),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_120),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_108),
.A3(n_120),
.B1(n_119),
.B2(n_118),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_120),
.B1(n_119),
.B2(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_116),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

NAND2x1_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_116),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_136),
.B1(n_128),
.B2(n_130),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_143),
.B(n_134),
.C(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_128),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_103),
.C(n_90),
.Y(n_147)
);

BUFx4f_ASAP7_75t_SL g148 ( 
.A(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_140),
.A2(n_130),
.B(n_106),
.C(n_74),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_116),
.Y(n_152)
);

AOI211xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_73),
.B(n_132),
.C(n_109),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_127),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

NOR2xp67_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_129),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_127),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_150),
.C(n_129),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_R g164 ( 
.A(n_159),
.B(n_10),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_150),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_127),
.B1(n_116),
.B2(n_83),
.Y(n_166)
);

OAI221xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_87),
.B1(n_116),
.B2(n_11),
.C(n_82),
.Y(n_167)
);

AND2x4_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_116),
.Y(n_168)
);

AOI221x1_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_87),
.B1(n_97),
.B2(n_104),
.C(n_82),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_83),
.B1(n_98),
.B2(n_82),
.Y(n_170)
);

AND3x4_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_14),
.C(n_15),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_162),
.A3(n_87),
.B1(n_154),
.B2(n_27),
.C1(n_28),
.C2(n_29),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_167),
.C(n_163),
.Y(n_173)
);

AOI221xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_97),
.B1(n_110),
.B2(n_23),
.C(n_16),
.Y(n_174)
);

OAI221xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_124),
.B1(n_125),
.B2(n_22),
.C(n_105),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_170),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_125),
.B1(n_124),
.B2(n_83),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_169),
.B1(n_125),
.B2(n_124),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_124),
.B1(n_83),
.B2(n_98),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

NAND2x2_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_98),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_124),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_180),
.A2(n_98),
.B1(n_124),
.B2(n_181),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_185),
.Y(n_187)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_186),
.B1(n_184),
.B2(n_182),
.C(n_179),
.Y(n_188)
);


endmodule