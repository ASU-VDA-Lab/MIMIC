module fake_jpeg_9058_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_0),
.B(n_7),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_3),
.Y(n_12)
);

BUFx2_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_8),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_21),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_20),
.Y(n_36)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_25),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_1),
.C(n_2),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_18),
.C(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_5),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_35),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_9),
.B1(n_16),
.B2(n_14),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_33),
.B1(n_23),
.B2(n_25),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_14),
.B1(n_16),
.B2(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

AOI22x1_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_26),
.B1(n_22),
.B2(n_23),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_36),
.B(n_31),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_46),
.C(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_39),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_43),
.C(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_29),
.Y(n_52)
);

AO21x1_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_52),
.B(n_47),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_54),
.C(n_38),
.Y(n_56)
);


endmodule