module real_jpeg_206_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_215;
wire n_249;
wire n_292;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_197;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_285;
wire n_45;
wire n_160;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_297;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_1),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_86),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_86),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_86),
.Y(n_166)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_3),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_3),
.A2(n_63),
.B1(n_64),
.B2(n_105),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_105),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_105),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_4),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_73),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_73),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_5),
.B(n_151),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_5),
.B(n_64),
.C(n_82),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_5),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_5),
.B(n_81),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_5),
.B(n_29),
.C(n_66),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_186),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_5),
.B(n_33),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_5),
.B(n_99),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_186),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_54),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_6),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_54),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_9),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_71),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_71),
.Y(n_143)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_12),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_150),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_150),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_150),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_14),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_14),
.A2(n_43),
.B1(n_63),
.B2(n_64),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_15),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_126),
.B1(n_300),
.B2(n_301),
.Y(n_18)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_19),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_124),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_109),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_21),
.B(n_109),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.C(n_90),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_22),
.A2(n_23),
.B1(n_75),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_58),
.B2(n_74),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_37),
.B1(n_38),
.B2(n_57),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_26),
.A2(n_38),
.B(n_74),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_26),
.A2(n_57),
.B1(n_59),
.B2(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_34),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_27),
.A2(n_33),
.B1(n_95),
.B2(n_143),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_27),
.A2(n_186),
.B(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_28),
.A2(n_32),
.B1(n_35),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_28),
.A2(n_32),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_28),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_28),
.A2(n_32),
.B1(n_166),
.B2(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_28),
.A2(n_211),
.B(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_28),
.A2(n_32),
.B1(n_211),
.B2(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_29),
.A2(n_30),
.B1(n_66),
.B2(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_29),
.B(n_232),
.Y(n_231)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_32),
.A2(n_165),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_32),
.B(n_180),
.Y(n_213)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_33),
.A2(n_179),
.B(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B(n_51),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_39),
.A2(n_44),
.B1(n_106),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_41),
.B1(n_48),
.B2(n_49),
.Y(n_56)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_41),
.A2(n_106),
.B(n_186),
.C(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_41),
.B(n_186),
.Y(n_187)
);

AOI32xp33_ASAP7_75t_L g198 ( 
.A1(n_41),
.A2(n_46),
.A3(n_48),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_44),
.B(n_53),
.Y(n_108)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_44),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_44),
.A2(n_51),
.B(n_272),
.Y(n_271)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_46),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_45),
.B(n_176),
.Y(n_175)
);

NAND2xp33_ASAP7_75t_SL g200 ( 
.A(n_45),
.B(n_49),
.Y(n_200)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_55),
.A2(n_104),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_59),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_68),
.B1(n_72),
.B2(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_60),
.A2(n_171),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_60),
.A2(n_68),
.B1(n_169),
.B2(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_70),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_61),
.A2(n_99),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_61),
.A2(n_98),
.B1(n_99),
.B2(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_61),
.A2(n_168),
.B(n_170),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_61),
.B(n_172),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_62)
);

AO22x2_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_64),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_64),
.B(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_68),
.A2(n_192),
.B(n_193),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_68),
.A2(n_193),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B(n_89),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_78),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_85),
.B1(n_87),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_87),
.B1(n_88),
.B2(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_79),
.A2(n_87),
.B1(n_159),
.B2(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_79),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_79),
.A2(n_190),
.B(n_252),
.Y(n_270)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_81),
.B(n_147),
.Y(n_252)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_87),
.A2(n_101),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_87),
.A2(n_146),
.B(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_100),
.C(n_102),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_92),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_93),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_99),
.B(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_102),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B(n_107),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_108),
.B(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_123),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_126),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_152),
.B(n_299),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_128),
.B(n_131),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.C(n_137),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_132),
.B(n_135),
.Y(n_297)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_137),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_144),
.C(n_148),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_138),
.A2(n_139),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_140),
.B(n_142),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_141),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_148),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_149),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_294),
.B(n_298),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_263),
.B(n_291),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_205),
.B(n_262),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_181),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_156),
.B(n_181),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_167),
.C(n_173),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_157),
.B(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_161),
.C(n_164),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_167),
.B(n_173),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_195),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_182),
.B(n_196),
.C(n_204),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_188),
.B2(n_194),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_183),
.B(n_189),
.C(n_191),
.Y(n_276)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_188),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_204),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_197),
.B(n_202),
.Y(n_267)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_257),
.B(n_261),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_246),
.B(n_256),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_228),
.B(n_245),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_222),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_222),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_214),
.B1(n_220),
.B2(n_221),
.Y(n_209)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_217),
.C(n_220),
.Y(n_247)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_239),
.B(n_244),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_234),
.B(n_238),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_237),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_236),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_242),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_248),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_253),
.C(n_254),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_260),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_278),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_277),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_277),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_274),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_275),
.C(n_276),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_269),
.C(n_273),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_273),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_290),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_290),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_284),
.C(n_286),
.Y(n_295)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_296),
.Y(n_298)
);


endmodule