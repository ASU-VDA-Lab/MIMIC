module fake_jpeg_22819_n_289 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_0),
.Y(n_48)
);

HAxp5_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_32),
.CON(n_63),
.SN(n_63)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_54),
.Y(n_99)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_18),
.B1(n_23),
.B2(n_20),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_27),
.Y(n_95)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_58),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_63),
.Y(n_96)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_62),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_19),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_68),
.Y(n_117)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_67),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_19),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_19),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_84),
.Y(n_118)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_77),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_18),
.B1(n_23),
.B2(n_36),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_80),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_22),
.B1(n_30),
.B2(n_20),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_18),
.B1(n_36),
.B2(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_38),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_20),
.B1(n_36),
.B2(n_32),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_38),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_33),
.B1(n_35),
.B2(n_34),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_33),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_37),
.B1(n_31),
.B2(n_26),
.Y(n_86)
);

AO22x2_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_87),
.B1(n_75),
.B2(n_72),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_31),
.B1(n_26),
.B2(n_25),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_25),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_63),
.B(n_24),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_107),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_1),
.Y(n_149)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_104),
.Y(n_143)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_106),
.Y(n_151)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_45),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_27),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_21),
.Y(n_124)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_116),
.B(n_1),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_51),
.A2(n_1),
.B(n_2),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_53),
.A3(n_46),
.B1(n_44),
.B2(n_40),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_46),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_131),
.B(n_104),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_65),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_127),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_78),
.B1(n_71),
.B2(n_76),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_65),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_129),
.B(n_135),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_65),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_101),
.C(n_111),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_97),
.C(n_44),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_89),
.Y(n_139)
);

NOR2x1_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_76),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_27),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_90),
.A2(n_114),
.B1(n_95),
.B2(n_96),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_96),
.A2(n_78),
.B1(n_71),
.B2(n_24),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_96),
.A2(n_120),
.B1(n_117),
.B2(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_147),
.A2(n_153),
.B1(n_106),
.B2(n_105),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_98),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_100),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_155),
.A2(n_164),
.B(n_169),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_134),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_170),
.C(n_184),
.Y(n_185)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_168),
.Y(n_186)
);

AO22x1_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_44),
.B1(n_40),
.B2(n_46),
.Y(n_162)
);

AO22x1_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_21),
.B1(n_123),
.B2(n_132),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_178),
.B1(n_141),
.B2(n_136),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_92),
.B(n_107),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_174),
.B1(n_103),
.B2(n_147),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_44),
.B(n_40),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_17),
.A3(n_16),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_175),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_126),
.A2(n_44),
.B(n_40),
.C(n_56),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_138),
.B(n_16),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_40),
.B(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_181),
.A2(n_130),
.B(n_21),
.Y(n_196)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_27),
.B(n_21),
.C(n_5),
.D(n_6),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_122),
.B1(n_152),
.B2(n_136),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_194),
.B1(n_198),
.B2(n_208),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_182),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_192),
.Y(n_227)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_144),
.A3(n_149),
.B1(n_146),
.B2(n_135),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_167),
.Y(n_216)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_200),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_191),
.A2(n_201),
.B1(n_160),
.B2(n_156),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_166),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_196),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_168),
.A2(n_149),
.B1(n_129),
.B2(n_142),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_157),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_161),
.B1(n_181),
.B2(n_162),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_123),
.C(n_56),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_169),
.Y(n_221)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_165),
.C(n_180),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_226),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_198),
.B(n_158),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_224),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_213),
.B(n_219),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_186),
.A2(n_208),
.B1(n_193),
.B2(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_222),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_177),
.B1(n_160),
.B2(n_179),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_206),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_186),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_156),
.B1(n_187),
.B2(n_165),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_235),
.Y(n_245)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_206),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_230),
.A2(n_205),
.B1(n_187),
.B2(n_154),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_237),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_197),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_215),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_164),
.B(n_178),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_210),
.B(n_185),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_211),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_185),
.C(n_155),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_243),
.C(n_211),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_189),
.C(n_201),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_247),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_214),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_251),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_3),
.B(n_4),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_220),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_243),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_212),
.C(n_187),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_255),
.C(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_205),
.Y(n_254)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_254),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_184),
.C(n_207),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_232),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_14),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_233),
.B1(n_234),
.B2(n_242),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_258),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_267),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_255),
.A2(n_240),
.B1(n_132),
.B2(n_199),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_4),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_244),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_265),
.A2(n_250),
.B(n_261),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_260),
.C(n_264),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_271),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_248),
.B1(n_253),
.B2(n_246),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_262),
.A2(n_246),
.B1(n_5),
.B2(n_7),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_273),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_274),
.B(n_258),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_276),
.B(n_269),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_260),
.C(n_266),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_273),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_278),
.B(n_266),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_10),
.C(n_13),
.Y(n_286)
);

NOR4xp25_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_269),
.C(n_272),
.D(n_268),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_279),
.B(n_11),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_286),
.B(n_10),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_285),
.C(n_13),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_13),
.Y(n_289)
);


endmodule