module real_jpeg_7267_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_1),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_1),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_1),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_1),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_1),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_1),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_1),
.B(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_2),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_2),
.B(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_3),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_3),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_3),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_3),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_3),
.B(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_4),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_5),
.B(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_5),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_5),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_5),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_5),
.B(n_240),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_5),
.B(n_281),
.Y(n_280)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_7),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_7),
.B(n_14),
.Y(n_125)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_7),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_8),
.Y(n_184)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_10),
.B(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_10),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_10),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_10),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_10),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_10),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_10),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_10),
.B(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_11),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_12),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_12),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_12),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_12),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_12),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_12),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_12),
.B(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_13),
.Y(n_240)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_14),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_15),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_15),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_15),
.B(n_143),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_192),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_190),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_146),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_19),
.B(n_146),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_100),
.C(n_130),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_20),
.B(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_68),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_21),
.B(n_69),
.C(n_85),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_45),
.C(n_57),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_22),
.B(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_30),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_23),
.B(n_31),
.C(n_44),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_38),
.B2(n_44),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_33),
.B(n_72),
.Y(n_71)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_36),
.Y(n_141)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_36),
.Y(n_213)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_37),
.Y(n_186)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_37),
.Y(n_237)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_37),
.Y(n_268)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_41),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_42),
.Y(n_208)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_43),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_45),
.A2(n_57),
.B1(n_58),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_45),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.C(n_52),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_46),
.A2(n_52),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_46),
.Y(n_201)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_48),
.Y(n_263)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_48),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_50),
.B(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_52),
.Y(n_202)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_55),
.Y(n_243)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_56),
.Y(n_153)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_59),
.A2(n_156),
.B1(n_157),
.B2(n_160),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_59),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_59),
.A2(n_63),
.B1(n_64),
.B2(n_156),
.Y(n_218)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_61),
.Y(n_257)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_62),
.Y(n_248)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_85),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_71),
.B(n_78),
.C(n_83),
.Y(n_189)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_75),
.Y(n_216)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_78),
.A2(n_79),
.B1(n_121),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_79),
.B(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_92),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_88),
.B(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_86),
.B(n_93),
.C(n_97),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_100),
.B(n_130),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_113),
.C(n_118),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_101),
.B(n_113),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_110),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_106),
.C(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_115),
.B(n_262),
.Y(n_261)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_118),
.B(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.C(n_126),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_119),
.A2(n_120),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_121),
.Y(n_300)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_122),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_123),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_145),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_163),
.C(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_138),
.Y(n_164)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_175),
.C(n_176),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_173),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_161),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_157),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_157),
.A2(n_160),
.B1(n_253),
.B2(n_258),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_157),
.B(n_258),
.Y(n_301)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_159),
.Y(n_251)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_159),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_189),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_180)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_185),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_224),
.B(n_326),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_222),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_195),
.B(n_222),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.C(n_219),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_196),
.B(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_198),
.B(n_219),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.C(n_217),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_199),
.B(n_317),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_203),
.A2(n_217),
.B1(n_218),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_203),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.C(n_214),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_204),
.A2(n_205),
.B1(n_214),
.B2(n_215),
.Y(n_305)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_209),
.B(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_321),
.B(n_325),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_307),
.B(n_320),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_293),
.B(n_306),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_269),
.B(n_292),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_259),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_230),
.B(n_259),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_244),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_231),
.B(n_245),
.C(n_252),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_232),
.B(n_239),
.C(n_241),
.Y(n_303)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_249),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_247),
.Y(n_281)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_253),
.Y(n_258)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.C(n_264),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_264),
.B1(n_265),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_286),
.B(n_291),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_279),
.B(n_285),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_278),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_278),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_276),
.Y(n_287)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_295),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_302),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_303),
.C(n_304),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_296),
.Y(n_329)
);

FAx1_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.CI(n_301),
.CON(n_296),
.SN(n_296)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_299),
.C(n_301),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_319),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_319),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_313),
.C(n_316),
.Y(n_322)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_323),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);


endmodule