module fake_ariane_2798_n_2738 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_410, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_350, n_291, n_344, n_381, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_413, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_2738);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_410;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_413;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_2738;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_817;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_524;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_2370;
wire n_2663;
wire n_495;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_2227;
wire n_1512;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_432;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_533;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1790;
wire n_1354;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1443;
wire n_1021;
wire n_491;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_468;
wire n_2703;
wire n_696;
wire n_1442;
wire n_482;
wire n_2620;
wire n_798;
wire n_1833;
wire n_577;
wire n_1691;
wire n_916;
wire n_1386;
wire n_1884;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1972;
wire n_2015;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_436;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2439;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_749;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1832;
wire n_767;
wire n_1392;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_489;
wire n_2294;
wire n_2274;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_471;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1563;
wire n_1020;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_1689;
wire n_970;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2483;
wire n_441;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2662;
wire n_1259;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_2640;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_2476;
wire n_1365;
wire n_553;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2122;
wire n_1611;
wire n_2399;
wire n_1414;
wire n_2067;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2599;
wire n_727;
wire n_699;
wire n_590;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_545;
wire n_2418;
wire n_1614;
wire n_1162;
wire n_536;
wire n_1377;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_501;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2707;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_710;
wire n_534;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_1800;
wire n_982;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_521;
wire n_2140;
wire n_873;
wire n_1748;
wire n_1301;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_2489;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1873;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_1476;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_649;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1759;
wire n_1557;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2525;
wire n_1815;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_473;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2613;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_2234;
wire n_1341;
wire n_1356;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1534;
wire n_453;
wire n_1948;
wire n_1065;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_2121;
wire n_1559;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_1454;
wire n_2592;
wire n_660;
wire n_464;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_519;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_540;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_493;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1758;
wire n_2503;
wire n_1110;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_969;
wire n_2028;
wire n_1663;
wire n_919;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_679;
wire n_663;
wire n_1720;
wire n_2409;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_2676;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_2206;
wire n_997;
wire n_635;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1806;
wire n_1533;
wire n_2372;
wire n_671;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_459;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_2188;
wire n_1777;
wire n_1019;
wire n_1477;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_2587;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_537;
wire n_1063;
wire n_2205;
wire n_2183;
wire n_991;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_1474;
wire n_2081;
wire n_937;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1722;
wire n_1001;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1644;
wire n_1002;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_431;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_1820;
wire n_2590;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_357),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_374),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_65),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_110),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_227),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_342),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_248),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_90),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_230),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_395),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_396),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_180),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_225),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_198),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_33),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_86),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_349),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_142),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_30),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_159),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_55),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_369),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_11),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_2),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_361),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_185),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_162),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_372),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_400),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_18),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_87),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_389),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_238),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_88),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_50),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_316),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_335),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_336),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_363),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_258),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_168),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_7),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_385),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_267),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_355),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_232),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_260),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_74),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_185),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_184),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_77),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_92),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_154),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_364),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_366),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_82),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_125),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_8),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_314),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_262),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_320),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_85),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_391),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_334),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_237),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_3),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_9),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_346),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_261),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_180),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_207),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_270),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_90),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_178),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_298),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_318),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_265),
.Y(n_491)
);

BUFx10_ASAP7_75t_L g492 ( 
.A(n_234),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_371),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_222),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_169),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_139),
.Y(n_496)
);

BUFx5_ASAP7_75t_L g497 ( 
.A(n_337),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_325),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_379),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_327),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_300),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_98),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_301),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_362),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_6),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_87),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_44),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_308),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_360),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_40),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_338),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_52),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_311),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_409),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_129),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_199),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_204),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_55),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_178),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_275),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_81),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_351),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_304),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_235),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_42),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_227),
.Y(n_526)
);

INVxp33_ASAP7_75t_SL g527 ( 
.A(n_352),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_333),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_268),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_297),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_220),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_356),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_162),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_413),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_122),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_115),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_82),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_30),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_197),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_393),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_402),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_75),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_330),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_136),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_399),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_322),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_152),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_343),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_156),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_219),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_112),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_121),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_394),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_386),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_408),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_79),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_313),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_60),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_404),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_291),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_67),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_35),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_290),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_49),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_228),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_365),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_75),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_359),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_299),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_388),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_256),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_410),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_384),
.Y(n_573)
);

INVxp67_ASAP7_75t_SL g574 ( 
.A(n_285),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_117),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_25),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_263),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_319),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_29),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_414),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_97),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_387),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_114),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_32),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_97),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_331),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_122),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_222),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_307),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_340),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_172),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_71),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_347),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_80),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_144),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_151),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_302),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_169),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_91),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_383),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_57),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_309),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_188),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_28),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_203),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_102),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_345),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_72),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_6),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_57),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_375),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_276),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_108),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_191),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_312),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_306),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_310),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_25),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_354),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_407),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_36),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_78),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_411),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_123),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_212),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_174),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_324),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_139),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_71),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_228),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_77),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_220),
.Y(n_632)
);

BUFx8_ASAP7_75t_SL g633 ( 
.A(n_116),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_370),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_63),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_323),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_145),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_317),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_21),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_194),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_99),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_81),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_332),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_339),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_54),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_28),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_133),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_20),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_159),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_134),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_272),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_69),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_168),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_183),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_121),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_63),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_5),
.Y(n_657)
);

BUFx2_ASAP7_75t_SL g658 ( 
.A(n_54),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_303),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_367),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_45),
.Y(n_661)
);

BUFx5_ASAP7_75t_L g662 ( 
.A(n_0),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_406),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_212),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_412),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_109),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_189),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_202),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_378),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_242),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_358),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_305),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_405),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_183),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_236),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_187),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_116),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_163),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_161),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_254),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_321),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_150),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_245),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_164),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_123),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_170),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_197),
.Y(n_687)
);

CKINVDCx14_ASAP7_75t_R g688 ( 
.A(n_22),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_353),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_133),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_392),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_377),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_124),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_64),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_233),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_214),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_127),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_373),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_218),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_160),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_368),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_136),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_47),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_202),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_341),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_195),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_380),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_119),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_328),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_241),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_72),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_287),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_35),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_160),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_315),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_43),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_229),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_88),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_381),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_166),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_350),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_132),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_284),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_170),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_0),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_191),
.Y(n_726)
);

BUFx10_ASAP7_75t_L g727 ( 
.A(n_257),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_401),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_79),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_292),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_26),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_390),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_102),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_348),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_100),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_329),
.Y(n_736)
);

CKINVDCx14_ASAP7_75t_R g737 ( 
.A(n_195),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_403),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_294),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_60),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_397),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_83),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_78),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_12),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_53),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_200),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_51),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_41),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_376),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_134),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_398),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_96),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_52),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_58),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_163),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_85),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_27),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_145),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_19),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_326),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_95),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_382),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_278),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_203),
.Y(n_764)
);

BUFx10_ASAP7_75t_L g765 ( 
.A(n_110),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_73),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_155),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_187),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_206),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_344),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_199),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_217),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_120),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_218),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_34),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_103),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_221),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_219),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_662),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_629),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_552),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_427),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_427),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_434),
.Y(n_784)
);

INVxp33_ASAP7_75t_SL g785 ( 
.A(n_725),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_688),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_419),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_434),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_750),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_662),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_440),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_642),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_537),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_537),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_606),
.Y(n_795)
);

INVxp33_ASAP7_75t_SL g796 ( 
.A(n_728),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_653),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_737),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_662),
.Y(n_799)
);

CKINVDCx14_ASAP7_75t_R g800 ( 
.A(n_482),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_606),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_704),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_463),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_704),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_758),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_653),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_758),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_662),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_658),
.Y(n_809)
);

INVxp33_ASAP7_75t_SL g810 ( 
.A(n_417),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_654),
.B(n_1),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_662),
.Y(n_812)
);

INVxp67_ASAP7_75t_SL g813 ( 
.A(n_653),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_662),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_662),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_633),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_462),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_762),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_417),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_482),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_662),
.Y(n_821)
);

INVxp33_ASAP7_75t_SL g822 ( 
.A(n_418),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_422),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_426),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_433),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_438),
.Y(n_826)
);

INVxp33_ASAP7_75t_SL g827 ( 
.A(n_418),
.Y(n_827)
);

NOR2xp67_ASAP7_75t_L g828 ( 
.A(n_462),
.B(n_1),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_449),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_609),
.B(n_2),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_546),
.Y(n_831)
);

INVxp67_ASAP7_75t_SL g832 ( 
.A(n_653),
.Y(n_832)
);

BUFx10_ASAP7_75t_L g833 ( 
.A(n_653),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_482),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_492),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_455),
.Y(n_836)
);

INVxp33_ASAP7_75t_SL g837 ( 
.A(n_428),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_456),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_470),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_702),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_702),
.Y(n_841)
);

INVxp67_ASAP7_75t_SL g842 ( 
.A(n_702),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_546),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_702),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_702),
.Y(n_845)
);

INVxp33_ASAP7_75t_L g846 ( 
.A(n_472),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_714),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_714),
.Y(n_848)
);

INVxp67_ASAP7_75t_SL g849 ( 
.A(n_714),
.Y(n_849)
);

INVxp33_ASAP7_75t_SL g850 ( 
.A(n_428),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_714),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_714),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_488),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_488),
.Y(n_854)
);

INVxp33_ASAP7_75t_SL g855 ( 
.A(n_429),
.Y(n_855)
);

INVxp33_ASAP7_75t_L g856 ( 
.A(n_494),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_439),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_517),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_594),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_644),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_521),
.Y(n_861)
);

INVxp33_ASAP7_75t_L g862 ( 
.A(n_531),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_533),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_429),
.Y(n_864)
);

INVx4_ASAP7_75t_R g865 ( 
.A(n_644),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_535),
.Y(n_866)
);

NOR2xp67_ASAP7_75t_L g867 ( 
.A(n_609),
.B(n_3),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_639),
.B(n_4),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_542),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_556),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_558),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_421),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_430),
.Y(n_873)
);

CKINVDCx14_ASAP7_75t_R g874 ( 
.A(n_492),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_562),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_423),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_639),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_564),
.Y(n_878)
);

NOR2xp67_ASAP7_75t_L g879 ( 
.A(n_743),
.B(n_4),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_492),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_581),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_641),
.Y(n_882)
);

INVxp67_ASAP7_75t_SL g883 ( 
.A(n_594),
.Y(n_883)
);

INVxp33_ASAP7_75t_L g884 ( 
.A(n_575),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_636),
.Y(n_885)
);

INVxp67_ASAP7_75t_SL g886 ( 
.A(n_637),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_584),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_585),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_636),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_592),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_599),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_636),
.Y(n_892)
);

INVxp33_ASAP7_75t_L g893 ( 
.A(n_603),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_727),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_424),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_645),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_604),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_610),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_678),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_439),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_727),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_614),
.Y(n_902)
);

INVxp67_ASAP7_75t_SL g903 ( 
.A(n_637),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_624),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_625),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_727),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_415),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_646),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_647),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_650),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_656),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_661),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_516),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_415),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_666),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_425),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_682),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_431),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_684),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_693),
.Y(n_920)
);

INVxp33_ASAP7_75t_SL g921 ( 
.A(n_430),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_743),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_446),
.Y(n_923)
);

INVxp67_ASAP7_75t_SL g924 ( 
.A(n_640),
.Y(n_924)
);

INVxp33_ASAP7_75t_SL g925 ( 
.A(n_432),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_471),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_699),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_451),
.Y(n_928)
);

INVxp33_ASAP7_75t_L g929 ( 
.A(n_703),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_708),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_432),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_471),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_711),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_718),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_726),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_640),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_740),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_420),
.Y(n_938)
);

INVxp33_ASAP7_75t_L g939 ( 
.A(n_744),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_747),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_452),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_748),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_753),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_754),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_468),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_764),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_767),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_690),
.B(n_5),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_778),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_435),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_690),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_420),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_436),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_773),
.Y(n_954)
);

INVxp33_ASAP7_75t_L g955 ( 
.A(n_459),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_436),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_439),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_773),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_435),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_474),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_471),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_676),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_676),
.Y(n_963)
);

NOR2xp67_ASAP7_75t_L g964 ( 
.A(n_437),
.B(n_441),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_676),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_685),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_685),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_437),
.B(n_7),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_685),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_735),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_735),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_735),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_765),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_479),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_439),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_765),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_765),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_483),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_489),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_498),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_508),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_513),
.Y(n_982)
);

INVxp33_ASAP7_75t_L g983 ( 
.A(n_459),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_501),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_520),
.Y(n_985)
);

CKINVDCx16_ASAP7_75t_R g986 ( 
.A(n_416),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_530),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_441),
.Y(n_988)
);

INVxp67_ASAP7_75t_SL g989 ( 
.A(n_501),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_444),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_532),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_540),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_444),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_541),
.Y(n_994)
);

INVxp67_ASAP7_75t_SL g995 ( 
.A(n_589),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_548),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_557),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_570),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_580),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_586),
.Y(n_1000)
);

INVxp33_ASAP7_75t_SL g1001 ( 
.A(n_445),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_447),
.Y(n_1002)
);

INVxp33_ASAP7_75t_SL g1003 ( 
.A(n_445),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_590),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_442),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_442),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_615),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_620),
.Y(n_1008)
);

BUFx2_ASAP7_75t_SL g1009 ( 
.A(n_453),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_623),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_448),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_443),
.Y(n_1012)
);

INVxp67_ASAP7_75t_SL g1013 ( 
.A(n_589),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_638),
.Y(n_1014)
);

CKINVDCx16_ASAP7_75t_R g1015 ( 
.A(n_461),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_659),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_669),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_681),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_689),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_717),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_721),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_723),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_448),
.Y(n_1023)
);

INVxp67_ASAP7_75t_SL g1024 ( 
.A(n_627),
.Y(n_1024)
);

INVxp33_ASAP7_75t_L g1025 ( 
.A(n_627),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_491),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_734),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_741),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_464),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_559),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_464),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_643),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_465),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_643),
.B(n_8),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_663),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_465),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_663),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_466),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_466),
.Y(n_1039)
);

INVxp33_ASAP7_75t_L g1040 ( 
.A(n_760),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_760),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_698),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_497),
.Y(n_1043)
);

INVxp67_ASAP7_75t_SL g1044 ( 
.A(n_698),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_467),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_497),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_439),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_467),
.Y(n_1048)
);

INVxp67_ASAP7_75t_SL g1049 ( 
.A(n_527),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_476),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_612),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_476),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_497),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_443),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_619),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_715),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_480),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_480),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_497),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_481),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_481),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_484),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_739),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_484),
.Y(n_1064)
);

INVxp67_ASAP7_75t_SL g1065 ( 
.A(n_617),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_503),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_485),
.Y(n_1067)
);

INVx5_ASAP7_75t_L g1068 ( 
.A(n_857),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_SL g1069 ( 
.A(n_913),
.B(n_550),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_813),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_1044),
.B(n_500),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_857),
.Y(n_1072)
);

BUFx12f_ASAP7_75t_L g1073 ( 
.A(n_816),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_857),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_797),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_800),
.B(n_485),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_857),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_831),
.B(n_712),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_831),
.B(n_574),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_843),
.B(n_598),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_1009),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_832),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_874),
.B(n_955),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_797),
.Y(n_1084)
);

BUFx12f_ASAP7_75t_L g1085 ( 
.A(n_816),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_983),
.B(n_504),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_842),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_803),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_857),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_819),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_849),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_779),
.A2(n_812),
.B(n_790),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_823),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_796),
.B(n_450),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_797),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_806),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_900),
.Y(n_1097)
);

OAI22x1_ASAP7_75t_SL g1098 ( 
.A1(n_787),
.A2(n_495),
.B1(n_496),
.B2(n_487),
.Y(n_1098)
);

OAI22x1_ASAP7_75t_L g1099 ( 
.A1(n_818),
.A2(n_755),
.B1(n_757),
.B2(n_652),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_819),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_806),
.Y(n_1101)
);

NOR2x1_ASAP7_75t_L g1102 ( 
.A(n_1066),
.B(n_617),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_900),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_824),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_806),
.Y(n_1105)
);

OA22x2_ASAP7_75t_SL g1106 ( 
.A1(n_1049),
.A2(n_495),
.B1(n_496),
.B2(n_487),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_796),
.A2(n_776),
.B1(n_769),
.B2(n_696),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_833),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1047),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_900),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_825),
.Y(n_1111)
);

AOI22x1_ASAP7_75t_SL g1112 ( 
.A1(n_1002),
.A2(n_696),
.B1(n_697),
.B2(n_694),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_826),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1047),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1025),
.B(n_509),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1009),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_907),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_907),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1029),
.B(n_1036),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_864),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_818),
.A2(n_505),
.B1(n_506),
.B2(n_502),
.Y(n_1121)
);

INVx5_ASAP7_75t_L g1122 ( 
.A(n_900),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_840),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_840),
.Y(n_1124)
);

INVx5_ASAP7_75t_L g1125 ( 
.A(n_900),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_841),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_833),
.Y(n_1127)
);

OA21x2_ASAP7_75t_L g1128 ( 
.A1(n_814),
.A2(n_454),
.B(n_450),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_833),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_829),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1040),
.B(n_511),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_841),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_957),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_844),
.Y(n_1134)
);

INVx5_ASAP7_75t_L g1135 ( 
.A(n_957),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_820),
.B(n_454),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_957),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_914),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_844),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_845),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_785),
.A2(n_510),
.B1(n_512),
.B2(n_507),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_845),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_836),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_786),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_957),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_914),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_938),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_1032),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_957),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_838),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_847),
.Y(n_1151)
);

INVx5_ASAP7_75t_L g1152 ( 
.A(n_975),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_846),
.B(n_694),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_839),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_975),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_864),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1038),
.B(n_457),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_858),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_938),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1066),
.B(n_514),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_975),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_847),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_975),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1032),
.Y(n_1164)
);

BUFx8_ASAP7_75t_SL g1165 ( 
.A(n_787),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_784),
.B(n_522),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_931),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_861),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_975),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_952),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_843),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_848),
.Y(n_1172)
);

BUFx12f_ASAP7_75t_L g1173 ( 
.A(n_786),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1037),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_876),
.B(n_617),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1037),
.Y(n_1176)
);

AND2x2_ASAP7_75t_SL g1177 ( 
.A(n_948),
.B(n_617),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_848),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_851),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_851),
.Y(n_1180)
);

AND2x2_ASAP7_75t_R g1181 ( 
.A(n_1002),
.B(n_697),
.Y(n_1181)
);

OAI22x1_ASAP7_75t_SL g1182 ( 
.A1(n_791),
.A2(n_706),
.B1(n_713),
.B2(n_700),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_860),
.B(n_523),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_863),
.Y(n_1184)
);

INVx5_ASAP7_75t_L g1185 ( 
.A(n_1035),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_798),
.Y(n_1186)
);

BUFx12f_ASAP7_75t_L g1187 ( 
.A(n_798),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_866),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_876),
.B(n_617),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_856),
.B(n_700),
.Y(n_1190)
);

AND2x6_ASAP7_75t_L g1191 ( 
.A(n_1043),
.B(n_763),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_869),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1039),
.B(n_1048),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_860),
.B(n_984),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_862),
.B(n_884),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_870),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_852),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_895),
.B(n_916),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_989),
.B(n_524),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_931),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_952),
.Y(n_1201)
);

OAI22x1_ASAP7_75t_R g1202 ( 
.A1(n_791),
.A2(n_777),
.B1(n_713),
.B2(n_716),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_852),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_895),
.B(n_763),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_871),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_875),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_953),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1035),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_820),
.B(n_457),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_878),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_785),
.A2(n_777),
.B1(n_716),
.B2(n_720),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_893),
.B(n_706),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_779),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_953),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_887),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_790),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_881),
.Y(n_1217)
);

INVx4_ASAP7_75t_L g1218 ( 
.A(n_1035),
.Y(n_1218)
);

INVx6_ASAP7_75t_L g1219 ( 
.A(n_916),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_888),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_995),
.B(n_528),
.Y(n_1221)
);

BUFx12f_ASAP7_75t_L g1222 ( 
.A(n_834),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_956),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_890),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_872),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_821),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_891),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_956),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_821),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1013),
.B(n_529),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_897),
.Y(n_1231)
);

BUFx8_ASAP7_75t_L g1232 ( 
.A(n_1031),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_815),
.Y(n_1233)
);

INVx6_ASAP7_75t_L g1234 ( 
.A(n_945),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_834),
.B(n_458),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_872),
.Y(n_1236)
);

BUFx12f_ASAP7_75t_L g1237 ( 
.A(n_835),
.Y(n_1237)
);

BUFx12f_ASAP7_75t_L g1238 ( 
.A(n_835),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1046),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_799),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1046),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_918),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1050),
.B(n_458),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1024),
.B(n_534),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1005),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_898),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1031),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_945),
.B(n_763),
.Y(n_1248)
);

BUFx8_ASAP7_75t_L g1249 ( 
.A(n_1045),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1005),
.Y(n_1250)
);

AND2x6_ASAP7_75t_L g1251 ( 
.A(n_1083),
.B(n_763),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1071),
.B(n_880),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1093),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1239),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1104),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1198),
.B(n_961),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1239),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1239),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1111),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1113),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1130),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1198),
.B(n_962),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1239),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_1195),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1092),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1092),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1143),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1241),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1153),
.B(n_1045),
.Y(n_1269)
);

NAND2xp33_ASAP7_75t_L g1270 ( 
.A(n_1223),
.B(n_1117),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1150),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1166),
.B(n_1006),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1177),
.B(n_859),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1213),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1177),
.B(n_883),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1213),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1216),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1154),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1158),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_SL g1280 ( 
.A(n_1069),
.B(n_810),
.Y(n_1280)
);

INVx6_ASAP7_75t_L g1281 ( 
.A(n_1219),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1168),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1184),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1188),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1127),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1073),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1071),
.B(n_885),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1198),
.B(n_886),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1071),
.B(n_885),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1199),
.B(n_1006),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1218),
.B(n_889),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1218),
.B(n_889),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1192),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1196),
.Y(n_1294)
);

INVx6_ASAP7_75t_L g1295 ( 
.A(n_1219),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1205),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1240),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1206),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1171),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1218),
.B(n_892),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1241),
.Y(n_1301)
);

OR2x6_ASAP7_75t_L g1302 ( 
.A(n_1073),
.B(n_811),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1210),
.Y(n_1303)
);

OAI22x1_ASAP7_75t_SL g1304 ( 
.A1(n_1217),
.A2(n_882),
.B1(n_896),
.B2(n_881),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1215),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1220),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1222),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1127),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1224),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1227),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1190),
.B(n_903),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1241),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1240),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1127),
.B(n_894),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1233),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1171),
.B(n_1079),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1078),
.B(n_894),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1226),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1231),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1246),
.Y(n_1320)
);

AND2x6_ASAP7_75t_L g1321 ( 
.A(n_1175),
.B(n_763),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1070),
.Y(n_1322)
);

AND2x6_ASAP7_75t_L g1323 ( 
.A(n_1175),
.B(n_1034),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1222),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1233),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1212),
.B(n_924),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1078),
.B(n_960),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1217),
.A2(n_896),
.B1(n_899),
.B2(n_882),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1082),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1087),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1226),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1091),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1088),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1208),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1208),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1208),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1225),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1226),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1225),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1225),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1236),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1079),
.B(n_1012),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1146),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1117),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1229),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1078),
.B(n_880),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1080),
.B(n_960),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1079),
.B(n_963),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1236),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1229),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1236),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1242),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1118),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1242),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1133),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1229),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1242),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1223),
.B(n_1054),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1109),
.A2(n_808),
.B(n_1053),
.Y(n_1359)
);

OR2x6_ASAP7_75t_L g1360 ( 
.A(n_1085),
.B(n_811),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_SL g1361 ( 
.A(n_1237),
.B(n_810),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1133),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1229),
.Y(n_1363)
);

CKINVDCx8_ASAP7_75t_R g1364 ( 
.A(n_1118),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1197),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1133),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1080),
.B(n_1000),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1080),
.B(n_965),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1148),
.Y(n_1369)
);

BUFx8_ASAP7_75t_L g1370 ( 
.A(n_1085),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1109),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1148),
.Y(n_1372)
);

CKINVDCx16_ASAP7_75t_R g1373 ( 
.A(n_1237),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1148),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1197),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1100),
.B(n_986),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1164),
.Y(n_1377)
);

CKINVDCx8_ASAP7_75t_R g1378 ( 
.A(n_1138),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1119),
.B(n_906),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1114),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1114),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1090),
.B(n_972),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1075),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1197),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1194),
.B(n_966),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1164),
.Y(n_1386)
);

INVx6_ASAP7_75t_L g1387 ( 
.A(n_1219),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1075),
.Y(n_1388)
);

AND2x6_ASAP7_75t_L g1389 ( 
.A(n_1175),
.B(n_918),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1076),
.B(n_1000),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1084),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1164),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1084),
.Y(n_1393)
);

AND2x6_ASAP7_75t_L g1394 ( 
.A(n_1189),
.B(n_923),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1174),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1119),
.B(n_967),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1174),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1197),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1193),
.B(n_906),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1174),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1176),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1176),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_SL g1403 ( 
.A1(n_1094),
.A2(n_899),
.B1(n_1030),
.B2(n_1026),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1095),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1138),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1203),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1176),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1193),
.B(n_969),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1274),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1333),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1322),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1379),
.B(n_1159),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1329),
.Y(n_1413)
);

INVx6_ASAP7_75t_L g1414 ( 
.A(n_1281),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1399),
.B(n_1094),
.C(n_1159),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1343),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1330),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1355),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1302),
.B(n_1238),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1252),
.B(n_1136),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1290),
.B(n_1157),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1269),
.B(n_1147),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1332),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1287),
.B(n_1136),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1327),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1270),
.B(n_1214),
.C(n_1207),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1274),
.Y(n_1427)
);

INVx5_ASAP7_75t_L g1428 ( 
.A(n_1321),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1253),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_1316),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1285),
.B(n_1214),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1290),
.B(n_1273),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1355),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1276),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1285),
.B(n_1207),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1289),
.B(n_1235),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1255),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1259),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1276),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1273),
.A2(n_1275),
.B1(n_1323),
.B2(n_1311),
.Y(n_1440)
);

INVx4_ASAP7_75t_L g1441 ( 
.A(n_1281),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1285),
.B(n_1228),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1270),
.B(n_1054),
.C(n_1012),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1286),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1275),
.B(n_1157),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1272),
.B(n_1243),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1254),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1277),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1260),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1342),
.B(n_1235),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1323),
.A2(n_1128),
.B1(n_948),
.B2(n_928),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1261),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1286),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1281),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1267),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1271),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1342),
.B(n_1209),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1278),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1272),
.B(n_1243),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1355),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1362),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1279),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1317),
.B(n_1209),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1282),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1277),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1308),
.B(n_1245),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1376),
.B(n_1015),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1344),
.Y(n_1468)
);

AND3x2_ASAP7_75t_L g1469 ( 
.A(n_1361),
.B(n_1201),
.C(n_1170),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1283),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1280),
.A2(n_1141),
.B1(n_1121),
.B2(n_1250),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1362),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1284),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1307),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1307),
.Y(n_1475)
);

AOI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1265),
.A2(n_1183),
.B(n_1128),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1362),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1327),
.B(n_1086),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1293),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1353),
.B(n_1120),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1294),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1296),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1254),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1323),
.A2(n_1116),
.B1(n_1081),
.B2(n_1167),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1308),
.B(n_1081),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1405),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1323),
.A2(n_1128),
.B1(n_928),
.B2(n_941),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1298),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1382),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1366),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1303),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1305),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1347),
.B(n_1367),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1323),
.A2(n_1396),
.B1(n_1408),
.B2(n_1316),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1308),
.B(n_1314),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1306),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1366),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1347),
.B(n_1115),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1309),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1264),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_L g1501 ( 
.A(n_1265),
.B(n_1116),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1310),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1324),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1396),
.B(n_1108),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1367),
.B(n_1131),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1366),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_SL g1507 ( 
.A1(n_1403),
.A2(n_1030),
.B1(n_1051),
.B2(n_1026),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1346),
.B(n_1358),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1295),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1319),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1390),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1258),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1320),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1358),
.B(n_1221),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1258),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_SL g1516 ( 
.A(n_1302),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1396),
.B(n_1108),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1408),
.B(n_1230),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1408),
.B(n_1244),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1324),
.Y(n_1520)
);

OAI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1364),
.A2(n_1238),
.B1(n_1107),
.B2(n_827),
.Y(n_1521)
);

NAND2xp33_ASAP7_75t_R g1522 ( 
.A(n_1302),
.B(n_892),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1316),
.B(n_1291),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1390),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1311),
.B(n_901),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1297),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1292),
.B(n_1160),
.Y(n_1527)
);

NAND2xp33_ASAP7_75t_L g1528 ( 
.A(n_1266),
.B(n_1200),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1258),
.Y(n_1529)
);

NAND2xp33_ASAP7_75t_L g1530 ( 
.A(n_1266),
.B(n_1247),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1313),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1326),
.B(n_1156),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1300),
.B(n_1234),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1370),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1313),
.Y(n_1535)
);

INVxp33_ASAP7_75t_L g1536 ( 
.A(n_1328),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1373),
.B(n_1211),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1383),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1326),
.B(n_901),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1295),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1383),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1268),
.B(n_1129),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_R g1543 ( 
.A(n_1364),
.B(n_1144),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1288),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1268),
.B(n_1129),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1315),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1348),
.B(n_1234),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1315),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1388),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1325),
.A2(n_941),
.B1(n_974),
.B2(n_923),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1388),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1325),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1268),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1359),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1288),
.Y(n_1555)
);

INVxp67_ASAP7_75t_SL g1556 ( 
.A(n_1254),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1254),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1391),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1391),
.Y(n_1559)
);

INVx8_ASAP7_75t_L g1560 ( 
.A(n_1360),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1348),
.B(n_1234),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1560),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1432),
.B(n_1378),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1409),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1494),
.B(n_1378),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1416),
.Y(n_1566)
);

BUFx4f_ASAP7_75t_L g1567 ( 
.A(n_1560),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1447),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1409),
.Y(n_1569)
);

OAI21xp33_ASAP7_75t_L g1570 ( 
.A1(n_1421),
.A2(n_827),
.B(n_822),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1446),
.B(n_1249),
.C(n_1232),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1459),
.B(n_1385),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1445),
.B(n_1368),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1450),
.B(n_1257),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1422),
.B(n_1368),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1560),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_L g1577 ( 
.A(n_1420),
.B(n_1249),
.C(n_1232),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1532),
.B(n_1368),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1427),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1447),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1420),
.B(n_1385),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1411),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1424),
.B(n_1436),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1440),
.A2(n_1099),
.B1(n_1394),
.B2(n_1389),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1424),
.B(n_1385),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1450),
.B(n_1257),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1413),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1417),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1440),
.A2(n_1394),
.B1(n_1389),
.B2(n_1380),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1489),
.B(n_1348),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1543),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1410),
.Y(n_1592)
);

AND2x2_ASAP7_75t_SL g1593 ( 
.A(n_1451),
.B(n_1487),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1427),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1423),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1468),
.B(n_1256),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1436),
.B(n_1256),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1486),
.B(n_1256),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1434),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1544),
.B(n_1262),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1429),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1463),
.B(n_1262),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1430),
.B(n_1299),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1434),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1447),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1463),
.B(n_1262),
.Y(n_1606)
);

NAND2xp33_ASAP7_75t_L g1607 ( 
.A(n_1543),
.B(n_1334),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1437),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1447),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1555),
.B(n_1360),
.Y(n_1610)
);

AOI22x1_ASAP7_75t_L g1611 ( 
.A1(n_1418),
.A2(n_1335),
.B1(n_1336),
.B2(n_1337),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1518),
.B(n_1389),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1483),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1525),
.B(n_1360),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1539),
.B(n_873),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1415),
.B(n_1249),
.C(n_1232),
.Y(n_1616)
);

AO22x2_ASAP7_75t_L g1617 ( 
.A1(n_1507),
.A2(n_1112),
.B1(n_1202),
.B2(n_1304),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1519),
.B(n_1389),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1438),
.Y(n_1619)
);

INVx4_ASAP7_75t_L g1620 ( 
.A(n_1428),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1449),
.Y(n_1621)
);

NOR2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1474),
.B(n_1144),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1483),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1508),
.B(n_1389),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1454),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1428),
.Y(n_1626)
);

NAND2x1p5_ASAP7_75t_L g1627 ( 
.A(n_1428),
.B(n_1299),
.Y(n_1627)
);

INVx4_ASAP7_75t_L g1628 ( 
.A(n_1428),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1454),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1475),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1528),
.B(n_990),
.C(n_988),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1419),
.B(n_1394),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1452),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1457),
.B(n_1295),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1419),
.B(n_1173),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1480),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1540),
.Y(n_1637)
);

INVx4_ASAP7_75t_L g1638 ( 
.A(n_1414),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1455),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1540),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1456),
.Y(n_1641)
);

BUFx10_ASAP7_75t_L g1642 ( 
.A(n_1503),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1508),
.B(n_1394),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1439),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1483),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1439),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1514),
.B(n_1394),
.Y(n_1647)
);

INVx4_ASAP7_75t_L g1648 ( 
.A(n_1414),
.Y(n_1648)
);

INVx4_ASAP7_75t_L g1649 ( 
.A(n_1414),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1467),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1448),
.Y(n_1651)
);

NAND2x1p5_ASAP7_75t_L g1652 ( 
.A(n_1441),
.B(n_1312),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1523),
.B(n_1514),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1419),
.B(n_1339),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1441),
.B(n_1312),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1458),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1493),
.B(n_1340),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1483),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1425),
.B(n_1511),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1448),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1500),
.B(n_950),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1524),
.B(n_959),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1469),
.B(n_1341),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1462),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1528),
.B(n_1058),
.C(n_1033),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1547),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1464),
.Y(n_1667)
);

INVx4_ASAP7_75t_L g1668 ( 
.A(n_1509),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1520),
.B(n_993),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1537),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1478),
.B(n_1011),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1465),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1470),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1498),
.B(n_1387),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1473),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1479),
.Y(n_1676)
);

BUFx4f_ASAP7_75t_L g1677 ( 
.A(n_1481),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1482),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1471),
.B(n_1064),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1444),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1505),
.B(n_1387),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1488),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1491),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1523),
.B(n_1257),
.Y(n_1684)
);

INVxp67_ASAP7_75t_SL g1685 ( 
.A(n_1554),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1492),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1583),
.B(n_1484),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1562),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1583),
.B(n_1547),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1568),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1593),
.A2(n_1536),
.B1(n_1055),
.B2(n_1056),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1564),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1653),
.A2(n_1495),
.B(n_1527),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_SL g1694 ( 
.A(n_1591),
.B(n_1534),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1597),
.A2(n_1521),
.B1(n_1530),
.B2(n_1561),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1592),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1563),
.B(n_1426),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1564),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1563),
.B(n_1051),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1569),
.Y(n_1700)
);

O2A1O1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1570),
.A2(n_1530),
.B(n_822),
.C(n_850),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1573),
.B(n_1561),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1573),
.B(n_1572),
.Y(n_1703)
);

AND2x6_ASAP7_75t_L g1704 ( 
.A(n_1632),
.B(n_1418),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1597),
.B(n_1606),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1606),
.A2(n_1435),
.B1(n_1431),
.B2(n_1527),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1562),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1569),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1579),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_1685),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1581),
.B(n_1496),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1636),
.B(n_1055),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1579),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1593),
.A2(n_1679),
.B1(n_1536),
.B2(n_1590),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1594),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1620),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1585),
.B(n_1499),
.Y(n_1717)
);

O2A1O1Ixp5_ASAP7_75t_L g1718 ( 
.A1(n_1653),
.A2(n_1435),
.B(n_1431),
.C(n_1485),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1602),
.B(n_1502),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1594),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1677),
.B(n_1443),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1671),
.B(n_1510),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1578),
.B(n_1550),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1599),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1576),
.B(n_1509),
.Y(n_1725)
);

OAI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1650),
.A2(n_1106),
.B1(n_809),
.B2(n_781),
.C(n_1412),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1677),
.B(n_1412),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1596),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1666),
.B(n_1575),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1598),
.Y(n_1730)
);

INVx3_ASAP7_75t_L g1731 ( 
.A(n_1620),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1666),
.B(n_1513),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1603),
.B(n_1485),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1615),
.B(n_1504),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1565),
.B(n_1056),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1634),
.B(n_1504),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1634),
.B(n_1550),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1566),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1669),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1603),
.B(n_1614),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1603),
.B(n_1517),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1657),
.B(n_1451),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1626),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1624),
.A2(n_1487),
.B(n_1495),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1599),
.Y(n_1745)
);

AND2x6_ASAP7_75t_L g1746 ( 
.A(n_1632),
.B(n_1433),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1582),
.A2(n_1460),
.B1(n_1461),
.B2(n_1433),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1600),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1674),
.B(n_1517),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1657),
.B(n_1546),
.Y(n_1750)
);

AND2x2_ASAP7_75t_SL g1751 ( 
.A(n_1589),
.B(n_1501),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1674),
.B(n_1063),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1617),
.A2(n_1063),
.B1(n_926),
.B2(n_932),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1604),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1604),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1644),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1644),
.Y(n_1757)
);

AND2x6_ASAP7_75t_SL g1758 ( 
.A(n_1635),
.B(n_830),
.Y(n_1758)
);

BUFx12f_ASAP7_75t_L g1759 ( 
.A(n_1642),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1681),
.B(n_837),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1730),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1698),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1722),
.B(n_1670),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1699),
.B(n_1165),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1692),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1739),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1692),
.Y(n_1767)
);

BUFx4f_ASAP7_75t_L g1768 ( 
.A(n_1704),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1700),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1705),
.B(n_1689),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1698),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1708),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1700),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1708),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1690),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1720),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1709),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_R g1778 ( 
.A(n_1694),
.B(n_1630),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1720),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_SL g1780 ( 
.A1(n_1726),
.A2(n_1635),
.B1(n_932),
.B2(n_926),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1752),
.B(n_1165),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1760),
.B(n_837),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1695),
.B(n_1565),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1709),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1713),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1713),
.Y(n_1786)
);

BUFx3_ASAP7_75t_L g1787 ( 
.A(n_1704),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1695),
.B(n_1654),
.Y(n_1788)
);

AO22x1_ASAP7_75t_L g1789 ( 
.A1(n_1687),
.A2(n_1370),
.B1(n_1632),
.B2(n_1453),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1710),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1703),
.B(n_1661),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1715),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1751),
.A2(n_1617),
.B1(n_1522),
.B2(n_1607),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1759),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1690),
.Y(n_1795)
);

INVx4_ASAP7_75t_L g1796 ( 
.A(n_1704),
.Y(n_1796)
);

INVx5_ASAP7_75t_L g1797 ( 
.A(n_1704),
.Y(n_1797)
);

INVx3_ASAP7_75t_L g1798 ( 
.A(n_1690),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_1690),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1704),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1696),
.B(n_850),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1688),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1715),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1738),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1745),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1712),
.B(n_855),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1745),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1754),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1691),
.A2(n_1617),
.B1(n_1584),
.B2(n_1577),
.Y(n_1809)
);

INVx2_ASAP7_75t_SL g1810 ( 
.A(n_1688),
.Y(n_1810)
);

BUFx4f_ASAP7_75t_L g1811 ( 
.A(n_1775),
.Y(n_1811)
);

NAND2xp33_ASAP7_75t_SL g1812 ( 
.A(n_1778),
.B(n_1622),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1806),
.B(n_1680),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1793),
.A2(n_1735),
.B1(n_1522),
.B2(n_1751),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1768),
.A2(n_1706),
.B(n_1751),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1791),
.B(n_1728),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1770),
.B(n_1711),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1765),
.Y(n_1818)
);

OAI21xp33_ASAP7_75t_L g1819 ( 
.A1(n_1782),
.A2(n_921),
.B(n_855),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1761),
.Y(n_1820)
);

NOR3xp33_ASAP7_75t_SL g1821 ( 
.A(n_1794),
.B(n_1680),
.C(n_1697),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1764),
.B(n_921),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1763),
.B(n_1728),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1765),
.Y(n_1824)
);

AO21x2_ASAP7_75t_L g1825 ( 
.A1(n_1767),
.A2(n_1744),
.B(n_1684),
.Y(n_1825)
);

INVx4_ASAP7_75t_L g1826 ( 
.A(n_1775),
.Y(n_1826)
);

A2O1A1Ixp33_ASAP7_75t_L g1827 ( 
.A1(n_1793),
.A2(n_1701),
.B(n_1702),
.C(n_1717),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1780),
.A2(n_1753),
.B1(n_1723),
.B2(n_1740),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1767),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1775),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1768),
.A2(n_1693),
.B(n_1719),
.Y(n_1831)
);

O2A1O1Ixp5_ASAP7_75t_L g1832 ( 
.A1(n_1783),
.A2(n_1727),
.B(n_1721),
.C(n_1718),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1769),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1766),
.B(n_1748),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1769),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1773),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1787),
.B(n_1707),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1781),
.B(n_925),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1773),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1801),
.A2(n_1736),
.B(n_1734),
.C(n_1607),
.Y(n_1840)
);

A2O1A1Ixp33_ASAP7_75t_L g1841 ( 
.A1(n_1788),
.A2(n_1584),
.B(n_1681),
.C(n_1616),
.Y(n_1841)
);

INVx6_ASAP7_75t_L g1842 ( 
.A(n_1797),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_SL g1843 ( 
.A1(n_1780),
.A2(n_1635),
.B1(n_1571),
.B2(n_1714),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1777),
.B(n_1807),
.Y(n_1844)
);

OAI21x1_ASAP7_75t_L g1845 ( 
.A1(n_1795),
.A2(n_1586),
.B(n_1574),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1804),
.B(n_1729),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1802),
.B(n_925),
.Y(n_1847)
);

AO32x1_ASAP7_75t_L g1848 ( 
.A1(n_1777),
.A2(n_1786),
.A3(n_1792),
.B1(n_1785),
.B2(n_1784),
.Y(n_1848)
);

A2O1A1Ixp33_ASAP7_75t_L g1849 ( 
.A1(n_1809),
.A2(n_1732),
.B(n_1665),
.C(n_1631),
.Y(n_1849)
);

INVx1_ASAP7_75t_SL g1850 ( 
.A(n_1790),
.Y(n_1850)
);

O2A1O1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1802),
.A2(n_1749),
.B(n_877),
.C(n_922),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1810),
.B(n_1001),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1790),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1787),
.B(n_1707),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1810),
.Y(n_1855)
);

INVx1_ASAP7_75t_SL g1856 ( 
.A(n_1775),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1784),
.Y(n_1857)
);

AOI33xp33_ASAP7_75t_L g1858 ( 
.A1(n_1785),
.A2(n_1023),
.A3(n_958),
.B1(n_954),
.B2(n_1662),
.B3(n_1057),
.Y(n_1858)
);

O2A1O1Ixp5_ASAP7_75t_L g1859 ( 
.A1(n_1789),
.A2(n_1733),
.B(n_1684),
.C(n_1586),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1818),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1824),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1814),
.A2(n_1768),
.B1(n_1796),
.B2(n_1797),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1811),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1829),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1833),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1835),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1817),
.B(n_1758),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1839),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1811),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1843),
.A2(n_1819),
.B1(n_1822),
.B2(n_1838),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1820),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1836),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1857),
.Y(n_1873)
);

BUFx12f_ASAP7_75t_L g1874 ( 
.A(n_1830),
.Y(n_1874)
);

AOI33xp33_ASAP7_75t_L g1875 ( 
.A1(n_1834),
.A2(n_1023),
.A3(n_1060),
.B1(n_1062),
.B2(n_1061),
.B3(n_1052),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1815),
.A2(n_1685),
.B(n_1797),
.Y(n_1876)
);

AND2x6_ASAP7_75t_L g1877 ( 
.A(n_1837),
.B(n_1787),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1844),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1844),
.Y(n_1879)
);

INVxp67_ASAP7_75t_SL g1880 ( 
.A(n_1850),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1850),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1846),
.B(n_1795),
.Y(n_1882)
);

INVx4_ASAP7_75t_L g1883 ( 
.A(n_1830),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1828),
.A2(n_1789),
.B1(n_1516),
.B2(n_1737),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1837),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1854),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1816),
.B(n_1786),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1853),
.Y(n_1888)
);

OAI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1827),
.A2(n_1796),
.B1(n_1797),
.B2(n_1800),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1853),
.B(n_1800),
.Y(n_1890)
);

INVx3_ASAP7_75t_L g1891 ( 
.A(n_1830),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1847),
.A2(n_1516),
.B1(n_1737),
.B2(n_1723),
.Y(n_1892)
);

INVx1_ASAP7_75t_SL g1893 ( 
.A(n_1812),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1854),
.B(n_1800),
.Y(n_1894)
);

OAI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1817),
.A2(n_1796),
.B1(n_1797),
.B2(n_1741),
.Y(n_1895)
);

A2O1A1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1841),
.A2(n_1742),
.B(n_1501),
.C(n_1797),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1823),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1848),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1855),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1848),
.Y(n_1900)
);

INVx5_ASAP7_75t_L g1901 ( 
.A(n_1842),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1840),
.B(n_1792),
.Y(n_1902)
);

BUFx12f_ASAP7_75t_L g1903 ( 
.A(n_1826),
.Y(n_1903)
);

AND2x2_ASAP7_75t_SL g1904 ( 
.A(n_1858),
.B(n_1796),
.Y(n_1904)
);

CKINVDCx20_ASAP7_75t_R g1905 ( 
.A(n_1821),
.Y(n_1905)
);

OA21x2_ASAP7_75t_L g1906 ( 
.A1(n_1845),
.A2(n_1805),
.B(n_1803),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1849),
.B(n_1803),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1826),
.B(n_1856),
.Y(n_1908)
);

AND2x6_ASAP7_75t_L g1909 ( 
.A(n_1856),
.B(n_1742),
.Y(n_1909)
);

BUFx2_ASAP7_75t_L g1910 ( 
.A(n_1842),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1852),
.B(n_1758),
.Y(n_1911)
);

BUFx3_ASAP7_75t_L g1912 ( 
.A(n_1813),
.Y(n_1912)
);

BUFx2_ASAP7_75t_L g1913 ( 
.A(n_1825),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1832),
.A2(n_867),
.B(n_828),
.Y(n_1914)
);

CKINVDCx6p67_ASAP7_75t_R g1915 ( 
.A(n_1851),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1859),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1831),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1829),
.Y(n_1918)
);

BUFx2_ASAP7_75t_L g1919 ( 
.A(n_1820),
.Y(n_1919)
);

NAND2x1p5_ASAP7_75t_L g1920 ( 
.A(n_1850),
.B(n_1795),
.Y(n_1920)
);

A2O1A1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1815),
.A2(n_879),
.B(n_868),
.C(n_1589),
.Y(n_1921)
);

AOI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1814),
.A2(n_1610),
.B1(n_1746),
.B2(n_1704),
.Y(n_1922)
);

NOR2x1_ASAP7_75t_SL g1923 ( 
.A(n_1885),
.B(n_1759),
.Y(n_1923)
);

AO31x2_ASAP7_75t_L g1924 ( 
.A1(n_1913),
.A2(n_1807),
.A3(n_1808),
.B(n_1805),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1882),
.B(n_1795),
.Y(n_1925)
);

O2A1O1Ixp33_ASAP7_75t_SL g1926 ( 
.A1(n_1905),
.A2(n_1001),
.B(n_1003),
.C(n_1067),
.Y(n_1926)
);

O2A1O1Ixp33_ASAP7_75t_SL g1927 ( 
.A1(n_1905),
.A2(n_1003),
.B(n_817),
.C(n_1042),
.Y(n_1927)
);

OAI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1876),
.A2(n_1798),
.B(n_1808),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1881),
.Y(n_1929)
);

AOI22x1_ASAP7_75t_L g1930 ( 
.A1(n_1893),
.A2(n_722),
.B1(n_724),
.B2(n_720),
.Y(n_1930)
);

AO21x1_ASAP7_75t_L g1931 ( 
.A1(n_1867),
.A2(n_1042),
.B(n_854),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1864),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1897),
.B(n_1798),
.Y(n_1933)
);

BUFx2_ASAP7_75t_L g1934 ( 
.A(n_1881),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1871),
.B(n_1798),
.Y(n_1935)
);

O2A1O1Ixp33_ASAP7_75t_SL g1936 ( 
.A1(n_1870),
.A2(n_1642),
.B(n_1588),
.C(n_1595),
.Y(n_1936)
);

O2A1O1Ixp33_ASAP7_75t_L g1937 ( 
.A1(n_1914),
.A2(n_968),
.B(n_792),
.C(n_789),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1871),
.B(n_1919),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1872),
.Y(n_1939)
);

BUFx10_ASAP7_75t_L g1940 ( 
.A(n_1867),
.Y(n_1940)
);

O2A1O1Ixp33_ASAP7_75t_SL g1941 ( 
.A1(n_1911),
.A2(n_1601),
.B(n_1608),
.C(n_1587),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1921),
.A2(n_964),
.B(n_1654),
.Y(n_1942)
);

AOI211xp5_ASAP7_75t_L g1943 ( 
.A1(n_1911),
.A2(n_724),
.B(n_729),
.C(n_722),
.Y(n_1943)
);

NOR2xp67_ASAP7_75t_L g1944 ( 
.A(n_1917),
.B(n_1775),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1918),
.Y(n_1945)
);

BUFx12f_ASAP7_75t_L g1946 ( 
.A(n_1874),
.Y(n_1946)
);

OAI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1884),
.A2(n_733),
.B1(n_742),
.B2(n_731),
.C(n_729),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1873),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1921),
.A2(n_1747),
.B(n_1799),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1909),
.A2(n_1750),
.B1(n_1663),
.B2(n_1724),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1860),
.Y(n_1951)
);

CKINVDCx14_ASAP7_75t_R g1952 ( 
.A(n_1912),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1887),
.B(n_1799),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1909),
.A2(n_1750),
.B1(n_1663),
.B2(n_1724),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1892),
.A2(n_1746),
.B1(n_1654),
.B2(n_1647),
.Y(n_1955)
);

INVx2_ASAP7_75t_SL g1956 ( 
.A(n_1899),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1912),
.B(n_1098),
.Y(n_1957)
);

AO31x2_ASAP7_75t_L g1958 ( 
.A1(n_1916),
.A2(n_1772),
.A3(n_1774),
.B(n_1762),
.Y(n_1958)
);

AOI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1896),
.A2(n_1799),
.B(n_1643),
.Y(n_1959)
);

O2A1O1Ixp33_ASAP7_75t_L g1960 ( 
.A1(n_1896),
.A2(n_780),
.B(n_979),
.C(n_978),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1880),
.B(n_1799),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1885),
.Y(n_1962)
);

INVxp67_ASAP7_75t_L g1963 ( 
.A(n_1888),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1861),
.Y(n_1964)
);

AOI221xp5_ASAP7_75t_L g1965 ( 
.A1(n_1907),
.A2(n_1182),
.B1(n_519),
.B2(n_525),
.C(n_518),
.Y(n_1965)
);

BUFx3_ASAP7_75t_L g1966 ( 
.A(n_1903),
.Y(n_1966)
);

AO32x2_ASAP7_75t_L g1967 ( 
.A1(n_1886),
.A2(n_1181),
.A3(n_1649),
.B1(n_1648),
.B2(n_1638),
.Y(n_1967)
);

O2A1O1Ixp33_ASAP7_75t_SL g1968 ( 
.A1(n_1880),
.A2(n_1902),
.B(n_1865),
.C(n_1868),
.Y(n_1968)
);

AOI32xp33_ASAP7_75t_L g1969 ( 
.A1(n_1875),
.A2(n_742),
.A3(n_745),
.B1(n_733),
.B2(n_731),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_L g1970 ( 
.A(n_1915),
.B(n_9),
.Y(n_1970)
);

O2A1O1Ixp5_ASAP7_75t_L g1971 ( 
.A1(n_1889),
.A2(n_854),
.B(n_853),
.C(n_951),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1895),
.A2(n_1799),
.B(n_1466),
.Y(n_1972)
);

OAI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1904),
.A2(n_1102),
.B(n_939),
.Y(n_1973)
);

O2A1O1Ixp33_ASAP7_75t_SL g1974 ( 
.A1(n_1866),
.A2(n_1621),
.B(n_1633),
.C(n_1619),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1890),
.B(n_1690),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1873),
.B(n_936),
.Y(n_1976)
);

O2A1O1Ixp33_ASAP7_75t_SL g1977 ( 
.A1(n_1878),
.A2(n_1641),
.B(n_1656),
.C(n_1639),
.Y(n_1977)
);

OAI21x1_ASAP7_75t_L g1978 ( 
.A1(n_1862),
.A2(n_1476),
.B(n_1771),
.Y(n_1978)
);

AOI21xp5_ASAP7_75t_L g1979 ( 
.A1(n_1895),
.A2(n_1466),
.B(n_1442),
.Y(n_1979)
);

INVx5_ASAP7_75t_L g1980 ( 
.A(n_1877),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1920),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1879),
.Y(n_1982)
);

A2O1A1Ixp33_ASAP7_75t_L g1983 ( 
.A1(n_1875),
.A2(n_1663),
.B(n_974),
.C(n_929),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1904),
.A2(n_1442),
.B(n_1716),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1910),
.Y(n_1985)
);

AND2x6_ASAP7_75t_L g1986 ( 
.A(n_1894),
.B(n_1772),
.Y(n_1986)
);

A2O1A1Ixp33_ASAP7_75t_L g1987 ( 
.A1(n_1922),
.A2(n_746),
.B(n_768),
.C(n_752),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1863),
.B(n_1370),
.Y(n_1988)
);

OAI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1920),
.A2(n_981),
.B(n_980),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1906),
.Y(n_1990)
);

CKINVDCx6p67_ASAP7_75t_R g1991 ( 
.A(n_1863),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1908),
.A2(n_1731),
.B(n_1716),
.Y(n_1992)
);

O2A1O1Ixp33_ASAP7_75t_SL g1993 ( 
.A1(n_1891),
.A2(n_1667),
.B(n_1673),
.C(n_1664),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1906),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1863),
.A2(n_746),
.B1(n_752),
.B2(n_745),
.Y(n_1995)
);

O2A1O1Ixp33_ASAP7_75t_SL g1996 ( 
.A1(n_1891),
.A2(n_1676),
.B(n_1675),
.C(n_1678),
.Y(n_1996)
);

OAI21x1_ASAP7_75t_L g1997 ( 
.A1(n_1906),
.A2(n_1900),
.B(n_1898),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1908),
.Y(n_1998)
);

AOI221xp5_ASAP7_75t_L g1999 ( 
.A1(n_1894),
.A2(n_536),
.B1(n_538),
.B2(n_526),
.C(n_515),
.Y(n_1999)
);

OAI31xp33_ASAP7_75t_SL g2000 ( 
.A1(n_1909),
.A2(n_12),
.A3(n_10),
.B(n_11),
.Y(n_2000)
);

NAND2x1p5_ASAP7_75t_L g2001 ( 
.A(n_1863),
.B(n_1567),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1909),
.B(n_1883),
.Y(n_2002)
);

O2A1O1Ixp33_ASAP7_75t_SL g2003 ( 
.A1(n_1883),
.A2(n_1683),
.B(n_1686),
.C(n_1682),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1909),
.B(n_1776),
.Y(n_2004)
);

AOI22xp33_ASAP7_75t_L g2005 ( 
.A1(n_1942),
.A2(n_1877),
.B1(n_1755),
.B2(n_1756),
.Y(n_2005)
);

OAI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1937),
.A2(n_759),
.B(n_756),
.Y(n_2006)
);

INVxp67_ASAP7_75t_L g2007 ( 
.A(n_1934),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1929),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1940),
.B(n_1901),
.Y(n_2009)
);

AOI22xp33_ASAP7_75t_L g2010 ( 
.A1(n_1931),
.A2(n_1877),
.B1(n_1041),
.B2(n_1659),
.Y(n_2010)
);

BUFx12f_ASAP7_75t_L g2011 ( 
.A(n_1946),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_SL g2012 ( 
.A1(n_1940),
.A2(n_1877),
.B1(n_1186),
.B2(n_1187),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1951),
.Y(n_2013)
);

NAND2xp33_ASAP7_75t_L g2014 ( 
.A(n_1969),
.B(n_1869),
.Y(n_2014)
);

AOI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1947),
.A2(n_1877),
.B1(n_1755),
.B2(n_1756),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1963),
.B(n_1938),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1964),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1962),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1982),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_1952),
.B(n_1869),
.Y(n_2020)
);

INVx3_ASAP7_75t_L g2021 ( 
.A(n_1962),
.Y(n_2021)
);

AOI22xp33_ASAP7_75t_L g2022 ( 
.A1(n_1970),
.A2(n_1041),
.B1(n_1659),
.B2(n_1657),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1948),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1956),
.B(n_1901),
.Y(n_2024)
);

INVx2_ASAP7_75t_SL g2025 ( 
.A(n_1985),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1935),
.B(n_936),
.Y(n_2026)
);

OAI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1955),
.A2(n_1901),
.B1(n_1869),
.B2(n_759),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1976),
.Y(n_2028)
);

INVx6_ASAP7_75t_L g2029 ( 
.A(n_1980),
.Y(n_2029)
);

INVx6_ASAP7_75t_L g2030 ( 
.A(n_1980),
.Y(n_2030)
);

HB1xp67_ASAP7_75t_L g2031 ( 
.A(n_1997),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1924),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1987),
.A2(n_1869),
.B1(n_1901),
.B2(n_771),
.Y(n_2033)
);

AOI221xp5_ASAP7_75t_L g2034 ( 
.A1(n_1969),
.A2(n_766),
.B1(n_768),
.B2(n_761),
.C(n_756),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_1998),
.B(n_936),
.Y(n_2035)
);

OAI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1955),
.A2(n_774),
.B1(n_766),
.B2(n_771),
.Y(n_2036)
);

INVx4_ASAP7_75t_L g2037 ( 
.A(n_1966),
.Y(n_2037)
);

INVx4_ASAP7_75t_L g2038 ( 
.A(n_1991),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1957),
.Y(n_2039)
);

AOI22xp33_ASAP7_75t_L g2040 ( 
.A1(n_1950),
.A2(n_1954),
.B1(n_1965),
.B2(n_2004),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1924),
.Y(n_2041)
);

NAND2x1p5_ASAP7_75t_L g2042 ( 
.A(n_1980),
.B(n_1567),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_2004),
.A2(n_1973),
.B1(n_1986),
.B2(n_1932),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1924),
.Y(n_2044)
);

INVx2_ASAP7_75t_SL g2045 ( 
.A(n_1925),
.Y(n_2045)
);

AND2x2_ASAP7_75t_SL g2046 ( 
.A(n_2000),
.B(n_1725),
.Y(n_2046)
);

AOI221xp5_ASAP7_75t_L g2047 ( 
.A1(n_1943),
.A2(n_774),
.B1(n_775),
.B2(n_772),
.C(n_761),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1939),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1986),
.A2(n_1945),
.B1(n_1999),
.B2(n_1930),
.Y(n_2049)
);

HB1xp67_ASAP7_75t_L g2050 ( 
.A(n_1994),
.Y(n_2050)
);

AOI22xp33_ASAP7_75t_SL g2051 ( 
.A1(n_2000),
.A2(n_1186),
.B1(n_1187),
.B2(n_1173),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1986),
.A2(n_1757),
.B1(n_1754),
.B2(n_1776),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1953),
.B(n_982),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1968),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1961),
.B(n_902),
.Y(n_2055)
);

BUFx4_ASAP7_75t_SL g2056 ( 
.A(n_1926),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_1986),
.A2(n_1757),
.B1(n_1779),
.B2(n_1651),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1949),
.A2(n_1779),
.B1(n_1651),
.B2(n_1660),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1958),
.Y(n_2059)
);

NAND2xp33_ASAP7_75t_L g2060 ( 
.A(n_2002),
.B(n_772),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1958),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_1959),
.A2(n_1660),
.B1(n_1672),
.B2(n_1646),
.Y(n_2062)
);

INVx6_ASAP7_75t_L g2063 ( 
.A(n_1975),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1933),
.B(n_985),
.Y(n_2064)
);

HB1xp67_ASAP7_75t_L g2065 ( 
.A(n_2050),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_2037),
.B(n_1936),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2050),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2032),
.Y(n_2068)
);

AO21x2_ASAP7_75t_L g2069 ( 
.A1(n_2041),
.A2(n_1990),
.B(n_1944),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_2011),
.Y(n_2070)
);

INVxp67_ASAP7_75t_SL g2071 ( 
.A(n_2031),
.Y(n_2071)
);

OAI21x1_ASAP7_75t_L g2072 ( 
.A1(n_2044),
.A2(n_2054),
.B(n_2031),
.Y(n_2072)
);

CKINVDCx20_ASAP7_75t_R g2073 ( 
.A(n_2039),
.Y(n_2073)
);

BUFx2_ASAP7_75t_L g2074 ( 
.A(n_2007),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_2051),
.A2(n_1943),
.B1(n_1960),
.B2(n_1983),
.Y(n_2075)
);

CKINVDCx16_ASAP7_75t_R g2076 ( 
.A(n_2037),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2008),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2059),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2013),
.Y(n_2079)
);

INVx1_ASAP7_75t_SL g2080 ( 
.A(n_2026),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_2061),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2017),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2019),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_2007),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2028),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2035),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2023),
.Y(n_2087)
);

CKINVDCx20_ASAP7_75t_R g2088 ( 
.A(n_2025),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2016),
.B(n_1981),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2055),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2045),
.B(n_1981),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2053),
.Y(n_2092)
);

OAI21x1_ASAP7_75t_L g2093 ( 
.A1(n_2043),
.A2(n_1928),
.B(n_1978),
.Y(n_2093)
);

AOI21x1_ASAP7_75t_L g2094 ( 
.A1(n_2064),
.A2(n_1944),
.B(n_1972),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_2020),
.B(n_1927),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2048),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2018),
.Y(n_2097)
);

OAI21xp5_ASAP7_75t_L g2098 ( 
.A1(n_2051),
.A2(n_1941),
.B(n_1971),
.Y(n_2098)
);

HB1xp67_ASAP7_75t_L g2099 ( 
.A(n_2018),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_2070),
.Y(n_2100)
);

BUFx3_ASAP7_75t_L g2101 ( 
.A(n_2070),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_2073),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2078),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2080),
.B(n_2021),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2074),
.B(n_2021),
.Y(n_2105)
);

AOI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_2075),
.A2(n_2014),
.B1(n_2046),
.B2(n_2036),
.Y(n_2106)
);

OAI221xp5_ASAP7_75t_L g2107 ( 
.A1(n_2075),
.A2(n_2006),
.B1(n_2012),
.B2(n_2049),
.C(n_2022),
.Y(n_2107)
);

INVx11_ASAP7_75t_L g2108 ( 
.A(n_2070),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2074),
.B(n_2024),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2080),
.B(n_2024),
.Y(n_2110)
);

AOI221xp5_ASAP7_75t_L g2111 ( 
.A1(n_2092),
.A2(n_2034),
.B1(n_2047),
.B2(n_2022),
.C(n_775),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2092),
.B(n_1977),
.Y(n_2112)
);

AOI22xp33_ASAP7_75t_L g2113 ( 
.A1(n_2086),
.A2(n_2046),
.B1(n_2098),
.B2(n_2090),
.Y(n_2113)
);

AND2x4_ASAP7_75t_L g2114 ( 
.A(n_2072),
.B(n_2009),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2079),
.Y(n_2115)
);

AOI22xp33_ASAP7_75t_L g2116 ( 
.A1(n_2086),
.A2(n_2005),
.B1(n_2040),
.B2(n_2012),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_2098),
.A2(n_2027),
.B1(n_2010),
.B2(n_2057),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2090),
.B(n_1974),
.Y(n_2118)
);

NAND2x1_ASAP7_75t_L g2119 ( 
.A(n_2067),
.B(n_2029),
.Y(n_2119)
);

OAI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_2076),
.A2(n_2038),
.B1(n_2063),
.B2(n_2027),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_2094),
.Y(n_2121)
);

HB1xp67_ASAP7_75t_L g2122 ( 
.A(n_2084),
.Y(n_2122)
);

OA21x2_ASAP7_75t_L g2123 ( 
.A1(n_2072),
.A2(n_2052),
.B(n_2058),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2096),
.A2(n_2095),
.B1(n_2085),
.B2(n_2087),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2109),
.B(n_2084),
.Y(n_2125)
);

AND2x4_ASAP7_75t_L g2126 ( 
.A(n_2114),
.B(n_2072),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2112),
.B(n_2085),
.Y(n_2127)
);

AOI22xp33_ASAP7_75t_L g2128 ( 
.A1(n_2107),
.A2(n_2096),
.B1(n_2087),
.B2(n_2083),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2115),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2115),
.Y(n_2130)
);

AOI21xp5_ASAP7_75t_SL g2131 ( 
.A1(n_2106),
.A2(n_2066),
.B(n_1923),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2109),
.B(n_2105),
.Y(n_2132)
);

INVxp67_ASAP7_75t_L g2133 ( 
.A(n_2101),
.Y(n_2133)
);

BUFx6f_ASAP7_75t_L g2134 ( 
.A(n_2100),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2105),
.B(n_2099),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2122),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2124),
.B(n_2079),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2100),
.B(n_2076),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2118),
.B(n_2082),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_2104),
.B(n_2067),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2100),
.B(n_2091),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2110),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2121),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2106),
.A2(n_2010),
.B1(n_2060),
.B2(n_2015),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2100),
.B(n_2091),
.Y(n_2145)
);

INVx3_ASAP7_75t_L g2146 ( 
.A(n_2121),
.Y(n_2146)
);

AOI221xp5_ASAP7_75t_L g2147 ( 
.A1(n_2113),
.A2(n_2071),
.B1(n_2083),
.B2(n_2065),
.C(n_2068),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2100),
.B(n_2065),
.Y(n_2148)
);

INVx2_ASAP7_75t_SL g2149 ( 
.A(n_2108),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2121),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2114),
.B(n_2119),
.Y(n_2151)
);

INVxp67_ASAP7_75t_L g2152 ( 
.A(n_2101),
.Y(n_2152)
);

AOI22xp33_ASAP7_75t_L g2153 ( 
.A1(n_2121),
.A2(n_2096),
.B1(n_2068),
.B2(n_2069),
.Y(n_2153)
);

HB1xp67_ASAP7_75t_L g2154 ( 
.A(n_2121),
.Y(n_2154)
);

NOR2xp67_ASAP7_75t_L g2155 ( 
.A(n_2114),
.B(n_2038),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_2119),
.B(n_2077),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2134),
.Y(n_2157)
);

AOI22xp33_ASAP7_75t_L g2158 ( 
.A1(n_2128),
.A2(n_2123),
.B1(n_2117),
.B2(n_2116),
.Y(n_2158)
);

OR2x2_ASAP7_75t_L g2159 ( 
.A(n_2142),
.B(n_2089),
.Y(n_2159)
);

HB1xp67_ASAP7_75t_L g2160 ( 
.A(n_2125),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_2138),
.B(n_2088),
.Y(n_2161)
);

AOI221xp5_ASAP7_75t_L g2162 ( 
.A1(n_2137),
.A2(n_2071),
.B1(n_2111),
.B2(n_2120),
.C(n_2103),
.Y(n_2162)
);

AOI33xp33_ASAP7_75t_L g2163 ( 
.A1(n_2147),
.A2(n_2082),
.A3(n_2077),
.B1(n_2097),
.B2(n_2056),
.B3(n_909),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2134),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_2138),
.B(n_2102),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2142),
.B(n_2089),
.Y(n_2166)
);

NOR3xp33_ASAP7_75t_L g2167 ( 
.A(n_2146),
.B(n_2033),
.C(n_2102),
.Y(n_2167)
);

AOI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_2144),
.A2(n_2123),
.B1(n_2069),
.B2(n_2068),
.Y(n_2168)
);

AOI32xp33_ASAP7_75t_L g2169 ( 
.A1(n_2126),
.A2(n_2093),
.A3(n_2103),
.B1(n_2056),
.B2(n_1995),
.Y(n_2169)
);

AO31x2_ASAP7_75t_L g2170 ( 
.A1(n_2150),
.A2(n_2081),
.A3(n_2078),
.B(n_2108),
.Y(n_2170)
);

INVxp67_ASAP7_75t_L g2171 ( 
.A(n_2149),
.Y(n_2171)
);

AOI221xp5_ASAP7_75t_L g2172 ( 
.A1(n_2153),
.A2(n_908),
.B1(n_910),
.B2(n_905),
.C(n_904),
.Y(n_2172)
);

INVxp67_ASAP7_75t_L g2173 ( 
.A(n_2149),
.Y(n_2173)
);

OAI221xp5_ASAP7_75t_SL g2174 ( 
.A1(n_2144),
.A2(n_2097),
.B1(n_1984),
.B2(n_2062),
.C(n_1979),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_2134),
.Y(n_2175)
);

OAI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_2155),
.A2(n_2123),
.B1(n_2094),
.B2(n_2030),
.Y(n_2176)
);

AOI211xp5_ASAP7_75t_SL g2177 ( 
.A1(n_2131),
.A2(n_2003),
.B(n_1996),
.C(n_1993),
.Y(n_2177)
);

OAI221xp5_ASAP7_75t_L g2178 ( 
.A1(n_2127),
.A2(n_2131),
.B1(n_2139),
.B2(n_2155),
.C(n_2150),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2160),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2163),
.B(n_2133),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2165),
.B(n_2132),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_2171),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2165),
.B(n_2152),
.Y(n_2183)
);

INVxp67_ASAP7_75t_SL g2184 ( 
.A(n_2167),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2166),
.B(n_2136),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2161),
.B(n_2125),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2161),
.B(n_2132),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2173),
.B(n_2141),
.Y(n_2188)
);

AND2x4_ASAP7_75t_L g2189 ( 
.A(n_2175),
.B(n_2151),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2162),
.B(n_2136),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_2170),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2159),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2157),
.B(n_2141),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2168),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2170),
.Y(n_2195)
);

INVx2_ASAP7_75t_SL g2196 ( 
.A(n_2181),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2179),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_2182),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2187),
.B(n_2134),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2179),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2184),
.B(n_2158),
.Y(n_2201)
);

OAI33xp33_ASAP7_75t_L g2202 ( 
.A1(n_2190),
.A2(n_2176),
.A3(n_2143),
.B1(n_2164),
.B2(n_2130),
.B3(n_2129),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2192),
.Y(n_2203)
);

INVx1_ASAP7_75t_SL g2204 ( 
.A(n_2181),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2199),
.B(n_2187),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2198),
.B(n_2188),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2196),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2199),
.B(n_2188),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2200),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_2204),
.B(n_2183),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2196),
.B(n_2186),
.Y(n_2211)
);

AND2x2_ASAP7_75t_SL g2212 ( 
.A(n_2206),
.B(n_2201),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2208),
.B(n_2203),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2205),
.B(n_2193),
.Y(n_2214)
);

AOI211xp5_ASAP7_75t_L g2215 ( 
.A1(n_2210),
.A2(n_2202),
.B(n_2178),
.C(n_2194),
.Y(n_2215)
);

NAND2x1_ASAP7_75t_L g2216 ( 
.A(n_2207),
.B(n_2189),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2214),
.Y(n_2217)
);

AOI33xp33_ASAP7_75t_L g2218 ( 
.A1(n_2215),
.A2(n_2197),
.A3(n_2200),
.B1(n_2209),
.B2(n_2211),
.B3(n_2194),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2212),
.B(n_2210),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2219),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2217),
.Y(n_2221)
);

O2A1O1Ixp33_ASAP7_75t_L g2222 ( 
.A1(n_2220),
.A2(n_2206),
.B(n_2213),
.C(n_2216),
.Y(n_2222)
);

OAI221xp5_ASAP7_75t_L g2223 ( 
.A1(n_2220),
.A2(n_2169),
.B1(n_2191),
.B2(n_2195),
.C(n_2180),
.Y(n_2223)
);

OA22x2_ASAP7_75t_L g2224 ( 
.A1(n_2222),
.A2(n_2221),
.B1(n_2189),
.B2(n_2218),
.Y(n_2224)
);

AOI22xp33_ASAP7_75t_SL g2225 ( 
.A1(n_2223),
.A2(n_2191),
.B1(n_2195),
.B2(n_2218),
.Y(n_2225)
);

INVx2_ASAP7_75t_SL g2226 ( 
.A(n_2224),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2225),
.Y(n_2227)
);

INVxp67_ASAP7_75t_SL g2228 ( 
.A(n_2224),
.Y(n_2228)
);

NAND2x1_ASAP7_75t_L g2229 ( 
.A(n_2226),
.B(n_2189),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2228),
.Y(n_2230)
);

XOR2x2_ASAP7_75t_L g2231 ( 
.A(n_2227),
.B(n_2177),
.Y(n_2231)
);

AOI221xp5_ASAP7_75t_L g2232 ( 
.A1(n_2227),
.A2(n_2143),
.B1(n_2146),
.B2(n_2154),
.C(n_2172),
.Y(n_2232)
);

NAND4xp75_ASAP7_75t_L g2233 ( 
.A(n_2230),
.B(n_971),
.C(n_973),
.D(n_970),
.Y(n_2233)
);

OR2x2_ASAP7_75t_L g2234 ( 
.A(n_2229),
.B(n_2185),
.Y(n_2234)
);

AND3x1_ASAP7_75t_L g2235 ( 
.A(n_2232),
.B(n_2146),
.C(n_2193),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2234),
.B(n_2233),
.Y(n_2236)
);

AOI221xp5_ASAP7_75t_L g2237 ( 
.A1(n_2235),
.A2(n_2231),
.B1(n_2146),
.B2(n_2175),
.C(n_2185),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2234),
.Y(n_2238)
);

AOI221xp5_ASAP7_75t_L g2239 ( 
.A1(n_2235),
.A2(n_2126),
.B1(n_977),
.B2(n_976),
.C(n_2134),
.Y(n_2239)
);

XNOR2xp5_ASAP7_75t_L g2240 ( 
.A(n_2233),
.B(n_1988),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2234),
.B(n_2170),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2234),
.Y(n_2242)
);

NOR4xp75_ASAP7_75t_L g2243 ( 
.A(n_2233),
.B(n_2151),
.C(n_2148),
.D(n_2145),
.Y(n_2243)
);

AOI21xp33_ASAP7_75t_L g2244 ( 
.A1(n_2234),
.A2(n_783),
.B(n_782),
.Y(n_2244)
);

XNOR2x1_ASAP7_75t_L g2245 ( 
.A(n_2233),
.B(n_1659),
.Y(n_2245)
);

AOI22xp33_ASAP7_75t_L g2246 ( 
.A1(n_2234),
.A2(n_2126),
.B1(n_2148),
.B2(n_2130),
.Y(n_2246)
);

AOI211xp5_ASAP7_75t_L g2247 ( 
.A1(n_2234),
.A2(n_912),
.B(n_915),
.C(n_911),
.Y(n_2247)
);

AOI31xp33_ASAP7_75t_L g2248 ( 
.A1(n_2234),
.A2(n_608),
.A3(n_628),
.B(n_595),
.Y(n_2248)
);

AOI322xp5_ASAP7_75t_L g2249 ( 
.A1(n_2235),
.A2(n_2126),
.A3(n_2174),
.B1(n_2145),
.B2(n_2129),
.C1(n_930),
.C2(n_927),
.Y(n_2249)
);

NAND3xp33_ASAP7_75t_L g2250 ( 
.A(n_2238),
.B(n_2242),
.C(n_2247),
.Y(n_2250)
);

NOR2x1_ASAP7_75t_L g2251 ( 
.A(n_2248),
.B(n_917),
.Y(n_2251)
);

NAND3x1_ASAP7_75t_L g2252 ( 
.A(n_2236),
.B(n_2135),
.C(n_920),
.Y(n_2252)
);

NAND3xp33_ASAP7_75t_L g2253 ( 
.A(n_2244),
.B(n_933),
.C(n_919),
.Y(n_2253)
);

NOR3xp33_ASAP7_75t_L g2254 ( 
.A(n_2239),
.B(n_942),
.C(n_935),
.Y(n_2254)
);

AOI211x1_ASAP7_75t_L g2255 ( 
.A1(n_2243),
.A2(n_2135),
.B(n_937),
.C(n_940),
.Y(n_2255)
);

NOR2x1_ASAP7_75t_L g2256 ( 
.A(n_2241),
.B(n_934),
.Y(n_2256)
);

NAND3xp33_ASAP7_75t_L g2257 ( 
.A(n_2237),
.B(n_944),
.C(n_943),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2245),
.Y(n_2258)
);

NOR2x1_ASAP7_75t_L g2259 ( 
.A(n_2240),
.B(n_946),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2246),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2249),
.B(n_947),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2248),
.B(n_949),
.Y(n_2262)
);

NOR3xp33_ASAP7_75t_L g2263 ( 
.A(n_2238),
.B(n_805),
.C(n_793),
.Y(n_2263)
);

NAND4xp75_ASAP7_75t_L g2264 ( 
.A(n_2238),
.B(n_794),
.C(n_795),
.D(n_788),
.Y(n_2264)
);

NOR2x1_ASAP7_75t_L g2265 ( 
.A(n_2238),
.B(n_801),
.Y(n_2265)
);

NAND3x1_ASAP7_75t_L g2266 ( 
.A(n_2238),
.B(n_1989),
.C(n_804),
.Y(n_2266)
);

AND2x4_ASAP7_75t_L g2267 ( 
.A(n_2238),
.B(n_2156),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_2238),
.B(n_802),
.Y(n_2268)
);

XNOR2x1_ASAP7_75t_L g2269 ( 
.A(n_2238),
.B(n_1576),
.Y(n_2269)
);

NAND3xp33_ASAP7_75t_SL g2270 ( 
.A(n_2238),
.B(n_807),
.C(n_613),
.Y(n_2270)
);

NAND3xp33_ASAP7_75t_L g2271 ( 
.A(n_2238),
.B(n_544),
.C(n_539),
.Y(n_2271)
);

NOR2x1_ASAP7_75t_L g2272 ( 
.A(n_2238),
.B(n_987),
.Y(n_2272)
);

NOR2x1p5_ASAP7_75t_L g2273 ( 
.A(n_2238),
.B(n_547),
.Y(n_2273)
);

NOR3xp33_ASAP7_75t_L g2274 ( 
.A(n_2238),
.B(n_551),
.C(n_549),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2238),
.B(n_2140),
.Y(n_2275)
);

HB1xp67_ASAP7_75t_L g2276 ( 
.A(n_2238),
.Y(n_2276)
);

NOR2x1_ASAP7_75t_L g2277 ( 
.A(n_2238),
.B(n_991),
.Y(n_2277)
);

NAND4xp25_ASAP7_75t_L g2278 ( 
.A(n_2238),
.B(n_994),
.C(n_996),
.D(n_992),
.Y(n_2278)
);

NAND3x2_ASAP7_75t_L g2279 ( 
.A(n_2238),
.B(n_2156),
.C(n_2140),
.Y(n_2279)
);

OAI22xp33_ASAP7_75t_L g2280 ( 
.A1(n_2238),
.A2(n_565),
.B1(n_567),
.B2(n_561),
.Y(n_2280)
);

XOR2xp5_ASAP7_75t_L g2281 ( 
.A(n_2238),
.B(n_576),
.Y(n_2281)
);

INVx1_ASAP7_75t_SL g2282 ( 
.A(n_2238),
.Y(n_2282)
);

NOR3xp33_ASAP7_75t_L g2283 ( 
.A(n_2238),
.B(n_583),
.C(n_579),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2238),
.B(n_2123),
.Y(n_2284)
);

NOR3xp33_ASAP7_75t_L g2285 ( 
.A(n_2238),
.B(n_588),
.C(n_587),
.Y(n_2285)
);

AOI211xp5_ASAP7_75t_L g2286 ( 
.A1(n_2238),
.A2(n_596),
.B(n_601),
.C(n_591),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_2238),
.B(n_10),
.Y(n_2287)
);

NOR3xp33_ASAP7_75t_L g2288 ( 
.A(n_2238),
.B(n_618),
.C(n_605),
.Y(n_2288)
);

NOR3xp33_ASAP7_75t_SL g2289 ( 
.A(n_2238),
.B(n_622),
.C(n_621),
.Y(n_2289)
);

NOR3x1_ASAP7_75t_L g2290 ( 
.A(n_2238),
.B(n_998),
.C(n_997),
.Y(n_2290)
);

AOI211xp5_ASAP7_75t_L g2291 ( 
.A1(n_2238),
.A2(n_630),
.B(n_631),
.C(n_626),
.Y(n_2291)
);

NOR2x1p5_ASAP7_75t_L g2292 ( 
.A(n_2238),
.B(n_632),
.Y(n_2292)
);

NAND3xp33_ASAP7_75t_SL g2293 ( 
.A(n_2238),
.B(n_668),
.C(n_649),
.Y(n_2293)
);

NOR2xp67_ASAP7_75t_L g2294 ( 
.A(n_2238),
.B(n_13),
.Y(n_2294)
);

AOI22xp33_ASAP7_75t_SL g2295 ( 
.A1(n_2276),
.A2(n_648),
.B1(n_655),
.B2(n_635),
.Y(n_2295)
);

HB1xp67_ASAP7_75t_L g2296 ( 
.A(n_2294),
.Y(n_2296)
);

AOI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_2282),
.A2(n_664),
.B1(n_667),
.B2(n_657),
.Y(n_2297)
);

NOR2xp67_ASAP7_75t_L g2298 ( 
.A(n_2293),
.B(n_13),
.Y(n_2298)
);

NAND5xp2_ASAP7_75t_L g2299 ( 
.A(n_2289),
.B(n_2001),
.C(n_2042),
.D(n_1008),
.E(n_1010),
.Y(n_2299)
);

NOR3xp33_ASAP7_75t_L g2300 ( 
.A(n_2250),
.B(n_677),
.C(n_674),
.Y(n_2300)
);

AOI322xp5_ASAP7_75t_L g2301 ( 
.A1(n_2275),
.A2(n_686),
.A3(n_687),
.B1(n_679),
.B2(n_1967),
.C1(n_1014),
.C2(n_1004),
.Y(n_2301)
);

XNOR2xp5_ASAP7_75t_L g2302 ( 
.A(n_2269),
.B(n_14),
.Y(n_2302)
);

AOI211xp5_ASAP7_75t_L g2303 ( 
.A1(n_2260),
.A2(n_1016),
.B(n_1017),
.C(n_999),
.Y(n_2303)
);

AO22x2_ASAP7_75t_L g2304 ( 
.A1(n_2281),
.A2(n_1018),
.B1(n_1020),
.B2(n_1019),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2251),
.Y(n_2305)
);

AO22x2_ASAP7_75t_L g2306 ( 
.A1(n_2270),
.A2(n_1021),
.B1(n_1027),
.B2(n_1022),
.Y(n_2306)
);

OAI221xp5_ASAP7_75t_L g2307 ( 
.A1(n_2286),
.A2(n_1028),
.B1(n_1007),
.B2(n_1629),
.C(n_1625),
.Y(n_2307)
);

XNOR2xp5_ASAP7_75t_L g2308 ( 
.A(n_2252),
.B(n_14),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2267),
.Y(n_2309)
);

AOI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_2267),
.A2(n_1625),
.B1(n_1637),
.B2(n_1629),
.Y(n_2310)
);

AO22x2_ASAP7_75t_L g2311 ( 
.A1(n_2264),
.A2(n_1007),
.B1(n_1648),
.B2(n_1638),
.Y(n_2311)
);

OAI211xp5_ASAP7_75t_SL g2312 ( 
.A1(n_2291),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_2312)
);

NOR4xp75_ASAP7_75t_L g2313 ( 
.A(n_2262),
.B(n_17),
.C(n_15),
.D(n_16),
.Y(n_2313)
);

AOI322xp5_ASAP7_75t_L g2314 ( 
.A1(n_2284),
.A2(n_1967),
.A3(n_1725),
.B1(n_1640),
.B2(n_1637),
.C1(n_2081),
.C2(n_2078),
.Y(n_2314)
);

OAI22xp5_ASAP7_75t_SL g2315 ( 
.A1(n_2255),
.A2(n_1649),
.B1(n_469),
.B2(n_473),
.Y(n_2315)
);

OAI211xp5_ASAP7_75t_SL g2316 ( 
.A1(n_2258),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_2316)
);

AOI21xp5_ASAP7_75t_L g2317 ( 
.A1(n_2280),
.A2(n_469),
.B(n_460),
.Y(n_2317)
);

A2O1A1Ixp33_ASAP7_75t_L g2318 ( 
.A1(n_2271),
.A2(n_1640),
.B(n_473),
.C(n_475),
.Y(n_2318)
);

AOI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_2274),
.A2(n_1725),
.B1(n_1387),
.B2(n_1251),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2287),
.Y(n_2320)
);

AOI211xp5_ASAP7_75t_L g2321 ( 
.A1(n_2283),
.A2(n_475),
.B(n_477),
.C(n_460),
.Y(n_2321)
);

AOI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2285),
.A2(n_1251),
.B1(n_1533),
.B2(n_478),
.Y(n_2322)
);

AOI311xp33_ASAP7_75t_L g2323 ( 
.A1(n_2288),
.A2(n_26),
.A3(n_23),
.B(n_24),
.C(n_27),
.Y(n_2323)
);

AOI211xp5_ASAP7_75t_L g2324 ( 
.A1(n_2257),
.A2(n_478),
.B(n_486),
.C(n_477),
.Y(n_2324)
);

AOI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_2273),
.A2(n_1251),
.B1(n_1533),
.B2(n_490),
.Y(n_2325)
);

OAI211xp5_ASAP7_75t_L g2326 ( 
.A1(n_2261),
.A2(n_490),
.B(n_493),
.C(n_486),
.Y(n_2326)
);

AOI322xp5_ASAP7_75t_L g2327 ( 
.A1(n_2268),
.A2(n_2259),
.A3(n_2272),
.B1(n_2277),
.B2(n_2265),
.C1(n_2256),
.C2(n_2263),
.Y(n_2327)
);

NOR4xp25_ASAP7_75t_L g2328 ( 
.A(n_2278),
.B(n_1545),
.C(n_1542),
.D(n_32),
.Y(n_2328)
);

BUFx2_ASAP7_75t_L g2329 ( 
.A(n_2287),
.Y(n_2329)
);

AOI211xp5_ASAP7_75t_L g2330 ( 
.A1(n_2254),
.A2(n_499),
.B(n_692),
.C(n_493),
.Y(n_2330)
);

AOI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2292),
.A2(n_1251),
.B1(n_499),
.B2(n_695),
.Y(n_2331)
);

O2A1O1Ixp33_ASAP7_75t_L g2332 ( 
.A1(n_2253),
.A2(n_1545),
.B(n_1542),
.C(n_1204),
.Y(n_2332)
);

AOI21xp5_ASAP7_75t_L g2333 ( 
.A1(n_2290),
.A2(n_695),
.B(n_692),
.Y(n_2333)
);

AOI22xp5_ASAP7_75t_L g2334 ( 
.A1(n_2279),
.A2(n_1251),
.B1(n_705),
.B2(n_707),
.Y(n_2334)
);

INVx1_ASAP7_75t_SL g2335 ( 
.A(n_2266),
.Y(n_2335)
);

AOI21xp5_ASAP7_75t_L g2336 ( 
.A1(n_2282),
.A2(n_705),
.B(n_701),
.Y(n_2336)
);

OAI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2276),
.A2(n_1204),
.B(n_1189),
.Y(n_2337)
);

XNOR2xp5_ASAP7_75t_L g2338 ( 
.A(n_2276),
.B(n_29),
.Y(n_2338)
);

AOI21xp33_ASAP7_75t_SL g2339 ( 
.A1(n_2276),
.A2(n_31),
.B(n_33),
.Y(n_2339)
);

O2A1O1Ixp33_ASAP7_75t_L g2340 ( 
.A1(n_2276),
.A2(n_1204),
.B(n_1248),
.C(n_1189),
.Y(n_2340)
);

AOI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2282),
.A2(n_707),
.B1(n_709),
.B2(n_701),
.Y(n_2341)
);

HB1xp67_ASAP7_75t_L g2342 ( 
.A(n_2294),
.Y(n_2342)
);

OAI322xp33_ASAP7_75t_L g2343 ( 
.A1(n_2282),
.A2(n_732),
.A3(n_719),
.B1(n_736),
.B2(n_738),
.C1(n_730),
.C2(n_710),
.Y(n_2343)
);

AND4x1_ASAP7_75t_L g2344 ( 
.A(n_2289),
.B(n_36),
.C(n_31),
.D(n_34),
.Y(n_2344)
);

OA22x2_ASAP7_75t_L g2345 ( 
.A1(n_2282),
.A2(n_732),
.B1(n_736),
.B2(n_730),
.Y(n_2345)
);

NOR2xp33_ASAP7_75t_SL g2346 ( 
.A(n_2276),
.B(n_1668),
.Y(n_2346)
);

OAI211xp5_ASAP7_75t_SL g2347 ( 
.A1(n_2282),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_2347)
);

AOI211xp5_ASAP7_75t_L g2348 ( 
.A1(n_2282),
.A2(n_751),
.B(n_770),
.C(n_749),
.Y(n_2348)
);

OAI211xp5_ASAP7_75t_L g2349 ( 
.A1(n_2276),
.A2(n_770),
.B(n_39),
.C(n_37),
.Y(n_2349)
);

O2A1O1Ixp33_ASAP7_75t_L g2350 ( 
.A1(n_2276),
.A2(n_1248),
.B(n_41),
.C(n_38),
.Y(n_2350)
);

AOI221x1_ASAP7_75t_L g2351 ( 
.A1(n_2274),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.C(n_44),
.Y(n_2351)
);

AOI211x1_ASAP7_75t_L g2352 ( 
.A1(n_2275),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_2352)
);

AOI211xp5_ASAP7_75t_L g2353 ( 
.A1(n_2282),
.A2(n_1248),
.B(n_49),
.C(n_46),
.Y(n_2353)
);

OAI221xp5_ASAP7_75t_L g2354 ( 
.A1(n_2282),
.A2(n_1668),
.B1(n_2042),
.B2(n_51),
.C(n_48),
.Y(n_2354)
);

NOR2xp67_ASAP7_75t_SL g2355 ( 
.A(n_2276),
.B(n_1185),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2276),
.Y(n_2356)
);

AOI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_2282),
.A2(n_545),
.B(n_543),
.Y(n_2357)
);

OAI22xp5_ASAP7_75t_SL g2358 ( 
.A1(n_2281),
.A2(n_53),
.B1(n_48),
.B2(n_50),
.Y(n_2358)
);

AOI221xp5_ASAP7_75t_L g2359 ( 
.A1(n_2282),
.A2(n_555),
.B1(n_560),
.B2(n_554),
.C(n_553),
.Y(n_2359)
);

AOI211xp5_ASAP7_75t_L g2360 ( 
.A1(n_2282),
.A2(n_59),
.B(n_56),
.C(n_58),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2294),
.B(n_56),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2276),
.Y(n_2362)
);

AOI221xp5_ASAP7_75t_L g2363 ( 
.A1(n_2282),
.A2(n_568),
.B1(n_569),
.B2(n_566),
.C(n_563),
.Y(n_2363)
);

AOI211x1_ASAP7_75t_L g2364 ( 
.A1(n_2275),
.A2(n_62),
.B(n_59),
.C(n_61),
.Y(n_2364)
);

NOR4xp25_ASAP7_75t_L g2365 ( 
.A(n_2282),
.B(n_64),
.C(n_61),
.D(n_62),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_2282),
.B(n_497),
.Y(n_2366)
);

NAND4xp75_ASAP7_75t_L g2367 ( 
.A(n_2251),
.B(n_67),
.C(n_65),
.D(n_66),
.Y(n_2367)
);

AOI21xp5_ASAP7_75t_L g2368 ( 
.A1(n_2282),
.A2(n_572),
.B(n_571),
.Y(n_2368)
);

OAI21xp5_ASAP7_75t_SL g2369 ( 
.A1(n_2282),
.A2(n_66),
.B(n_68),
.Y(n_2369)
);

INVxp67_ASAP7_75t_L g2370 ( 
.A(n_2276),
.Y(n_2370)
);

OR2x2_ASAP7_75t_L g2371 ( 
.A(n_2282),
.B(n_68),
.Y(n_2371)
);

INVxp67_ASAP7_75t_SL g2372 ( 
.A(n_2276),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2276),
.B(n_1967),
.Y(n_2373)
);

AOI21xp5_ASAP7_75t_L g2374 ( 
.A1(n_2282),
.A2(n_577),
.B(n_573),
.Y(n_2374)
);

OAI211xp5_ASAP7_75t_SL g2375 ( 
.A1(n_2282),
.A2(n_73),
.B(n_69),
.C(n_70),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2276),
.B(n_2093),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2276),
.B(n_2093),
.Y(n_2377)
);

OAI211xp5_ASAP7_75t_L g2378 ( 
.A1(n_2276),
.A2(n_76),
.B(n_70),
.C(n_74),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2251),
.Y(n_2379)
);

A2O1A1Ixp33_ASAP7_75t_L g2380 ( 
.A1(n_2282),
.A2(n_865),
.B(n_582),
.C(n_593),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2294),
.B(n_76),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2282),
.A2(n_2030),
.B1(n_2029),
.B2(n_578),
.Y(n_2382)
);

NOR3xp33_ASAP7_75t_L g2383 ( 
.A(n_2276),
.B(n_600),
.C(n_597),
.Y(n_2383)
);

OAI22xp33_ASAP7_75t_L g2384 ( 
.A1(n_2282),
.A2(n_2030),
.B1(n_2029),
.B2(n_1618),
.Y(n_2384)
);

OAI221xp5_ASAP7_75t_SL g2385 ( 
.A1(n_2282),
.A2(n_86),
.B1(n_83),
.B2(n_84),
.C(n_89),
.Y(n_2385)
);

AND2x4_ASAP7_75t_L g2386 ( 
.A(n_2372),
.B(n_89),
.Y(n_2386)
);

OR2x2_ASAP7_75t_L g2387 ( 
.A(n_2296),
.B(n_91),
.Y(n_2387)
);

BUFx2_ASAP7_75t_L g2388 ( 
.A(n_2370),
.Y(n_2388)
);

OR2x2_ASAP7_75t_L g2389 ( 
.A(n_2342),
.B(n_92),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_SL g2390 ( 
.A(n_2356),
.B(n_602),
.Y(n_2390)
);

NOR3xp33_ASAP7_75t_L g2391 ( 
.A(n_2362),
.B(n_611),
.C(n_607),
.Y(n_2391)
);

INVxp67_ASAP7_75t_L g2392 ( 
.A(n_2329),
.Y(n_2392)
);

INVx1_ASAP7_75t_SL g2393 ( 
.A(n_2371),
.Y(n_2393)
);

NOR4xp25_ASAP7_75t_L g2394 ( 
.A(n_2309),
.B(n_95),
.C(n_93),
.D(n_94),
.Y(n_2394)
);

AND2x4_ASAP7_75t_L g2395 ( 
.A(n_2298),
.B(n_93),
.Y(n_2395)
);

NAND4xp25_ASAP7_75t_L g2396 ( 
.A(n_2323),
.B(n_98),
.C(n_94),
.D(n_96),
.Y(n_2396)
);

NAND3xp33_ASAP7_75t_L g2397 ( 
.A(n_2348),
.B(n_1185),
.C(n_634),
.Y(n_2397)
);

OR2x2_ASAP7_75t_L g2398 ( 
.A(n_2361),
.B(n_99),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2381),
.Y(n_2399)
);

NAND4xp75_ASAP7_75t_L g2400 ( 
.A(n_2352),
.B(n_103),
.C(n_100),
.D(n_101),
.Y(n_2400)
);

NOR2xp67_ASAP7_75t_L g2401 ( 
.A(n_2378),
.B(n_101),
.Y(n_2401)
);

NAND4xp75_ASAP7_75t_L g2402 ( 
.A(n_2364),
.B(n_106),
.C(n_104),
.D(n_105),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2320),
.B(n_2063),
.Y(n_2403)
);

INVxp67_ASAP7_75t_SL g2404 ( 
.A(n_2338),
.Y(n_2404)
);

NAND4xp75_ASAP7_75t_L g2405 ( 
.A(n_2305),
.B(n_106),
.C(n_104),
.D(n_105),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2304),
.Y(n_2406)
);

NAND5xp2_ASAP7_75t_L g2407 ( 
.A(n_2327),
.B(n_109),
.C(n_107),
.D(n_108),
.E(n_111),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2304),
.Y(n_2408)
);

AOI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2369),
.A2(n_616),
.B1(n_660),
.B2(n_651),
.Y(n_2409)
);

O2A1O1Ixp33_ASAP7_75t_L g2410 ( 
.A1(n_2380),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_2410)
);

NOR3xp33_ASAP7_75t_L g2411 ( 
.A(n_2379),
.B(n_670),
.C(n_665),
.Y(n_2411)
);

A2O1A1Ixp33_ASAP7_75t_L g2412 ( 
.A1(n_2357),
.A2(n_672),
.B(n_673),
.C(n_671),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2345),
.Y(n_2413)
);

AOI221xp5_ASAP7_75t_L g2414 ( 
.A1(n_2365),
.A2(n_683),
.B1(n_691),
.B2(n_680),
.C(n_675),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2313),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2344),
.B(n_2373),
.Y(n_2416)
);

NAND4xp25_ASAP7_75t_SL g2417 ( 
.A(n_2354),
.B(n_115),
.C(n_113),
.D(n_114),
.Y(n_2417)
);

NOR2x1p5_ASAP7_75t_L g2418 ( 
.A(n_2367),
.B(n_117),
.Y(n_2418)
);

OAI222xp33_ASAP7_75t_L g2419 ( 
.A1(n_2308),
.A2(n_1627),
.B1(n_1655),
.B2(n_1652),
.C1(n_120),
.C2(n_125),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2335),
.B(n_118),
.Y(n_2420)
);

BUFx2_ASAP7_75t_L g2421 ( 
.A(n_2311),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2315),
.Y(n_2422)
);

NOR3x2_ASAP7_75t_L g2423 ( 
.A(n_2295),
.B(n_118),
.C(n_119),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2376),
.B(n_2063),
.Y(n_2424)
);

OAI221xp5_ASAP7_75t_SL g2425 ( 
.A1(n_2334),
.A2(n_127),
.B1(n_124),
.B2(n_126),
.C(n_128),
.Y(n_2425)
);

OAI22xp5_ASAP7_75t_L g2426 ( 
.A1(n_2297),
.A2(n_1185),
.B1(n_1627),
.B2(n_2081),
.Y(n_2426)
);

OAI211xp5_ASAP7_75t_SL g2427 ( 
.A1(n_2366),
.A2(n_129),
.B(n_126),
.C(n_128),
.Y(n_2427)
);

BUFx2_ASAP7_75t_L g2428 ( 
.A(n_2311),
.Y(n_2428)
);

BUFx2_ASAP7_75t_L g2429 ( 
.A(n_2306),
.Y(n_2429)
);

NOR3xp33_ASAP7_75t_L g2430 ( 
.A(n_2337),
.B(n_1065),
.C(n_1123),
.Y(n_2430)
);

OAI22xp5_ASAP7_75t_L g2431 ( 
.A1(n_2382),
.A2(n_1185),
.B1(n_1351),
.B2(n_1349),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2377),
.B(n_130),
.Y(n_2432)
);

NOR2x1_ASAP7_75t_L g2433 ( 
.A(n_2343),
.B(n_131),
.Y(n_2433)
);

OAI21xp5_ASAP7_75t_SL g2434 ( 
.A1(n_2347),
.A2(n_131),
.B(n_132),
.Y(n_2434)
);

INVx1_ASAP7_75t_SL g2435 ( 
.A(n_2358),
.Y(n_2435)
);

OR2x2_ASAP7_75t_L g2436 ( 
.A(n_2299),
.B(n_135),
.Y(n_2436)
);

NOR3xp33_ASAP7_75t_SL g2437 ( 
.A(n_2326),
.B(n_135),
.C(n_137),
.Y(n_2437)
);

AO22x1_ASAP7_75t_L g2438 ( 
.A1(n_2300),
.A2(n_140),
.B1(n_137),
.B2(n_138),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2339),
.B(n_138),
.Y(n_2439)
);

NOR2x1p5_ASAP7_75t_L g2440 ( 
.A(n_2312),
.B(n_140),
.Y(n_2440)
);

OAI21xp33_ASAP7_75t_SL g2441 ( 
.A1(n_2336),
.A2(n_141),
.B(n_142),
.Y(n_2441)
);

NOR2x1_ASAP7_75t_L g2442 ( 
.A(n_2333),
.B(n_141),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2306),
.Y(n_2443)
);

AOI211xp5_ASAP7_75t_L g2444 ( 
.A1(n_2349),
.A2(n_146),
.B(n_143),
.C(n_144),
.Y(n_2444)
);

NOR2x1_ASAP7_75t_L g2445 ( 
.A(n_2375),
.B(n_143),
.Y(n_2445)
);

AND2x4_ASAP7_75t_L g2446 ( 
.A(n_2351),
.B(n_146),
.Y(n_2446)
);

AOI21xp5_ASAP7_75t_L g2447 ( 
.A1(n_2368),
.A2(n_1354),
.B(n_1352),
.Y(n_2447)
);

NOR5xp2_ASAP7_75t_L g2448 ( 
.A(n_2307),
.B(n_149),
.C(n_147),
.D(n_148),
.E(n_150),
.Y(n_2448)
);

INVxp67_ASAP7_75t_L g2449 ( 
.A(n_2302),
.Y(n_2449)
);

XNOR2xp5_ASAP7_75t_L g2450 ( 
.A(n_2360),
.B(n_147),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2331),
.Y(n_2451)
);

OR2x2_ASAP7_75t_L g2452 ( 
.A(n_2328),
.B(n_148),
.Y(n_2452)
);

AND3x4_ASAP7_75t_L g2453 ( 
.A(n_2383),
.B(n_149),
.C(n_151),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2325),
.B(n_2310),
.Y(n_2454)
);

NOR4xp75_ASAP7_75t_L g2455 ( 
.A(n_2321),
.B(n_154),
.C(n_152),
.D(n_153),
.Y(n_2455)
);

XOR2x2_ASAP7_75t_L g2456 ( 
.A(n_2385),
.B(n_153),
.Y(n_2456)
);

NOR2xp33_ASAP7_75t_L g2457 ( 
.A(n_2316),
.B(n_155),
.Y(n_2457)
);

NOR2x1_ASAP7_75t_L g2458 ( 
.A(n_2374),
.B(n_156),
.Y(n_2458)
);

NOR3xp33_ASAP7_75t_L g2459 ( 
.A(n_2359),
.B(n_1126),
.C(n_1124),
.Y(n_2459)
);

NOR2xp67_ASAP7_75t_L g2460 ( 
.A(n_2317),
.B(n_157),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_R g2461 ( 
.A(n_2346),
.B(n_157),
.Y(n_2461)
);

AOI31xp33_ASAP7_75t_SL g2462 ( 
.A1(n_2353),
.A2(n_164),
.A3(n_158),
.B(n_161),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2318),
.B(n_158),
.Y(n_2463)
);

AOI221xp5_ASAP7_75t_L g2464 ( 
.A1(n_2392),
.A2(n_2388),
.B1(n_2415),
.B2(n_2393),
.C(n_2396),
.Y(n_2464)
);

NAND3xp33_ASAP7_75t_L g2465 ( 
.A(n_2421),
.B(n_2330),
.C(n_2324),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_SL g2466 ( 
.A(n_2394),
.B(n_2303),
.Y(n_2466)
);

NAND5xp2_ASAP7_75t_L g2467 ( 
.A(n_2434),
.B(n_2350),
.C(n_2332),
.D(n_2319),
.E(n_2322),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2420),
.A2(n_2404),
.B(n_2390),
.Y(n_2468)
);

NOR2x1_ASAP7_75t_L g2469 ( 
.A(n_2387),
.B(n_2340),
.Y(n_2469)
);

NOR4xp25_ASAP7_75t_L g2470 ( 
.A(n_2435),
.B(n_2363),
.C(n_2355),
.D(n_2384),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_SL g2471 ( 
.A(n_2446),
.B(n_2341),
.Y(n_2471)
);

OAI22xp5_ASAP7_75t_SL g2472 ( 
.A1(n_2453),
.A2(n_2301),
.B1(n_2314),
.B2(n_167),
.Y(n_2472)
);

OAI21xp33_ASAP7_75t_SL g2473 ( 
.A1(n_2417),
.A2(n_165),
.B(n_166),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2446),
.Y(n_2474)
);

NAND4xp25_ASAP7_75t_L g2475 ( 
.A(n_2407),
.B(n_171),
.C(n_165),
.D(n_167),
.Y(n_2475)
);

AOI311xp33_ASAP7_75t_L g2476 ( 
.A1(n_2422),
.A2(n_173),
.A3(n_171),
.B(n_172),
.C(n_175),
.Y(n_2476)
);

NAND3xp33_ASAP7_75t_L g2477 ( 
.A(n_2428),
.B(n_1203),
.C(n_1134),
.Y(n_2477)
);

NAND2x1p5_ASAP7_75t_L g2478 ( 
.A(n_2429),
.B(n_1375),
.Y(n_2478)
);

OAI222xp33_ASAP7_75t_L g2479 ( 
.A1(n_2452),
.A2(n_1652),
.B1(n_1655),
.B2(n_176),
.C1(n_177),
.C2(n_179),
.Y(n_2479)
);

NOR3xp33_ASAP7_75t_L g2480 ( 
.A(n_2449),
.B(n_1134),
.C(n_1132),
.Y(n_2480)
);

NAND3xp33_ASAP7_75t_L g2481 ( 
.A(n_2414),
.B(n_1203),
.C(n_1139),
.Y(n_2481)
);

INVxp67_ASAP7_75t_L g2482 ( 
.A(n_2395),
.Y(n_2482)
);

AOI22xp5_ASAP7_75t_L g2483 ( 
.A1(n_2416),
.A2(n_1357),
.B1(n_1132),
.B2(n_1140),
.Y(n_2483)
);

OAI222xp33_ASAP7_75t_L g2484 ( 
.A1(n_2432),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.C1(n_177),
.C2(n_179),
.Y(n_2484)
);

AOI21xp5_ASAP7_75t_L g2485 ( 
.A1(n_2438),
.A2(n_808),
.B(n_1139),
.Y(n_2485)
);

NAND3xp33_ASAP7_75t_SL g2486 ( 
.A(n_2406),
.B(n_1142),
.C(n_1140),
.Y(n_2486)
);

NAND3xp33_ASAP7_75t_SL g2487 ( 
.A(n_2408),
.B(n_1151),
.C(n_1142),
.Y(n_2487)
);

AOI222xp33_ASAP7_75t_L g2488 ( 
.A1(n_2395),
.A2(n_181),
.B1(n_182),
.B2(n_184),
.C1(n_186),
.C2(n_188),
.Y(n_2488)
);

BUFx3_ASAP7_75t_L g2489 ( 
.A(n_2386),
.Y(n_2489)
);

BUFx2_ASAP7_75t_L g2490 ( 
.A(n_2445),
.Y(n_2490)
);

AOI22xp33_ASAP7_75t_L g2491 ( 
.A1(n_2418),
.A2(n_1203),
.B1(n_497),
.B2(n_1162),
.Y(n_2491)
);

AOI22xp5_ASAP7_75t_L g2492 ( 
.A1(n_2413),
.A2(n_1151),
.B1(n_1172),
.B2(n_1162),
.Y(n_2492)
);

NAND4xp25_ASAP7_75t_L g2493 ( 
.A(n_2457),
.B(n_186),
.C(n_181),
.D(n_182),
.Y(n_2493)
);

NAND4xp25_ASAP7_75t_L g2494 ( 
.A(n_2436),
.B(n_192),
.C(n_189),
.D(n_190),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2440),
.Y(n_2495)
);

NAND4xp25_ASAP7_75t_SL g2496 ( 
.A(n_2444),
.B(n_2441),
.C(n_2410),
.D(n_2433),
.Y(n_2496)
);

AOI211xp5_ASAP7_75t_L g2497 ( 
.A1(n_2425),
.A2(n_193),
.B(n_190),
.C(n_192),
.Y(n_2497)
);

AOI22xp5_ASAP7_75t_L g2498 ( 
.A1(n_2456),
.A2(n_1172),
.B1(n_1179),
.B2(n_1178),
.Y(n_2498)
);

OAI22xp33_ASAP7_75t_SL g2499 ( 
.A1(n_2398),
.A2(n_196),
.B1(n_193),
.B2(n_194),
.Y(n_2499)
);

NOR2x1_ASAP7_75t_L g2500 ( 
.A(n_2389),
.B(n_196),
.Y(n_2500)
);

BUFx2_ASAP7_75t_L g2501 ( 
.A(n_2386),
.Y(n_2501)
);

O2A1O1Ixp33_ASAP7_75t_L g2502 ( 
.A1(n_2412),
.A2(n_201),
.B(n_198),
.C(n_200),
.Y(n_2502)
);

NAND3xp33_ASAP7_75t_SL g2503 ( 
.A(n_2399),
.B(n_1179),
.C(n_1178),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2439),
.Y(n_2504)
);

AOI211xp5_ASAP7_75t_L g2505 ( 
.A1(n_2462),
.A2(n_205),
.B(n_201),
.C(n_204),
.Y(n_2505)
);

AOI22xp5_ASAP7_75t_L g2506 ( 
.A1(n_2450),
.A2(n_1180),
.B1(n_1612),
.B2(n_1321),
.Y(n_2506)
);

INVxp33_ASAP7_75t_L g2507 ( 
.A(n_2458),
.Y(n_2507)
);

NOR4xp25_ASAP7_75t_L g2508 ( 
.A(n_2443),
.B(n_2397),
.C(n_2451),
.D(n_2431),
.Y(n_2508)
);

AOI211xp5_ASAP7_75t_L g2509 ( 
.A1(n_2460),
.A2(n_208),
.B(n_205),
.C(n_207),
.Y(n_2509)
);

NOR4xp25_ASAP7_75t_L g2510 ( 
.A(n_2463),
.B(n_1180),
.C(n_210),
.D(n_208),
.Y(n_2510)
);

XOR2xp5_ASAP7_75t_L g2511 ( 
.A(n_2400),
.B(n_209),
.Y(n_2511)
);

AOI21xp33_ASAP7_75t_L g2512 ( 
.A1(n_2442),
.A2(n_209),
.B(n_210),
.Y(n_2512)
);

OR2x6_ASAP7_75t_L g2513 ( 
.A(n_2401),
.B(n_1095),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2402),
.Y(n_2514)
);

AOI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_2409),
.A2(n_1321),
.B1(n_1515),
.B2(n_1512),
.Y(n_2515)
);

OAI22xp5_ASAP7_75t_L g2516 ( 
.A1(n_2437),
.A2(n_1461),
.B1(n_1472),
.B2(n_1460),
.Y(n_2516)
);

OR2x2_ASAP7_75t_L g2517 ( 
.A(n_2424),
.B(n_211),
.Y(n_2517)
);

AOI22xp33_ASAP7_75t_L g2518 ( 
.A1(n_2427),
.A2(n_497),
.B1(n_1372),
.B2(n_1369),
.Y(n_2518)
);

NAND4xp25_ASAP7_75t_SL g2519 ( 
.A(n_2411),
.B(n_214),
.C(n_211),
.D(n_213),
.Y(n_2519)
);

OAI211xp5_ASAP7_75t_L g2520 ( 
.A1(n_2391),
.A2(n_2461),
.B(n_2447),
.C(n_2454),
.Y(n_2520)
);

NOR2x1_ASAP7_75t_L g2521 ( 
.A(n_2405),
.B(n_213),
.Y(n_2521)
);

NOR2x1p5_ASAP7_75t_L g2522 ( 
.A(n_2423),
.B(n_215),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2455),
.Y(n_2523)
);

INVxp67_ASAP7_75t_L g2524 ( 
.A(n_2403),
.Y(n_2524)
);

NOR3xp33_ASAP7_75t_SL g2525 ( 
.A(n_2419),
.B(n_215),
.C(n_216),
.Y(n_2525)
);

NOR3xp33_ASAP7_75t_L g2526 ( 
.A(n_2430),
.B(n_1059),
.C(n_1053),
.Y(n_2526)
);

NAND3xp33_ASAP7_75t_SL g2527 ( 
.A(n_2448),
.B(n_216),
.C(n_217),
.Y(n_2527)
);

OAI221xp5_ASAP7_75t_L g2528 ( 
.A1(n_2426),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.C(n_225),
.Y(n_2528)
);

NAND3xp33_ASAP7_75t_L g2529 ( 
.A(n_2459),
.B(n_1059),
.C(n_1096),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2501),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2489),
.B(n_224),
.Y(n_2531)
);

AOI21xp5_ASAP7_75t_L g2532 ( 
.A1(n_2471),
.A2(n_1377),
.B(n_1374),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2522),
.Y(n_2533)
);

XNOR2x1_ASAP7_75t_L g2534 ( 
.A(n_2500),
.B(n_226),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2482),
.B(n_226),
.Y(n_2535)
);

AO22x2_ASAP7_75t_L g2536 ( 
.A1(n_2474),
.A2(n_1392),
.B1(n_1395),
.B2(n_1386),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2490),
.Y(n_2537)
);

AOI22xp5_ASAP7_75t_L g2538 ( 
.A1(n_2524),
.A2(n_1321),
.B1(n_1515),
.B2(n_1512),
.Y(n_2538)
);

CKINVDCx20_ASAP7_75t_R g2539 ( 
.A(n_2523),
.Y(n_2539)
);

AND2x4_ASAP7_75t_L g2540 ( 
.A(n_2495),
.B(n_1096),
.Y(n_2540)
);

AOI22x1_ASAP7_75t_SL g2541 ( 
.A1(n_2514),
.A2(n_1400),
.B1(n_1401),
.B2(n_1397),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2513),
.Y(n_2542)
);

AND3x2_ASAP7_75t_L g2543 ( 
.A(n_2509),
.B(n_1407),
.C(n_1402),
.Y(n_2543)
);

NOR3xp33_ASAP7_75t_L g2544 ( 
.A(n_2504),
.B(n_1105),
.C(n_1101),
.Y(n_2544)
);

AOI21xp5_ASAP7_75t_L g2545 ( 
.A1(n_2468),
.A2(n_1105),
.B(n_1101),
.Y(n_2545)
);

NOR3xp33_ASAP7_75t_L g2546 ( 
.A(n_2465),
.B(n_1384),
.C(n_1375),
.Y(n_2546)
);

HB1xp67_ASAP7_75t_L g2547 ( 
.A(n_2517),
.Y(n_2547)
);

XOR2xp5_ASAP7_75t_L g2548 ( 
.A(n_2507),
.B(n_231),
.Y(n_2548)
);

OAI22x1_ASAP7_75t_L g2549 ( 
.A1(n_2511),
.A2(n_1626),
.B1(n_1628),
.B2(n_1611),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2478),
.B(n_2469),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2513),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2505),
.B(n_497),
.Y(n_2552)
);

AOI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2475),
.A2(n_1321),
.B1(n_1553),
.B2(n_1529),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_2499),
.B(n_1072),
.Y(n_2554)
);

AO22x2_ASAP7_75t_L g2555 ( 
.A1(n_2520),
.A2(n_1375),
.B1(n_1398),
.B2(n_1384),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2521),
.B(n_239),
.Y(n_2556)
);

AOI222xp33_ASAP7_75t_L g2557 ( 
.A1(n_2527),
.A2(n_1191),
.B1(n_1072),
.B2(n_1077),
.C1(n_1089),
.C2(n_1097),
.Y(n_2557)
);

AO221x1_ASAP7_75t_L g2558 ( 
.A1(n_2479),
.A2(n_1490),
.B1(n_1497),
.B2(n_1506),
.C(n_1477),
.Y(n_2558)
);

AOI221xp5_ASAP7_75t_L g2559 ( 
.A1(n_2512),
.A2(n_1072),
.B1(n_1074),
.B2(n_1077),
.C(n_1089),
.Y(n_2559)
);

AND2x4_ASAP7_75t_L g2560 ( 
.A(n_2525),
.B(n_240),
.Y(n_2560)
);

HB1xp67_ASAP7_75t_L g2561 ( 
.A(n_2496),
.Y(n_2561)
);

OAI22x1_ASAP7_75t_L g2562 ( 
.A1(n_2519),
.A2(n_1628),
.B1(n_1559),
.B2(n_1558),
.Y(n_2562)
);

OAI211xp5_ASAP7_75t_SL g2563 ( 
.A1(n_2491),
.A2(n_1398),
.B(n_1384),
.C(n_244),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2466),
.Y(n_2564)
);

BUFx3_ASAP7_75t_L g2565 ( 
.A(n_2498),
.Y(n_2565)
);

AOI222xp33_ASAP7_75t_L g2566 ( 
.A1(n_2473),
.A2(n_1191),
.B1(n_1074),
.B2(n_1077),
.C1(n_1089),
.C2(n_1097),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2472),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2494),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2493),
.Y(n_2569)
);

AOI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_2488),
.A2(n_1553),
.B1(n_1529),
.B2(n_1497),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2502),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2516),
.Y(n_2572)
);

A2O1A1Ixp33_ASAP7_75t_L g2573 ( 
.A1(n_2515),
.A2(n_1506),
.B(n_1398),
.C(n_1312),
.Y(n_2573)
);

AND2x4_ASAP7_75t_L g2574 ( 
.A(n_2480),
.B(n_2477),
.Y(n_2574)
);

OAI22x1_ASAP7_75t_L g2575 ( 
.A1(n_2506),
.A2(n_2483),
.B1(n_2492),
.B2(n_2529),
.Y(n_2575)
);

HB1xp67_ASAP7_75t_L g2576 ( 
.A(n_2484),
.Y(n_2576)
);

OAI22xp5_ASAP7_75t_L g2577 ( 
.A1(n_2518),
.A2(n_1557),
.B1(n_1580),
.B2(n_1605),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2497),
.Y(n_2578)
);

INVx3_ASAP7_75t_L g2579 ( 
.A(n_2470),
.Y(n_2579)
);

BUFx3_ASAP7_75t_L g2580 ( 
.A(n_2481),
.Y(n_2580)
);

CKINVDCx20_ASAP7_75t_R g2581 ( 
.A(n_2487),
.Y(n_2581)
);

BUFx2_ASAP7_75t_L g2582 ( 
.A(n_2476),
.Y(n_2582)
);

AOI22xp5_ASAP7_75t_L g2583 ( 
.A1(n_2528),
.A2(n_2508),
.B1(n_2510),
.B2(n_2526),
.Y(n_2583)
);

HB1xp67_ASAP7_75t_L g2584 ( 
.A(n_2485),
.Y(n_2584)
);

AOI22xp5_ASAP7_75t_L g2585 ( 
.A1(n_2486),
.A2(n_1746),
.B1(n_1557),
.B2(n_1556),
.Y(n_2585)
);

XOR2xp5_ASAP7_75t_L g2586 ( 
.A(n_2503),
.B(n_243),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2467),
.Y(n_2587)
);

XNOR2x1_ASAP7_75t_L g2588 ( 
.A(n_2489),
.B(n_246),
.Y(n_2588)
);

AOI221xp5_ASAP7_75t_L g2589 ( 
.A1(n_2464),
.A2(n_1169),
.B1(n_1072),
.B2(n_1074),
.C(n_1077),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2501),
.Y(n_2590)
);

CKINVDCx5p33_ASAP7_75t_R g2591 ( 
.A(n_2501),
.Y(n_2591)
);

INVxp67_ASAP7_75t_SL g2592 ( 
.A(n_2489),
.Y(n_2592)
);

AOI221xp5_ASAP7_75t_L g2593 ( 
.A1(n_2464),
.A2(n_1145),
.B1(n_1074),
.B2(n_1089),
.C(n_1097),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2501),
.Y(n_2594)
);

A2O1A1Ixp33_ASAP7_75t_L g2595 ( 
.A1(n_2464),
.A2(n_1338),
.B(n_1345),
.C(n_1363),
.Y(n_2595)
);

O2A1O1Ixp33_ASAP7_75t_L g2596 ( 
.A1(n_2474),
.A2(n_1338),
.B(n_1345),
.C(n_1356),
.Y(n_2596)
);

INVx2_ASAP7_75t_SL g2597 ( 
.A(n_2591),
.Y(n_2597)
);

INVx2_ASAP7_75t_SL g2598 ( 
.A(n_2530),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2592),
.Y(n_2599)
);

NAND3xp33_ASAP7_75t_L g2600 ( 
.A(n_2590),
.B(n_1103),
.C(n_1097),
.Y(n_2600)
);

OAI221xp5_ASAP7_75t_L g2601 ( 
.A1(n_2594),
.A2(n_2537),
.B1(n_2579),
.B2(n_2561),
.C(n_2582),
.Y(n_2601)
);

NAND5xp2_ASAP7_75t_L g2602 ( 
.A(n_2587),
.B(n_247),
.C(n_249),
.D(n_250),
.E(n_251),
.Y(n_2602)
);

NAND3xp33_ASAP7_75t_L g2603 ( 
.A(n_2547),
.B(n_1110),
.C(n_1103),
.Y(n_2603)
);

XOR2xp5_ASAP7_75t_L g2604 ( 
.A(n_2539),
.B(n_252),
.Y(n_2604)
);

XNOR2xp5_ASAP7_75t_L g2605 ( 
.A(n_2534),
.B(n_253),
.Y(n_2605)
);

AND2x4_ASAP7_75t_L g2606 ( 
.A(n_2533),
.B(n_255),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2550),
.Y(n_2607)
);

OAI22xp5_ASAP7_75t_L g2608 ( 
.A1(n_2564),
.A2(n_1568),
.B1(n_1580),
.B2(n_1605),
.Y(n_2608)
);

AOI22x1_ASAP7_75t_L g2609 ( 
.A1(n_2567),
.A2(n_1103),
.B1(n_1110),
.B2(n_1137),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2560),
.Y(n_2610)
);

AOI22xp33_ASAP7_75t_L g2611 ( 
.A1(n_2560),
.A2(n_1149),
.B1(n_1103),
.B2(n_1110),
.Y(n_2611)
);

AND3x1_ASAP7_75t_L g2612 ( 
.A(n_2556),
.B(n_259),
.C(n_264),
.Y(n_2612)
);

BUFx6f_ASAP7_75t_L g2613 ( 
.A(n_2540),
.Y(n_2613)
);

INVx4_ASAP7_75t_L g2614 ( 
.A(n_2542),
.Y(n_2614)
);

NAND3xp33_ASAP7_75t_SL g2615 ( 
.A(n_2551),
.B(n_1380),
.C(n_1371),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2576),
.Y(n_2616)
);

AOI22xp5_ASAP7_75t_L g2617 ( 
.A1(n_2568),
.A2(n_2569),
.B1(n_2571),
.B2(n_2578),
.Y(n_2617)
);

XNOR2x2_ASAP7_75t_L g2618 ( 
.A(n_2552),
.B(n_266),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2583),
.A2(n_1746),
.B1(n_1191),
.B2(n_1609),
.Y(n_2619)
);

AOI22xp5_ASAP7_75t_L g2620 ( 
.A1(n_2558),
.A2(n_1746),
.B1(n_1191),
.B2(n_1609),
.Y(n_2620)
);

NAND4xp25_ASAP7_75t_L g2621 ( 
.A(n_2557),
.B(n_269),
.C(n_271),
.D(n_273),
.Y(n_2621)
);

OAI222xp33_ASAP7_75t_L g2622 ( 
.A1(n_2553),
.A2(n_1645),
.B1(n_1743),
.B2(n_1731),
.C1(n_1716),
.C2(n_1992),
.Y(n_2622)
);

AOI22xp5_ASAP7_75t_L g2623 ( 
.A1(n_2563),
.A2(n_1746),
.B1(n_1191),
.B2(n_1645),
.Y(n_2623)
);

XNOR2xp5_ASAP7_75t_L g2624 ( 
.A(n_2588),
.B(n_274),
.Y(n_2624)
);

HB1xp67_ASAP7_75t_L g2625 ( 
.A(n_2548),
.Y(n_2625)
);

OAI221xp5_ASAP7_75t_L g2626 ( 
.A1(n_2584),
.A2(n_1155),
.B1(n_1110),
.B2(n_1137),
.C(n_1145),
.Y(n_2626)
);

AOI22xp5_ASAP7_75t_L g2627 ( 
.A1(n_2549),
.A2(n_1568),
.B1(n_1605),
.B2(n_1613),
.Y(n_2627)
);

CKINVDCx20_ASAP7_75t_R g2628 ( 
.A(n_2581),
.Y(n_2628)
);

AOI22xp33_ASAP7_75t_L g2629 ( 
.A1(n_2580),
.A2(n_1155),
.B1(n_1169),
.B2(n_1163),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2531),
.Y(n_2630)
);

OAI222xp33_ASAP7_75t_L g2631 ( 
.A1(n_2541),
.A2(n_1743),
.B1(n_1731),
.B2(n_1549),
.C1(n_1551),
.C2(n_1541),
.Y(n_2631)
);

XOR2xp5_ASAP7_75t_L g2632 ( 
.A(n_2586),
.B(n_277),
.Y(n_2632)
);

AOI221xp5_ASAP7_75t_L g2633 ( 
.A1(n_2559),
.A2(n_1163),
.B1(n_1169),
.B2(n_1161),
.C(n_1155),
.Y(n_2633)
);

NOR2x1p5_ASAP7_75t_L g2634 ( 
.A(n_2535),
.B(n_1137),
.Y(n_2634)
);

NOR3xp33_ASAP7_75t_L g2635 ( 
.A(n_2589),
.B(n_1381),
.C(n_1371),
.Y(n_2635)
);

OAI222xp33_ASAP7_75t_L g2636 ( 
.A1(n_2585),
.A2(n_1743),
.B1(n_1538),
.B2(n_1548),
.C1(n_1546),
.C2(n_1552),
.Y(n_2636)
);

OAI222xp33_ASAP7_75t_L g2637 ( 
.A1(n_2577),
.A2(n_1552),
.B1(n_1548),
.B2(n_1535),
.C1(n_1531),
.C2(n_1526),
.Y(n_2637)
);

NOR2x1p5_ASAP7_75t_L g2638 ( 
.A(n_2565),
.B(n_1137),
.Y(n_2638)
);

NAND3xp33_ASAP7_75t_SL g2639 ( 
.A(n_2566),
.B(n_1381),
.C(n_1356),
.Y(n_2639)
);

NAND3xp33_ASAP7_75t_L g2640 ( 
.A(n_2595),
.B(n_2544),
.C(n_2593),
.Y(n_2640)
);

AO22x2_ASAP7_75t_L g2641 ( 
.A1(n_2554),
.A2(n_2540),
.B1(n_2572),
.B2(n_2574),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2616),
.Y(n_2642)
);

XNOR2xp5_ASAP7_75t_L g2643 ( 
.A(n_2628),
.B(n_2543),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2618),
.Y(n_2644)
);

NOR2xp33_ASAP7_75t_R g2645 ( 
.A(n_2599),
.B(n_2574),
.Y(n_2645)
);

INVx1_ASAP7_75t_SL g2646 ( 
.A(n_2598),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2597),
.Y(n_2647)
);

OAI22xp5_ASAP7_75t_SL g2648 ( 
.A1(n_2601),
.A2(n_2562),
.B1(n_2575),
.B2(n_2570),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2605),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2612),
.Y(n_2650)
);

INVx3_ASAP7_75t_SL g2651 ( 
.A(n_2614),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2624),
.Y(n_2652)
);

AO21x2_ASAP7_75t_L g2653 ( 
.A1(n_2607),
.A2(n_2545),
.B(n_2532),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2625),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2632),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_SL g2656 ( 
.A(n_2610),
.B(n_2617),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2606),
.Y(n_2657)
);

XNOR2xp5_ASAP7_75t_L g2658 ( 
.A(n_2630),
.B(n_2546),
.Y(n_2658)
);

INVx3_ASAP7_75t_SL g2659 ( 
.A(n_2641),
.Y(n_2659)
);

INVx4_ASAP7_75t_L g2660 ( 
.A(n_2613),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2613),
.B(n_2555),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2641),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2604),
.Y(n_2663)
);

INVx2_ASAP7_75t_SL g2664 ( 
.A(n_2634),
.Y(n_2664)
);

OAI21x1_ASAP7_75t_L g2665 ( 
.A1(n_2611),
.A2(n_2596),
.B(n_2538),
.Y(n_2665)
);

AOI21xp33_ASAP7_75t_SL g2666 ( 
.A1(n_2640),
.A2(n_2536),
.B(n_2573),
.Y(n_2666)
);

AOI22xp5_ASAP7_75t_L g2667 ( 
.A1(n_2623),
.A2(n_2536),
.B1(n_1145),
.B2(n_1149),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2620),
.B(n_279),
.Y(n_2668)
);

XNOR2xp5_ASAP7_75t_L g2669 ( 
.A(n_2638),
.B(n_280),
.Y(n_2669)
);

NOR2xp33_ASAP7_75t_R g2670 ( 
.A(n_2615),
.B(n_281),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2609),
.Y(n_2671)
);

HB1xp67_ASAP7_75t_L g2672 ( 
.A(n_2659),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2651),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2642),
.Y(n_2674)
);

AO22x2_ASAP7_75t_L g2675 ( 
.A1(n_2646),
.A2(n_2600),
.B1(n_2603),
.B2(n_2639),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2662),
.Y(n_2676)
);

OAI222xp33_ASAP7_75t_L g2677 ( 
.A1(n_2656),
.A2(n_2608),
.B1(n_2626),
.B2(n_2627),
.C1(n_2629),
.C2(n_2619),
.Y(n_2677)
);

AO22x1_ASAP7_75t_L g2678 ( 
.A1(n_2647),
.A2(n_2635),
.B1(n_2602),
.B2(n_2621),
.Y(n_2678)
);

HB1xp67_ASAP7_75t_L g2679 ( 
.A(n_2654),
.Y(n_2679)
);

OR2x2_ASAP7_75t_L g2680 ( 
.A(n_2660),
.B(n_2631),
.Y(n_2680)
);

OAI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2644),
.A2(n_2633),
.B1(n_2636),
.B2(n_2637),
.Y(n_2681)
);

OAI22xp33_ASAP7_75t_L g2682 ( 
.A1(n_2652),
.A2(n_2622),
.B1(n_1658),
.B2(n_1623),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2657),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2650),
.Y(n_2684)
);

HB1xp67_ASAP7_75t_L g2685 ( 
.A(n_2645),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2643),
.Y(n_2686)
);

OAI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2664),
.A2(n_1155),
.B1(n_1169),
.B2(n_1163),
.Y(n_2687)
);

OAI222xp33_ASAP7_75t_L g2688 ( 
.A1(n_2649),
.A2(n_1068),
.B1(n_1122),
.B2(n_1125),
.C1(n_1135),
.C2(n_1152),
.Y(n_2688)
);

NOR3xp33_ASAP7_75t_L g2689 ( 
.A(n_2655),
.B(n_1404),
.C(n_1393),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2661),
.Y(n_2690)
);

OAI222xp33_ASAP7_75t_L g2691 ( 
.A1(n_2663),
.A2(n_1068),
.B1(n_1122),
.B2(n_1125),
.C1(n_1135),
.C2(n_1152),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2648),
.Y(n_2692)
);

OAI21xp5_ASAP7_75t_L g2693 ( 
.A1(n_2672),
.A2(n_2679),
.B(n_2685),
.Y(n_2693)
);

OAI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2674),
.A2(n_2668),
.B1(n_2669),
.B2(n_2667),
.Y(n_2694)
);

AOI21xp5_ASAP7_75t_L g2695 ( 
.A1(n_2673),
.A2(n_2658),
.B(n_2653),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2676),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2683),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2692),
.B(n_2658),
.Y(n_2698)
);

BUFx2_ASAP7_75t_L g2699 ( 
.A(n_2684),
.Y(n_2699)
);

HB1xp67_ASAP7_75t_L g2700 ( 
.A(n_2686),
.Y(n_2700)
);

OAI22xp5_ASAP7_75t_L g2701 ( 
.A1(n_2690),
.A2(n_2671),
.B1(n_2666),
.B2(n_2670),
.Y(n_2701)
);

INVx3_ASAP7_75t_L g2702 ( 
.A(n_2680),
.Y(n_2702)
);

OAI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2675),
.A2(n_2681),
.B1(n_2682),
.B2(n_2689),
.Y(n_2703)
);

CKINVDCx20_ASAP7_75t_R g2704 ( 
.A(n_2678),
.Y(n_2704)
);

OAI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_2675),
.A2(n_2665),
.B1(n_1145),
.B2(n_1149),
.Y(n_2705)
);

OAI22xp5_ASAP7_75t_L g2706 ( 
.A1(n_2687),
.A2(n_1163),
.B1(n_1149),
.B2(n_1161),
.Y(n_2706)
);

AOI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2700),
.A2(n_2677),
.B1(n_2691),
.B2(n_2688),
.Y(n_2707)
);

OAI22x1_ASAP7_75t_L g2708 ( 
.A1(n_2699),
.A2(n_1404),
.B1(n_1393),
.B2(n_1152),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2693),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2696),
.Y(n_2710)
);

AND2x4_ASAP7_75t_L g2711 ( 
.A(n_2697),
.B(n_282),
.Y(n_2711)
);

OAI22xp5_ASAP7_75t_SL g2712 ( 
.A1(n_2704),
.A2(n_1161),
.B1(n_1406),
.B2(n_1365),
.Y(n_2712)
);

AND3x4_ASAP7_75t_L g2713 ( 
.A(n_2695),
.B(n_283),
.C(n_286),
.Y(n_2713)
);

XNOR2xp5_ASAP7_75t_L g2714 ( 
.A(n_2698),
.B(n_288),
.Y(n_2714)
);

OR2x2_ASAP7_75t_L g2715 ( 
.A(n_2702),
.B(n_289),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2709),
.Y(n_2716)
);

XOR2xp5_ASAP7_75t_L g2717 ( 
.A(n_2710),
.B(n_2701),
.Y(n_2717)
);

NAND2xp33_ASAP7_75t_L g2718 ( 
.A(n_2707),
.B(n_2714),
.Y(n_2718)
);

AOI21xp5_ASAP7_75t_L g2719 ( 
.A1(n_2713),
.A2(n_2694),
.B(n_2703),
.Y(n_2719)
);

HB1xp67_ASAP7_75t_L g2720 ( 
.A(n_2715),
.Y(n_2720)
);

NAND2x1_ASAP7_75t_SL g2721 ( 
.A(n_2711),
.B(n_2705),
.Y(n_2721)
);

AND2x4_ASAP7_75t_L g2722 ( 
.A(n_2716),
.B(n_2720),
.Y(n_2722)
);

BUFx2_ASAP7_75t_L g2723 ( 
.A(n_2717),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2721),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2718),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2723),
.B(n_2719),
.Y(n_2726)
);

OAI21xp5_ASAP7_75t_L g2727 ( 
.A1(n_2722),
.A2(n_2706),
.B(n_2708),
.Y(n_2727)
);

NOR2x1_ASAP7_75t_L g2728 ( 
.A(n_2724),
.B(n_2712),
.Y(n_2728)
);

OR2x6_ASAP7_75t_L g2729 ( 
.A(n_2725),
.B(n_1365),
.Y(n_2729)
);

OAI22xp33_ASAP7_75t_L g2730 ( 
.A1(n_2726),
.A2(n_1406),
.B1(n_1350),
.B2(n_1331),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2728),
.Y(n_2731)
);

OAI21xp5_ASAP7_75t_L g2732 ( 
.A1(n_2727),
.A2(n_1135),
.B(n_1125),
.Y(n_2732)
);

AO21x1_ASAP7_75t_L g2733 ( 
.A1(n_2729),
.A2(n_1135),
.B(n_1125),
.Y(n_2733)
);

AOI221xp5_ASAP7_75t_L g2734 ( 
.A1(n_2731),
.A2(n_1068),
.B1(n_1122),
.B2(n_1318),
.C(n_1301),
.Y(n_2734)
);

OR2x6_ASAP7_75t_L g2735 ( 
.A(n_2733),
.B(n_1263),
.Y(n_2735)
);

OR2x2_ASAP7_75t_L g2736 ( 
.A(n_2732),
.B(n_2730),
.Y(n_2736)
);

AOI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2736),
.A2(n_2735),
.B(n_2734),
.Y(n_2737)
);

AOI211xp5_ASAP7_75t_L g2738 ( 
.A1(n_2737),
.A2(n_293),
.B(n_295),
.C(n_296),
.Y(n_2738)
);


endmodule