module real_jpeg_4856_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_19),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_2),
.B(n_58),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_30),
.B1(n_98),
.B2(n_103),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_2),
.B(n_64),
.C(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_2),
.B(n_134),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_3),
.Y(n_72)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_6),
.A2(n_45),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_7),
.A2(n_38),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_8),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_117),
.Y(n_9)
);

OAI21xp5_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_66),
.B(n_116),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_42),
.B(n_65),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_20),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_18),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_15),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_30),
.B(n_31),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_21),
.A2(n_31),
.B(n_70),
.Y(n_122)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_33),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_22),
.A2(n_68),
.B1(n_69),
.B2(n_77),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_25),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_57),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_57),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_53),
.B(n_56),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_58),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_59),
.A2(n_126),
.B(n_131),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_80),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_80),
.Y(n_116)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_109),
.B1(n_114),
.B2(n_115),
.Y(n_80)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_115),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_97),
.B(n_104),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_105),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B1(n_92),
.B2(n_94),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_SL g127 ( 
.A(n_94),
.Y(n_127)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_143),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_121),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_132),
.B2(n_133),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

AO22x2_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_135),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);


endmodule