module real_jpeg_32233_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_544, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_544;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_469;
wire n_98;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_487;
wire n_93;
wire n_493;
wire n_242;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_0),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_0),
.Y(n_196)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_0),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_0),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_1),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_1),
.Y(n_63)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_1),
.A2(n_63),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22x1_ASAP7_75t_SL g176 ( 
.A1(n_1),
.A2(n_63),
.B1(n_177),
.B2(n_180),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_1),
.A2(n_63),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_2),
.B(n_70),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_2),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_4),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_4),
.Y(n_153)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_5),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_5),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_5),
.Y(n_261)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_5),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_6),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_6),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_6),
.A2(n_119),
.B1(n_273),
.B2(n_369),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_L g435 ( 
.A1(n_6),
.A2(n_212),
.B1(n_273),
.B2(n_436),
.Y(n_435)
);

OAI22xp33_ASAP7_75t_SL g466 ( 
.A1(n_6),
.A2(n_273),
.B1(n_467),
.B2(n_469),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_7),
.A2(n_114),
.B1(n_118),
.B2(n_122),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_7),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_7),
.A2(n_122),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_7),
.A2(n_122),
.B1(n_225),
.B2(n_229),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_7),
.A2(n_122),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_8),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_8),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_8),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_10),
.Y(n_93)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_11),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_11),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_12),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_12),
.A2(n_47),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

AO22x1_ASAP7_75t_SL g201 ( 
.A1(n_12),
.A2(n_47),
.B1(n_202),
.B2(n_205),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_12),
.A2(n_47),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_SL g432 ( 
.A(n_12),
.B(n_177),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_12),
.B(n_170),
.Y(n_462)
);

OAI32xp33_ASAP7_75t_L g480 ( 
.A1(n_12),
.A2(n_427),
.A3(n_481),
.B1(n_486),
.B2(n_492),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_13),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_71),
.B(n_526),
.Y(n_14)
);

INVxp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g526 ( 
.A1(n_16),
.A2(n_527),
.B1(n_541),
.B2(n_542),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_69),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_51),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_18),
.A2(n_185),
.B1(n_188),
.B2(n_544),
.Y(n_184)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_19),
.B(n_188),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_19),
.B(n_52),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_42),
.B(n_43),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_20),
.B(n_43),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_20),
.B(n_270),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_20),
.Y(n_291)
);

NOR2x1p5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.B1(n_28),
.B2(n_31),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_23),
.Y(n_272)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_24),
.Y(n_228)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_24),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_24),
.Y(n_354)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_26),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_27),
.Y(n_351)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_33),
.B(n_270),
.Y(n_327)
);

AO22x2_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_35),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_35),
.Y(n_363)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_37),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_38),
.Y(n_137)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_42),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_42),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_47),
.B(n_48),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_47),
.B(n_56),
.Y(n_400)
);

AOI32xp33_ASAP7_75t_L g426 ( 
.A1(n_47),
.A2(n_427),
.A3(n_429),
.B1(n_431),
.B2(n_432),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_47),
.B(n_487),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_47),
.B(n_81),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_47),
.B(n_195),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_48),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_53),
.B(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_53),
.B(n_303),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_54),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_55),
.B(n_59),
.Y(n_164)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_57),
.A2(n_224),
.B(n_231),
.Y(n_223)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_57),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_58),
.B(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_66),
.Y(n_230)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVxp33_ASAP7_75t_L g541 ( 
.A(n_69),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_304),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_284),
.C(n_302),
.Y(n_72)
);

NOR2xp67_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_245),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_74),
.B(n_537),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_217),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_75),
.B(n_217),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_165),
.C(n_184),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_77),
.B(n_166),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_161),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_112),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_79),
.B(n_162),
.C(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_79),
.A2(n_233),
.B1(n_234),
.B2(n_244),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_79),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_79),
.B(n_298),
.C(n_301),
.Y(n_297)
);

MAJx2_ASAP7_75t_L g376 ( 
.A(n_79),
.B(n_377),
.C(n_378),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_79),
.A2(n_233),
.B1(n_378),
.B2(n_395),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_94),
.B(n_107),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_80),
.B(n_107),
.Y(n_174)
);

NAND2x1p5_ASAP7_75t_L g216 ( 
.A(n_80),
.B(n_176),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_80),
.B(n_209),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_80),
.B(n_435),
.Y(n_447)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_95),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_86),
.B1(n_89),
.B2(n_91),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_88),
.Y(n_199)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_93),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_94),
.B(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_94),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_94),
.B(n_107),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_94),
.B(n_435),
.Y(n_434)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_103),
.B2(n_106),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_99),
.Y(n_439)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_111),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_112),
.Y(n_219)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_123),
.B(n_154),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_114),
.Y(n_347)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_116),
.Y(n_240)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2x1_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_158),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_124),
.B(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_125),
.B(n_238),
.Y(n_266)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_125),
.A2(n_238),
.B(n_294),
.Y(n_293)
);

AO21x2_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_135),
.B(n_140),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_129),
.Y(n_430)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g431 ( 
.A(n_135),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_143),
.B1(n_147),
.B2(n_151),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_154),
.B(n_367),
.Y(n_399)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2x1_ASAP7_75t_L g265 ( 
.A(n_155),
.B(n_266),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_156),
.Y(n_294)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_161),
.A2(n_162),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_161),
.B(n_286),
.C(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_163),
.B(n_327),
.Y(n_377)
);

OAI21x1_ASAP7_75t_SL g290 ( 
.A1(n_164),
.A2(n_224),
.B(n_291),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_164),
.B(n_269),
.Y(n_371)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g277 ( 
.A1(n_167),
.A2(n_168),
.B(n_173),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B(n_171),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_170),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_170),
.B(n_368),
.Y(n_379)
);

NOR2x1_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_172),
.B(n_379),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_174),
.B(n_434),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_175),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_175),
.B(n_252),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_175),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_177),
.B(n_493),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_184),
.B(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_185),
.A2(n_186),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_207),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_187),
.A2(n_188),
.B1(n_426),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2x2_ASAP7_75t_SL g331 ( 
.A(n_188),
.B(n_207),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_188),
.B(n_426),
.Y(n_425)
);

AO21x2_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_193),
.B(n_200),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_193),
.A2(n_316),
.B(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_194),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_194),
.B(n_201),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_194),
.B(n_466),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_195),
.Y(n_503)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_199),
.Y(n_318)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_203),
.Y(n_468)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx4f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_215),
.B(n_216),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_216),
.A2(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_216),
.B(n_313),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_216),
.B(n_434),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_222),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_232),
.Y(n_222)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_224),
.Y(n_299)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_234),
.Y(n_301)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_236),
.B(n_367),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_282),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_246),
.B(n_282),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_277),
.C(n_278),
.Y(n_246)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_247),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_263),
.C(n_267),
.Y(n_247)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_249),
.B(n_330),
.Y(n_329)
);

OAI21x1_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B(n_253),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2x2_ASAP7_75t_SL g384 ( 
.A(n_254),
.B(n_385),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

AND2x4_ASAP7_75t_SL g464 ( 
.A(n_255),
.B(n_465),
.Y(n_464)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_258),
.A2(n_316),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_258),
.B(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_259),
.B(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_261),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_261),
.Y(n_470)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_261),
.Y(n_485)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_261),
.Y(n_491)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_265),
.B(n_268),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_266),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_284),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_285),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_288),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_297),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_292),
.B1(n_295),
.B2(n_296),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_290),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_295),
.C(n_297),
.Y(n_303)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_SL g311 ( 
.A(n_292),
.B(n_312),
.C(n_325),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_293),
.Y(n_388)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_302),
.Y(n_540)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_414),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_336),
.B(n_413),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NOR3xp33_ASAP7_75t_L g415 ( 
.A(n_308),
.B(n_407),
.C(n_416),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_332),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_309),
.B(n_332),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_328),
.C(n_331),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_311),
.B(n_411),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_312),
.B(n_387),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_313),
.B(n_447),
.Y(n_498)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_315),
.B(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_321),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_321),
.B(n_465),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2x1_ASAP7_75t_L g387 ( 
.A(n_326),
.B(n_388),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_329),
.B(n_331),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_389),
.B(n_407),
.C(n_412),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_380),
.Y(n_337)
);

NAND2x1_ASAP7_75t_L g390 ( 
.A(n_338),
.B(n_380),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_372),
.C(n_375),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_339),
.B(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_365),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_371),
.C(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_346),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_342),
.B(n_346),
.Y(n_396)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx4f_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI31xp33_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.A3(n_352),
.B(n_355),
.Y(n_346)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx11_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx12f_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_359),
.B(n_364),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_371),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_366),
.Y(n_382)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_376),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_394),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_378),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_379),
.B(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_384),
.C(n_409),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_390),
.B(n_417),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_405),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_392),
.B(n_405),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_396),
.C(n_397),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_393),
.B(n_441),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_396),
.B(n_398),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.C(n_401),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_399),
.B(n_423),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_400),
.A2(n_401),
.B1(n_402),
.B2(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_400),
.Y(n_424)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_403),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_408),
.B(n_410),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_418),
.Y(n_414)
);

AO21x1_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_442),
.B(n_525),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_440),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_420),
.B(n_440),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_425),
.C(n_433),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_421),
.A2(n_422),
.B1(n_455),
.B2(n_456),
.Y(n_454)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_433),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_426),
.Y(n_453)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx3_ASAP7_75t_SL g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

OAI21x1_ASAP7_75t_SL g442 ( 
.A1(n_443),
.A2(n_457),
.B(n_524),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_454),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_444),
.B(n_454),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_448),
.C(n_451),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_445),
.A2(n_446),
.B1(n_448),
.B2(n_449),
.Y(n_472)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_473),
.B(n_523),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_471),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_SL g523 ( 
.A(n_459),
.B(n_471),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.C(n_463),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_460),
.A2(n_461),
.B1(n_462),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_460),
.Y(n_477)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_464),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_466),
.B(n_503),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_470),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_474),
.A2(n_499),
.B(n_522),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_478),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_475),
.B(n_478),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_498),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_498),
.Y(n_504)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_505),
.B(n_521),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_504),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_501),
.B(n_504),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_511),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_506),
.A2(n_509),
.B(n_520),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_508),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_510),
.B(n_512),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_519),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.Y(n_527)
);

OAI21xp33_ASAP7_75t_L g529 ( 
.A1(n_530),
.A2(n_536),
.B(n_538),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_535),
.Y(n_530)
);

AOI21xp33_ASAP7_75t_L g538 ( 
.A1(n_531),
.A2(n_539),
.B(n_540),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_532),
.A2(n_533),
.B(n_534),
.Y(n_531)
);


endmodule