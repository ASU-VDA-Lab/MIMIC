module fake_jpeg_9049_n_253 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_35),
.Y(n_62)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_29),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_45),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_25),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_25),
.Y(n_47)
);

CKINVDCx9p33_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_58),
.B(n_32),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_25),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_22),
.C(n_38),
.Y(n_91)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_53),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_55),
.B1(n_56),
.B2(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_20),
.B1(n_21),
.B2(n_19),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_20),
.B1(n_19),
.B2(n_21),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_31),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_59),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_17),
.B1(n_34),
.B2(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_0),
.B(n_1),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_69),
.B(n_28),
.C(n_18),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_30),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_33),
.Y(n_98)
);

AO22x1_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_33),
.B1(n_31),
.B2(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_74),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_39),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_72),
.A2(n_58),
.B(n_76),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_22),
.C(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_75),
.Y(n_115)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_81),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_78),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_40),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_93),
.C(n_48),
.Y(n_109)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_91),
.Y(n_116)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_88),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_45),
.B1(n_28),
.B2(n_18),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_86),
.A2(n_94),
.B1(n_96),
.B2(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_27),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_80),
.B(n_83),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_63),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_40),
.C(n_38),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_48),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_40),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_69),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_64),
.A2(n_45),
.B1(n_33),
.B2(n_2),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_51),
.A2(n_44),
.B1(n_38),
.B2(n_40),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_66),
.B1(n_33),
.B2(n_2),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_113),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_64),
.B1(n_50),
.B2(n_44),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_120),
.B1(n_71),
.B2(n_85),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_112),
.C(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_128),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_40),
.C(n_61),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_47),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_47),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_124),
.C(n_3),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_81),
.A2(n_64),
.B1(n_61),
.B2(n_69),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_126),
.B1(n_129),
.B2(n_90),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_66),
.C(n_1),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_125),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_66),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_123),
.A2(n_89),
.B1(n_72),
.B2(n_91),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_132),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_74),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_101),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_139),
.Y(n_160)
);

OAI31xp33_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_72),
.A3(n_103),
.B(n_95),
.Y(n_136)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_153),
.Y(n_168)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_103),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_128),
.C(n_119),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_143),
.A2(n_152),
.B1(n_122),
.B2(n_127),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_88),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_148),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_145),
.B(n_115),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_124),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_116),
.B(n_118),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_101),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_154),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_115),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_105),
.A2(n_90),
.B1(n_95),
.B2(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_99),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_156),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_104),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_176),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_165),
.B(n_179),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_116),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_106),
.C(n_6),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_118),
.B1(n_121),
.B2(n_110),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_170),
.A2(n_152),
.B1(n_138),
.B2(n_135),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_116),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_122),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_16),
.B1(n_7),
.B2(n_10),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_154),
.B1(n_130),
.B2(n_143),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_168),
.B1(n_175),
.B2(n_171),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_179),
.B(n_145),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_191),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_189),
.B1(n_178),
.B2(n_164),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_137),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_197),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_173),
.A2(n_136),
.B1(n_140),
.B2(n_153),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_160),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_169),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_151),
.B(n_147),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_147),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_194),
.C(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_172),
.A2(n_5),
.B(n_6),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_5),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_5),
.B(n_7),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_208),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_194),
.C(n_188),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_205),
.A2(n_211),
.B(n_213),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_161),
.C(n_168),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_212),
.C(n_185),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_186),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_163),
.C(n_165),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_193),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_215),
.C(n_216),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_181),
.C(n_191),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_183),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_223),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_181),
.C(n_189),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_220),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_184),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_188),
.C(n_195),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_224),
.A2(n_201),
.B1(n_162),
.B2(n_11),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_218),
.A2(n_199),
.B1(n_200),
.B2(n_213),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_227),
.A2(n_228),
.B1(n_232),
.B2(n_234),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_225),
.A2(n_207),
.B1(n_200),
.B2(n_167),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_207),
.A3(n_205),
.B1(n_198),
.B2(n_208),
.C1(n_158),
.C2(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_215),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_221),
.A2(n_222),
.B(n_219),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_214),
.B(n_12),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_216),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_235),
.A2(n_239),
.B(n_226),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_231),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g238 ( 
.A(n_232),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_234),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_11),
.C(n_13),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_233),
.C(n_229),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_243),
.C(n_244),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_237),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_237),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_14),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_240),
.C(n_15),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_244),
.B(n_245),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_250),
.C(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_14),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_16),
.Y(n_253)
);


endmodule