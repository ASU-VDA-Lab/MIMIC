module fake_jpeg_20557_n_112 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_112);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx5p33_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_25),
.Y(n_27)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_9),
.Y(n_28)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_17),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_25),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_27),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_44),
.Y(n_48)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_19),
.C(n_21),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_27),
.B(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_51),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_15),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_30),
.B1(n_31),
.B2(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_13),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_63),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_43),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_67),
.C(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_32),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_23),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_48),
.C(n_49),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_77),
.C(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_59),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_37),
.A3(n_40),
.B1(n_39),
.B2(n_42),
.C1(n_26),
.C2(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_64),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_36),
.C(n_20),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_32),
.C(n_42),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_32),
.C(n_59),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_67),
.B1(n_62),
.B2(n_63),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_86),
.B1(n_38),
.B2(n_10),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_88),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_71),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_68),
.C(n_76),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_94),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_22),
.C(n_16),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_96),
.Y(n_99)
);

OAI322xp33_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_10),
.A3(n_9),
.B1(n_13),
.B2(n_14),
.C1(n_18),
.C2(n_25),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_89),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_18),
.C(n_14),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_88),
.B1(n_40),
.B2(n_39),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_93),
.B(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_84),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_37),
.A3(n_26),
.B1(n_3),
.B2(n_4),
.C1(n_1),
.C2(n_6),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_0),
.B(n_1),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_2),
.B(n_4),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_0),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_98),
.B1(n_2),
.B2(n_3),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_108),
.C(n_104),
.Y(n_110)
);

OAI321xp33_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_8),
.C(n_109),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_5),
.Y(n_112)
);


endmodule