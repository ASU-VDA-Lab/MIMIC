module fake_jpeg_7263_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

OR2x2_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_5),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_4),
.B(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_4),
.B(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_0),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_13),
.A2(n_16),
.B1(n_7),
.B2(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_17),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

AND2x6_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_1),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_19),
.A2(n_13),
.B1(n_7),
.B2(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_13),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_15),
.B1(n_18),
.B2(n_14),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_11),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_14),
.C(n_15),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_22),
.C(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_28),
.B1(n_14),
.B2(n_26),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_27),
.B1(n_24),
.B2(n_8),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_32),
.B(n_14),
.Y(n_33)
);

AOI322xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.A3(n_3),
.B1(n_6),
.B2(n_10),
.C1(n_12),
.C2(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_10),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_3),
.B(n_6),
.Y(n_36)
);

BUFx24_ASAP7_75t_SL g37 ( 
.A(n_36),
.Y(n_37)
);


endmodule