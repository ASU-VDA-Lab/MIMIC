module fake_jpeg_11276_n_532 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_532);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_532;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_54),
.B(n_55),
.Y(n_124)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_56),
.Y(n_130)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_69),
.Y(n_141)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_60),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_62),
.B(n_73),
.Y(n_125)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_65),
.Y(n_137)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_38),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_17),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_75),
.B(n_76),
.Y(n_149)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_77),
.B(n_87),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_81),
.B(n_89),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_82),
.Y(n_121)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_19),
.B(n_16),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_22),
.B(n_16),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_93),
.B(n_94),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_27),
.B(n_25),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_27),
.B(n_16),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_95),
.B(n_96),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_99),
.Y(n_112)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_100),
.B(n_101),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_46),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_52),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_105),
.A2(n_106),
.B1(n_110),
.B2(n_111),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_60),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_109),
.B(n_82),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_30),
.B1(n_33),
.B2(n_45),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_30),
.B1(n_33),
.B2(n_45),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_45),
.B1(n_33),
.B2(n_30),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_113),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_57),
.A2(n_23),
.B1(n_30),
.B2(n_33),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_117),
.A2(n_122),
.B1(n_123),
.B2(n_131),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_59),
.A2(n_64),
.B1(n_74),
.B2(n_72),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_63),
.A2(n_45),
.B1(n_43),
.B2(n_34),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_53),
.A2(n_34),
.B1(n_43),
.B2(n_41),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_67),
.A2(n_79),
.B1(n_97),
.B2(n_85),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_65),
.A2(n_50),
.B1(n_29),
.B2(n_44),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_147),
.B1(n_156),
.B2(n_157),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_88),
.A2(n_98),
.B1(n_99),
.B2(n_41),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_70),
.A2(n_37),
.B1(n_25),
.B2(n_36),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_58),
.B(n_42),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_142),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_66),
.B(n_42),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_90),
.A2(n_37),
.B1(n_36),
.B2(n_22),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_92),
.A2(n_29),
.B1(n_50),
.B2(n_47),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_61),
.A2(n_50),
.B1(n_47),
.B2(n_44),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_163),
.Y(n_238)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_164),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_87),
.B(n_29),
.C(n_44),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_165),
.A2(n_187),
.B(n_219),
.Y(n_222)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_166),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_76),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_167),
.B(n_180),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_124),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_172),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_169),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_159),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_173),
.B(n_213),
.Y(n_258)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_178),
.Y(n_256)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_179),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_76),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_103),
.B(n_84),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_211),
.C(n_121),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_125),
.B(n_47),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_193),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_195),
.Y(n_231)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

INVx5_ASAP7_75t_SL g186 ( 
.A(n_152),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_186),
.Y(n_239)
);

NAND2x1_ASAP7_75t_SL g187 ( 
.A(n_116),
.B(n_84),
.Y(n_187)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_188),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_82),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_112),
.Y(n_191)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_147),
.A2(n_135),
.B1(n_112),
.B2(n_127),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_110),
.B(n_111),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_109),
.B(n_0),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_15),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_131),
.A2(n_51),
.B1(n_96),
.B2(n_13),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_137),
.B1(n_158),
.B2(n_128),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_11),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_204),
.Y(n_246)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_200),
.Y(n_269)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_0),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_203),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_143),
.B(n_0),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_130),
.B(n_11),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_161),
.A2(n_51),
.B1(n_2),
.B2(n_3),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_205),
.A2(n_132),
.B1(n_108),
.B2(n_137),
.Y(n_252)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_143),
.B(n_1),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_217),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_130),
.B(n_11),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_208),
.B(n_209),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_108),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_118),
.B(n_2),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_218),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_103),
.B(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_151),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_214),
.B(n_216),
.Y(n_267)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_145),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_215),
.A2(n_199),
.B1(n_188),
.B2(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_104),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_104),
.B(n_3),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_133),
.B(n_3),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_221),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_164),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_226),
.B(n_232),
.C(n_211),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_227),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_181),
.B(n_132),
.Y(n_232)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_182),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_234),
.B(n_259),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_170),
.A2(n_148),
.B1(n_134),
.B2(n_107),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_240),
.A2(n_250),
.B1(n_251),
.B2(n_270),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_R g283 ( 
.A(n_242),
.B(n_211),
.Y(n_283)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_186),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_244),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_194),
.A2(n_108),
.B1(n_132),
.B2(n_134),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_194),
.A2(n_191),
.B1(n_196),
.B2(n_192),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_252),
.A2(n_209),
.B1(n_212),
.B2(n_216),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_182),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_200),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_214),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_174),
.A2(n_158),
.B1(n_114),
.B2(n_120),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_173),
.A2(n_148),
.B1(n_107),
.B2(n_127),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_193),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_271),
.B(n_273),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_165),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_224),
.B(n_183),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_274),
.B(n_275),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_228),
.B(n_207),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_276),
.B(n_289),
.Y(n_357)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_279),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_252),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_221),
.A2(n_171),
.B1(n_217),
.B2(n_203),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_281),
.A2(n_302),
.B1(n_305),
.B2(n_314),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_283),
.B(n_242),
.Y(n_321)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_222),
.A2(n_171),
.B(n_202),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_285),
.A2(n_311),
.B(n_258),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_287),
.B(n_247),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_223),
.A2(n_173),
.B1(n_218),
.B2(n_178),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_288),
.A2(n_308),
.B1(n_270),
.B2(n_220),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_228),
.B(n_163),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_290),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_232),
.B(n_213),
.C(n_206),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_309),
.C(n_316),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_267),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_294),
.Y(n_323)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_293),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_267),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_176),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_297),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_226),
.B(n_201),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_298),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_253),
.B(n_166),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_230),
.B(n_215),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_231),
.B(n_185),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_312),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_240),
.A2(n_177),
.B1(n_169),
.B2(n_162),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_230),
.B(n_119),
.Y(n_304)
);

XNOR2x2_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_310),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_223),
.A2(n_119),
.B1(n_154),
.B2(n_128),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_248),
.Y(n_306)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_225),
.A2(n_120),
.B1(n_114),
.B2(n_154),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_225),
.B(n_179),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_257),
.B(n_235),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_233),
.A2(n_189),
.B(n_121),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_246),
.B(n_4),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_229),
.Y(n_313)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_313),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_235),
.A2(n_96),
.B1(n_5),
.B2(n_6),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_239),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_315),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_258),
.B(n_4),
.C(n_5),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_241),
.B(n_7),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_317),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_307),
.A2(n_239),
.B1(n_241),
.B2(n_243),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_318),
.A2(n_282),
.B1(n_300),
.B2(n_308),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_321),
.B(n_276),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_341),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_329),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_298),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_330),
.B(n_346),
.Y(n_363)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_258),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_334),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_285),
.A2(n_261),
.B1(n_254),
.B2(n_236),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_335),
.A2(n_350),
.B1(n_305),
.B2(n_279),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_337),
.B(n_339),
.C(n_342),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_287),
.B(n_249),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_243),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_340),
.A2(n_345),
.B(n_303),
.Y(n_392)
);

OAI32xp33_ASAP7_75t_L g341 ( 
.A1(n_273),
.A2(n_236),
.A3(n_264),
.B1(n_256),
.B2(n_238),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_283),
.B(n_244),
.Y(n_342)
);

AO22x1_ASAP7_75t_L g345 ( 
.A1(n_299),
.A2(n_264),
.B1(n_256),
.B2(n_262),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_310),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_280),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_347),
.B(n_354),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_299),
.A2(n_266),
.B(n_260),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_349),
.A2(n_300),
.B(n_315),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_281),
.A2(n_261),
.B1(n_254),
.B2(n_237),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_266),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_356),
.C(n_309),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_304),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_296),
.B(n_262),
.C(n_260),
.Y(n_356)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_284),
.Y(n_359)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_359),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_343),
.A2(n_307),
.B1(n_272),
.B2(n_282),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_360),
.A2(n_371),
.B1(n_376),
.B2(n_378),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_364),
.A2(n_349),
.B(n_334),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_340),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_381),
.Y(n_396)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_359),
.Y(n_369)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_369),
.Y(n_398)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_370),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_372),
.B(n_321),
.Y(n_411)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_351),
.Y(n_373)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_336),
.Y(n_374)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_343),
.A2(n_272),
.B1(n_289),
.B2(n_292),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_320),
.A2(n_294),
.B1(n_271),
.B2(n_272),
.Y(n_377)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_357),
.A2(n_277),
.B1(n_288),
.B2(n_293),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_344),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_379),
.B(n_380),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_319),
.B(n_278),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_340),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_348),
.Y(n_382)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_382),
.Y(n_412)
);

OA21x2_ASAP7_75t_L g383 ( 
.A1(n_326),
.A2(n_277),
.B(n_302),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_386),
.Y(n_403)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_387),
.C(n_322),
.Y(n_420)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_332),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_337),
.B(n_316),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_350),
.A2(n_314),
.B1(n_306),
.B2(n_313),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_389),
.A2(n_324),
.B1(n_328),
.B2(n_357),
.Y(n_414)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_391),
.Y(n_405)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_392),
.B(n_345),
.Y(n_409)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_325),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_329),
.A2(n_237),
.B(n_9),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_394),
.A2(n_323),
.B(n_334),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_339),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_395),
.B(n_7),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_397),
.A2(n_364),
.B(n_394),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_401),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_363),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_421),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_408),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_409),
.A2(n_413),
.B(n_374),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_361),
.A2(n_390),
.B1(n_362),
.B2(n_367),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_410),
.A2(n_414),
.B1(n_417),
.B2(n_388),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_411),
.B(n_10),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_366),
.A2(n_355),
.B(n_335),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_333),
.Y(n_415)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_361),
.A2(n_355),
.B1(n_327),
.B2(n_356),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_392),
.B(n_333),
.Y(n_419)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_419),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_422),
.C(n_352),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_376),
.B(n_393),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_375),
.B(n_353),
.C(n_342),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_383),
.A2(n_326),
.B1(n_331),
.B2(n_327),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_423),
.A2(n_362),
.B1(n_366),
.B2(n_388),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_372),
.B(n_358),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_424),
.B(n_322),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_369),
.B(n_352),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_425),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_427),
.A2(n_404),
.B1(n_423),
.B2(n_402),
.Y(n_456)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_428),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_431),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_385),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_442),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_425),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_432),
.A2(n_409),
.B(n_396),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_416),
.A2(n_383),
.B1(n_360),
.B2(n_365),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_434),
.A2(n_436),
.B1(n_441),
.B2(n_404),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_435),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_416),
.A2(n_374),
.B1(n_373),
.B2(n_370),
.Y(n_436)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_439),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_397),
.B(n_384),
.Y(n_440)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_440),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_402),
.A2(n_382),
.B1(n_387),
.B2(n_391),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_395),
.B(n_386),
.C(n_389),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_443),
.B(n_444),
.C(n_408),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_345),
.C(n_9),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_413),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_407),
.B(n_9),
.Y(n_447)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_447),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_406),
.B(n_10),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_448),
.B(n_412),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_449),
.B(n_411),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_10),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_415),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_454),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_432),
.A2(n_451),
.B(n_440),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_463),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_437),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_457),
.B(n_458),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_414),
.Y(n_459)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_459),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_465),
.Y(n_475)
);

INVx13_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_466),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_405),
.Y(n_467)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_470),
.B(n_472),
.Y(n_485)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_471),
.Y(n_487)
);

NOR3xp33_ASAP7_75t_SL g472 ( 
.A(n_433),
.B(n_421),
.C(n_405),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_455),
.A2(n_442),
.B(n_443),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_481),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_453),
.A2(n_454),
.B(n_460),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_480),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_460),
.A2(n_439),
.B(n_440),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_430),
.C(n_441),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_482),
.B(n_484),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_427),
.C(n_446),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_403),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_469),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_464),
.B(n_450),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_488),
.B(n_444),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_463),
.B(n_445),
.C(n_428),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_465),
.C(n_470),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_493),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_487),
.A2(n_461),
.B1(n_471),
.B2(n_452),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_491),
.A2(n_500),
.B1(n_473),
.B2(n_398),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_452),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_492),
.B(n_496),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_485),
.A2(n_434),
.B1(n_467),
.B2(n_459),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_503),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_474),
.B(n_482),
.C(n_489),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_499),
.A2(n_473),
.B(n_480),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_477),
.A2(n_403),
.B1(n_398),
.B2(n_399),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_478),
.B(n_412),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_501),
.B(n_400),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_462),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_502),
.B(n_496),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_476),
.A2(n_472),
.B1(n_466),
.B2(n_419),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_514),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_507),
.B(n_508),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_499),
.B(n_481),
.C(n_486),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_483),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_509),
.B(n_511),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_513),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_497),
.A2(n_486),
.B(n_475),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_497),
.A2(n_399),
.B(n_400),
.Y(n_513)
);

AO21x1_ASAP7_75t_L g515 ( 
.A1(n_505),
.A2(n_493),
.B(n_491),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_515),
.A2(n_508),
.B(n_492),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_506),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_520),
.B(n_521),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_513),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_516),
.C(n_512),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_517),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_524),
.B(n_525),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_519),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_526),
.A2(n_522),
.B1(n_494),
.B2(n_518),
.Y(n_528)
);

OAI321xp33_ASAP7_75t_L g530 ( 
.A1(n_528),
.A2(n_529),
.A3(n_504),
.B1(n_502),
.B2(n_418),
.C(n_449),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_527),
.A2(n_518),
.B1(n_512),
.B2(n_418),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_10),
.Y(n_531)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_531),
.Y(n_532)
);


endmodule