module fake_jpeg_5397_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_5),
.B(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_30),
.B1(n_24),
.B2(n_32),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_22),
.B1(n_28),
.B2(n_25),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_65),
.B(n_23),
.Y(n_93)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_53),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_28),
.B1(n_22),
.B2(n_31),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_68),
.B1(n_47),
.B2(n_23),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_55),
.Y(n_89)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_60),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_28),
.B1(n_20),
.B2(n_31),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_42),
.Y(n_88)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_32),
.B1(n_18),
.B2(n_30),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_66),
.B(n_1),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_35),
.A2(n_32),
.B1(n_18),
.B2(n_34),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_29),
.B1(n_19),
.B2(n_27),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_44),
.B1(n_38),
.B2(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_38),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_76),
.Y(n_105)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_38),
.Y(n_76)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_41),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_96),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_41),
.B1(n_37),
.B2(n_35),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_78),
.A2(n_79),
.B1(n_93),
.B2(n_71),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_81),
.B1(n_56),
.B2(n_66),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_37),
.B1(n_43),
.B2(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_85),
.Y(n_108)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_46),
.B(n_40),
.C(n_27),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_86),
.A2(n_103),
.B(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_91),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_36),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_52),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_64),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_92),
.B(n_97),
.Y(n_117)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

OR2x2_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_12),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_40),
.Y(n_97)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_34),
.B1(n_27),
.B2(n_26),
.Y(n_98)
);

AO21x2_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_27),
.B(n_34),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_49),
.B(n_29),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_55),
.C(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_62),
.B(n_1),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_29),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_107),
.A2(n_114),
.B1(n_118),
.B2(n_127),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_49),
.B1(n_61),
.B2(n_56),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_112),
.B1(n_128),
.B2(n_130),
.Y(n_145)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_61),
.B1(n_66),
.B2(n_60),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_129),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_61),
.B1(n_60),
.B2(n_48),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_116),
.C(n_73),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_71),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_63),
.B1(n_53),
.B2(n_48),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_19),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_100),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_86),
.A2(n_55),
.B1(n_26),
.B2(n_34),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_26),
.B1(n_21),
.B2(n_29),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_84),
.B1(n_82),
.B2(n_75),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_87),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_87),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_67),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_133),
.B(n_92),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_115),
.C(n_126),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_93),
.B(n_88),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_120),
.B(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_144),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_118),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_106),
.Y(n_144)
);

AOI32xp33_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_79),
.A3(n_97),
.B1(n_80),
.B2(n_86),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_159),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_103),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_147),
.B(n_149),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_98),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_156),
.B(n_118),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_96),
.CI(n_104),
.CON(n_149),
.SN(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_104),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_151),
.B(n_152),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_89),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_67),
.B(n_29),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_160),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_89),
.B1(n_87),
.B2(n_26),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_73),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_101),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_85),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_19),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_122),
.A2(n_94),
.B1(n_91),
.B2(n_83),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_164),
.A2(n_165),
.B1(n_114),
.B2(n_118),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_83),
.B1(n_89),
.B2(n_72),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_192),
.C(n_199),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_133),
.B(n_120),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_172),
.A2(n_180),
.B(n_139),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_151),
.B(n_141),
.Y(n_201)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_145),
.A2(n_107),
.B1(n_146),
.B2(n_154),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_189),
.B1(n_193),
.B2(n_195),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_125),
.B(n_113),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_112),
.B1(n_125),
.B2(n_128),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_181),
.A2(n_186),
.B1(n_158),
.B2(n_149),
.Y(n_219)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_185),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_187),
.CI(n_200),
.CON(n_217),
.SN(n_217)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_128),
.B1(n_109),
.B2(n_113),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_128),
.B(n_121),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_128),
.A3(n_130),
.B1(n_121),
.B2(n_131),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_198),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_145),
.A2(n_21),
.B1(n_19),
.B2(n_16),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_134),
.A2(n_21),
.B1(n_15),
.B2(n_14),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_153),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_150),
.B1(n_138),
.B2(n_136),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_134),
.A2(n_135),
.B(n_160),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_149),
.B(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_15),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_159),
.B(n_14),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_201),
.B(n_205),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_208),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_184),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_204),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_169),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_144),
.B(n_148),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_218),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_169),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_223),
.B1(n_212),
.B2(n_222),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_222),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_219),
.A2(n_221),
.B1(n_224),
.B2(n_229),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_183),
.A2(n_175),
.B(n_194),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_176),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_181),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_227),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_167),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_225),
.A2(n_228),
.B1(n_173),
.B2(n_182),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_166),
.B(n_13),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_199),
.C(n_200),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_167),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_233),
.A2(n_253),
.B1(n_221),
.B2(n_229),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_166),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_192),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_243),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_247),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_190),
.B1(n_185),
.B2(n_174),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_249),
.A2(n_252),
.B1(n_254),
.B2(n_213),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_204),
.B(n_174),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_173),
.B1(n_170),
.B2(n_171),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_225),
.A2(n_168),
.B1(n_7),
.B2(n_8),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_219),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_238),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_256),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_232),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_257),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_220),
.C(n_201),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_260),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_231),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_207),
.C(n_206),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_266),
.C(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_251),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_255),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_240),
.C(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_271),
.B(n_210),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_205),
.C(n_208),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_202),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_276),
.C(n_252),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_210),
.C(n_217),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_272),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_279),
.A2(n_228),
.B(n_224),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_248),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_287),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_271),
.B(n_258),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_235),
.CI(n_248),
.CON(n_283),
.SN(n_283)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_283),
.B(n_285),
.Y(n_302)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_236),
.B1(n_230),
.B2(n_212),
.Y(n_286)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_253),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_255),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_261),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_244),
.C(n_217),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_261),
.C(n_276),
.Y(n_300)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_298),
.B(n_306),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_264),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_296),
.B(n_304),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_269),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_301),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_288),
.Y(n_304)
);

AOI32xp33_ASAP7_75t_L g305 ( 
.A1(n_280),
.A2(n_273),
.A3(n_267),
.B1(n_244),
.B2(n_259),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_282),
.B(n_279),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_273),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_282),
.C(n_291),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_303),
.A2(n_284),
.B1(n_277),
.B2(n_283),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_309),
.A2(n_310),
.B(n_315),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_277),
.B(n_283),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_316),
.C(n_318),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_302),
.A2(n_293),
.B1(n_292),
.B2(n_291),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_317),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_295),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_217),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_9),
.C(n_10),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_299),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_320),
.A2(n_324),
.B(n_326),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_328),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_307),
.B1(n_301),
.B2(n_300),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_319),
.C(n_10),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_9),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_9),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_10),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_322),
.B(n_314),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_329),
.A2(n_332),
.B(n_334),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_325),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_313),
.Y(n_333)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_333),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_321),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_327),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_337),
.B(n_331),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_335),
.B1(n_319),
.B2(n_13),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_11),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_11),
.B(n_12),
.Y(n_342)
);


endmodule