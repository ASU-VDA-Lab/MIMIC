module fake_jpeg_13161_n_574 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_574);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_574;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_9),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_54),
.B(n_67),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_60),
.Y(n_155)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_46),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_53),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_69),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_33),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_76),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_21),
.B(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_10),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_79),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_94),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_22),
.B(n_8),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_22),
.B(n_8),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_98),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_28),
.B(n_11),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_28),
.B(n_7),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_36),
.B(n_12),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_59),
.A2(n_27),
.B1(n_35),
.B2(n_29),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_122),
.A2(n_148),
.B1(n_80),
.B2(n_62),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_75),
.A2(n_52),
.B1(n_42),
.B2(n_29),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_128),
.A2(n_135),
.B1(n_154),
.B2(n_91),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g134 ( 
.A1(n_69),
.A2(n_36),
.B(n_43),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_49),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_73),
.A2(n_29),
.B1(n_52),
.B2(n_43),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_81),
.A2(n_35),
.B1(n_25),
.B2(n_34),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_152),
.B1(n_168),
.B2(n_104),
.Y(n_176)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_66),
.A2(n_27),
.B1(n_35),
.B2(n_52),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_105),
.A2(n_34),
.B1(n_44),
.B2(n_30),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_57),
.A2(n_34),
.B1(n_26),
.B2(n_30),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_55),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_64),
.A2(n_34),
.B1(n_44),
.B2(n_40),
.Y(n_168)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_56),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_82),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_174),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_51),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_175),
.B(n_182),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_176),
.A2(n_183),
.B1(n_202),
.B2(n_226),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_178),
.B(n_196),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_112),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_179),
.B(n_211),
.Y(n_255)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_181),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_132),
.B(n_69),
.CI(n_90),
.CON(n_182),
.SN(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_168),
.A2(n_70),
.B1(n_77),
.B2(n_86),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_114),
.B(n_40),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_187),
.Y(n_263)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_188),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_117),
.B(n_58),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_191),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_192),
.B(n_224),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_193),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_194),
.Y(n_271)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_195),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_140),
.B(n_39),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_198),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_119),
.B(n_51),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_0),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_116),
.B(n_14),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_200),
.B(n_223),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_201),
.A2(n_220),
.B1(n_231),
.B2(n_235),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_152),
.A2(n_102),
.B1(n_65),
.B2(n_60),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_203),
.Y(n_251)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_133),
.Y(n_204)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_207),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_164),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_146),
.B(n_93),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_118),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_137),
.Y(n_212)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_213),
.Y(n_281)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

INVx3_ASAP7_75t_SL g292 ( 
.A(n_214),
.Y(n_292)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_153),
.B(n_68),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_138),
.C(n_167),
.Y(n_237)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_219),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_143),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_154),
.A2(n_101),
.B1(n_72),
.B2(n_48),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_222),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_109),
.B(n_15),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_111),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_142),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_228),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_122),
.A2(n_48),
.B1(n_45),
.B2(n_49),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_111),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_227),
.Y(n_290)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_115),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_125),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_157),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_233),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_144),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_141),
.B(n_49),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_170),
.B(n_15),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_113),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_32),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_138),
.A2(n_49),
.B1(n_32),
.B2(n_24),
.Y(n_235)
);

AO22x2_ASAP7_75t_L g236 ( 
.A1(n_157),
.A2(n_103),
.B1(n_48),
.B2(n_45),
.Y(n_236)
);

AOI22x1_ASAP7_75t_L g275 ( 
.A1(n_236),
.A2(n_160),
.B1(n_149),
.B2(n_144),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_237),
.B(n_254),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_148),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_241),
.A2(n_254),
.B(n_235),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_201),
.A2(n_123),
.B(n_167),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_242),
.A2(n_275),
.B(n_177),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_246),
.B(n_278),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_113),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_249),
.B(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_182),
.B(n_130),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_172),
.B(n_159),
.C(n_103),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_184),
.B(n_150),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_267),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_180),
.B(n_150),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_183),
.A2(n_136),
.B1(n_120),
.B2(n_149),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_269),
.A2(n_273),
.B1(n_276),
.B2(n_277),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_192),
.A2(n_136),
.B1(n_120),
.B2(n_162),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_191),
.A2(n_160),
.B1(n_162),
.B2(n_48),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_191),
.A2(n_48),
.B1(n_49),
.B2(n_32),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_188),
.B(n_0),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_0),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_217),
.A2(n_32),
.B1(n_6),
.B2(n_12),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_284),
.A2(n_257),
.B(n_248),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_174),
.B1(n_214),
.B2(n_181),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_294),
.A2(n_334),
.B1(n_336),
.B2(n_339),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_251),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_303),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_297),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_189),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_298),
.B(n_320),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_272),
.Y(n_351)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_301),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_307),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_267),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_304),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_174),
.C(n_190),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_305),
.B(n_319),
.C(n_5),
.Y(n_387)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_306),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_258),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_279),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_312),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_260),
.A2(n_257),
.B1(n_248),
.B2(n_243),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_310),
.A2(n_314),
.B1(n_292),
.B2(n_283),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_241),
.A2(n_236),
.B1(n_219),
.B2(n_230),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_311),
.A2(n_315),
.B1(n_327),
.B2(n_332),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_246),
.B(n_195),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_238),
.Y(n_313)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_313),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_260),
.A2(n_177),
.B1(n_187),
.B2(n_209),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_241),
.A2(n_236),
.B1(n_218),
.B2(n_231),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_249),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_316),
.B(n_321),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_240),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_317),
.A2(n_326),
.B(n_13),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_263),
.Y(n_318)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_268),
.B(n_185),
.C(n_203),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_227),
.C(n_17),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_238),
.Y(n_322)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_322),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_274),
.B(n_236),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_325),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_204),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_261),
.A2(n_273),
.B1(n_247),
.B2(n_285),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_264),
.Y(n_329)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_329),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_268),
.B(n_215),
.C(n_206),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_290),
.C(n_256),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_287),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_261),
.A2(n_220),
.B1(n_228),
.B2(n_224),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_333),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_285),
.A2(n_216),
.B1(n_209),
.B2(n_193),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_266),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_335),
.B(n_338),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_285),
.A2(n_247),
.B1(n_286),
.B2(n_275),
.Y(n_336)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_287),
.Y(n_337)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_243),
.B(n_290),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_239),
.B(n_216),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_340),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_239),
.B(n_198),
.Y(n_341)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_270),
.C(n_259),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_244),
.A2(n_242),
.B1(n_275),
.B2(n_284),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_342),
.A2(n_263),
.B1(n_271),
.B2(n_289),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_291),
.A2(n_198),
.B1(n_194),
.B2(n_3),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_343),
.A2(n_292),
.B1(n_294),
.B2(n_326),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_296),
.A2(n_280),
.B(n_272),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_347),
.A2(n_373),
.B(n_383),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_352),
.C(n_355),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_293),
.B(n_250),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_353),
.A2(n_364),
.B1(n_366),
.B2(n_368),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_296),
.B(n_291),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_358),
.A2(n_372),
.B1(n_379),
.B2(n_6),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_370),
.C(n_330),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_336),
.A2(n_289),
.B1(n_282),
.B2(n_265),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_297),
.A2(n_271),
.B(n_283),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_SL g398 ( 
.A1(n_365),
.A2(n_311),
.B(n_327),
.C(n_323),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_316),
.A2(n_256),
.B1(n_282),
.B2(n_265),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_324),
.A2(n_270),
.B1(n_259),
.B2(n_292),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_299),
.B(n_250),
.C(n_252),
.Y(n_370)
);

MAJx2_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_370),
.C(n_320),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_338),
.A2(n_252),
.B(n_245),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_342),
.A2(n_194),
.B1(n_245),
.B2(n_3),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_301),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_382),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_303),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_385),
.A2(n_305),
.B(n_325),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_309),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_343),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_13),
.Y(n_421)
);

MAJx2_ASAP7_75t_L g433 ( 
.A(n_389),
.B(n_369),
.C(n_377),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_328),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_390),
.B(n_416),
.Y(n_451)
);

OA22x2_ASAP7_75t_L g392 ( 
.A1(n_346),
.A2(n_307),
.B1(n_334),
.B2(n_315),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_392),
.B(n_409),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_346),
.A2(n_378),
.B1(n_350),
.B2(n_345),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_394),
.A2(n_396),
.B1(n_382),
.B2(n_384),
.Y(n_434)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_349),
.Y(n_395)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_395),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_378),
.A2(n_350),
.B1(n_357),
.B2(n_358),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_360),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_397),
.A2(n_405),
.B1(n_415),
.B2(n_420),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_398),
.A2(n_401),
.B(n_403),
.Y(n_436)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_399),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_332),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_400),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_404),
.C(n_413),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_365),
.A2(n_300),
.B(n_319),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_351),
.B(n_300),
.Y(n_404)
);

AO21x1_ASAP7_75t_L g405 ( 
.A1(n_347),
.A2(n_312),
.B(n_340),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_344),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g427 ( 
.A(n_406),
.Y(n_427)
);

AO22x1_ASAP7_75t_L g407 ( 
.A1(n_373),
.A2(n_306),
.B1(n_304),
.B2(n_335),
.Y(n_407)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_407),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_408),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_366),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_410),
.B(n_412),
.Y(n_456)
);

OAI211xp5_ASAP7_75t_L g411 ( 
.A1(n_374),
.A2(n_302),
.B(n_333),
.C(n_329),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_386),
.Y(n_428)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_380),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_352),
.B(n_322),
.C(n_313),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_354),
.B(n_295),
.Y(n_414)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_414),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_353),
.A2(n_318),
.B1(n_337),
.B2(n_331),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_354),
.B(n_308),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_355),
.B(n_5),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_419),
.C(n_421),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_357),
.B(n_6),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_363),
.B(n_13),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_362),
.B(n_387),
.C(n_371),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_422),
.B(n_424),
.Y(n_437)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_380),
.Y(n_423)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_423),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_364),
.B(n_13),
.C(n_16),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_368),
.A2(n_17),
.B1(n_18),
.B2(n_385),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_425),
.A2(n_348),
.B1(n_376),
.B2(n_361),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_428),
.B(n_393),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_L g475 ( 
.A(n_433),
.B(n_458),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_434),
.A2(n_440),
.B1(n_442),
.B2(n_444),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_435),
.A2(n_409),
.B1(n_407),
.B2(n_415),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_396),
.A2(n_384),
.B1(n_356),
.B2(n_367),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_394),
.A2(n_356),
.B1(n_367),
.B2(n_348),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_388),
.A2(n_375),
.B1(n_381),
.B2(n_17),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_443),
.A2(n_450),
.B1(n_424),
.B2(n_393),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_400),
.A2(n_375),
.B1(n_17),
.B2(n_18),
.Y(n_444)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_414),
.Y(n_447)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_397),
.Y(n_448)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_448),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_388),
.A2(n_18),
.B1(n_401),
.B2(n_405),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_452),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_407),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_392),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_400),
.A2(n_408),
.B1(n_398),
.B2(n_392),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_455),
.A2(n_398),
.B1(n_425),
.B2(n_392),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_391),
.B(n_402),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_457),
.B(n_422),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_391),
.B(n_404),
.Y(n_458)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_459),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_461),
.B(n_463),
.C(n_465),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_469),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_457),
.B(n_413),
.C(n_389),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_403),
.C(n_398),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_467),
.B(n_426),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_427),
.B(n_419),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_468),
.B(n_479),
.Y(n_507)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_441),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_441),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_471),
.Y(n_488)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_447),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_472),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_473),
.A2(n_480),
.B1(n_443),
.B2(n_435),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_474),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_432),
.B(n_417),
.C(n_421),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_476),
.B(n_482),
.C(n_453),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_436),
.A2(n_423),
.B(n_412),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_477),
.B(n_481),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_448),
.B(n_451),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_478),
.B(n_484),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_430),
.B(n_439),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_450),
.A2(n_449),
.B1(n_426),
.B2(n_429),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_456),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_437),
.C(n_433),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_428),
.B(n_431),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_436),
.A2(n_455),
.B(n_449),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_485),
.A2(n_467),
.B(n_480),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_434),
.B(n_437),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_486),
.B(n_444),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_490),
.A2(n_485),
.B(n_473),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_494),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_465),
.B(n_440),
.Y(n_494)
);

INVx5_ASAP7_75t_L g496 ( 
.A(n_478),
.Y(n_496)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_496),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_475),
.B(n_439),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_497),
.B(n_498),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_475),
.B(n_453),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_442),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_500),
.B(n_509),
.C(n_483),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_504),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_502),
.A2(n_459),
.B1(n_462),
.B2(n_460),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_430),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_463),
.B(n_452),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_506),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_481),
.B(n_445),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_508),
.B(n_468),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_476),
.B(n_477),
.C(n_469),
.Y(n_509)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_511),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_512),
.A2(n_499),
.B(n_492),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_514),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_489),
.A2(n_479),
.B(n_464),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_515),
.A2(n_525),
.B(n_492),
.Y(n_531)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_488),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_519),
.Y(n_537)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_487),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_496),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_523),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_521),
.B(n_494),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_493),
.B(n_464),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_522),
.B(n_526),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_505),
.B(n_460),
.C(n_470),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_502),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_524),
.B(n_527),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_490),
.A2(n_471),
.B(n_466),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_504),
.B(n_483),
.C(n_466),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_507),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_521),
.B(n_509),
.C(n_495),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_529),
.B(n_533),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_524),
.A2(n_499),
.B1(n_503),
.B2(n_438),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_530),
.A2(n_514),
.B1(n_516),
.B2(n_520),
.Y(n_546)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_531),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_535),
.B(n_510),
.C(n_516),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_525),
.A2(n_491),
.B(n_500),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_541),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_512),
.A2(n_497),
.B(n_495),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_539),
.B(n_528),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_501),
.C(n_498),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_438),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_543),
.B(n_523),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_537),
.B(n_513),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_544),
.B(n_547),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_546),
.A2(n_550),
.B1(n_531),
.B2(n_536),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_534),
.B(n_519),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_549),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_532),
.B(n_517),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_552),
.B(n_553),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g554 ( 
.A(n_541),
.B(n_528),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_554),
.B(n_539),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_545),
.B(n_529),
.C(n_535),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_557),
.A2(n_560),
.B(n_549),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_550),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_559),
.B(n_561),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_557),
.A2(n_548),
.B(n_551),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_563),
.A2(n_564),
.B(n_565),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_556),
.B(n_538),
.C(n_542),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_562),
.B(n_558),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_566),
.B(n_568),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_555),
.C(n_540),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_R g569 ( 
.A(n_567),
.B(n_555),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_569),
.A2(n_533),
.B(n_518),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_571),
.A2(n_570),
.B(n_446),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_R g573 ( 
.A(n_572),
.B(n_515),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_573),
.A2(n_510),
.B(n_530),
.Y(n_574)
);


endmodule