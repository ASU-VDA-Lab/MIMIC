module fake_ariane_1074_n_996 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_996);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_996;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_731;
wire n_336;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_840;
wire n_426;
wire n_433;
wire n_600;
wire n_481;
wire n_721;
wire n_795;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_839;
wire n_821;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_677;
wire n_614;
wire n_604;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_988;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_699;
wire n_727;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_715;
wire n_512;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_658;
wire n_616;
wire n_705;
wire n_630;
wire n_617;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_741;
wire n_747;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_680;
wire n_571;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_76),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_125),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_104),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_39),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_153),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_163),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_157),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_4),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_0),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_93),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_106),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_73),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_152),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_150),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_94),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_166),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_13),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_53),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_84),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_161),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_54),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_95),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_17),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_137),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_174),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_115),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_60),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_116),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_63),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_197),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_136),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_75),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_192),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_17),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_147),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_196),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_180),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_44),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_4),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_118),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_24),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_67),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_46),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_131),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_112),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_77),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_88),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_160),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_162),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_37),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_34),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_35),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_188),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_117),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_24),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_83),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_176),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_109),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_144),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_64),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_199),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_191),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_151),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_74),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_35),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_56),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_145),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_127),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_156),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_101),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_31),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_23),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_178),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_179),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_78),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_66),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_69),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_211),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_224),
.Y(n_287)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_215),
.B(n_283),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_207),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_0),
.Y(n_291)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_215),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_207),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_1),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_1),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_217),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_2),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_218),
.B(n_40),
.Y(n_299)
);

BUFx12f_ASAP7_75t_L g300 ( 
.A(n_263),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_2),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_202),
.B(n_3),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_260),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_215),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g306 ( 
.A(n_212),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_283),
.Y(n_307)
);

BUFx12f_ASAP7_75t_L g308 ( 
.A(n_205),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_283),
.Y(n_309)
);

CKINVDCx6p67_ASAP7_75t_R g310 ( 
.A(n_225),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_217),
.B(n_3),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_208),
.B(n_5),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_213),
.B(n_5),
.Y(n_313)
);

NOR2x1_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_41),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_214),
.B(n_6),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_6),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_216),
.Y(n_317)
);

AND2x6_ASAP7_75t_L g318 ( 
.A(n_220),
.B(n_42),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_7),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_222),
.Y(n_320)
);

BUFx12f_ASAP7_75t_L g321 ( 
.A(n_205),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_229),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_241),
.B(n_7),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_231),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_247),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_235),
.B(n_8),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_239),
.B(n_8),
.Y(n_327)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_221),
.Y(n_328)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_221),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_242),
.B(n_43),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_248),
.B(n_9),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_227),
.B(n_9),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_249),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_258),
.B(n_10),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

BUFx12f_ASAP7_75t_L g336 ( 
.A(n_206),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_252),
.B(n_10),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_253),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_286),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_L g340 ( 
.A1(n_299),
.A2(n_278),
.B1(n_225),
.B2(n_259),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_227),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_287),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_293),
.B(n_273),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_310),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_308),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_206),
.Y(n_346)
);

AO22x2_ASAP7_75t_L g347 ( 
.A1(n_334),
.A2(n_267),
.B1(n_254),
.B2(n_257),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_332),
.A2(n_278),
.B1(n_236),
.B2(n_281),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_334),
.A2(n_264),
.B1(n_265),
.B2(n_268),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_333),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_L g351 ( 
.A1(n_300),
.A2(n_209),
.B1(n_282),
.B2(n_281),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_L g352 ( 
.A1(n_300),
.A2(n_209),
.B1(n_282),
.B2(n_269),
.Y(n_352)
);

INVx8_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_291),
.A2(n_285),
.B1(n_276),
.B2(n_275),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_291),
.A2(n_274),
.B1(n_272),
.B2(n_271),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_L g357 ( 
.A1(n_323),
.A2(n_270),
.B1(n_266),
.B2(n_261),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_296),
.A2(n_233),
.B1(n_255),
.B2(n_251),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_200),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_294),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_296),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_303),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_295),
.B(n_11),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_210),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_298),
.A2(n_237),
.B1(n_245),
.B2(n_244),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_304),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_298),
.A2(n_232),
.B1(n_243),
.B2(n_240),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_304),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_295),
.A2(n_219),
.B1(n_223),
.B2(n_226),
.Y(n_369)
);

AND2x2_ASAP7_75t_SL g370 ( 
.A(n_311),
.B(n_316),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_301),
.A2(n_238),
.B1(n_234),
.B2(n_228),
.Y(n_371)
);

AO22x2_ASAP7_75t_L g372 ( 
.A1(n_311),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_290),
.B(n_256),
.Y(n_373)
);

AOI22x1_ASAP7_75t_L g374 ( 
.A1(n_316),
.A2(n_256),
.B1(n_14),
.B2(n_15),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_290),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_302),
.A2(n_256),
.B1(n_14),
.B2(n_15),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_302),
.A2(n_256),
.B1(n_16),
.B2(n_18),
.Y(n_378)
);

OR2x6_ASAP7_75t_L g379 ( 
.A(n_321),
.B(n_12),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_L g380 ( 
.A1(n_321),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_328),
.B(n_256),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_297),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_328),
.B(n_256),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_304),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_305),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_336),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_L g388 ( 
.A1(n_336),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_388)
);

INVxp33_ASAP7_75t_L g389 ( 
.A(n_297),
.Y(n_389)
);

AO22x2_ASAP7_75t_L g390 ( 
.A1(n_319),
.A2(n_317),
.B1(n_337),
.B2(n_315),
.Y(n_390)
);

AO22x2_ASAP7_75t_L g391 ( 
.A1(n_319),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_320),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_328),
.B(n_256),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_317),
.B(n_22),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_376),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_342),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_350),
.B(n_329),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_353),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_373),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_382),
.B(n_329),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_383),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_389),
.Y(n_405)
);

BUFx5_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_394),
.Y(n_407)
);

NAND2x1p5_ASAP7_75t_L g408 ( 
.A(n_341),
.B(n_314),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_343),
.Y(n_409)
);

OR2x6_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_312),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_346),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_359),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_354),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_366),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_368),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_348),
.B(n_320),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_329),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_390),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_386),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_369),
.B(n_320),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_386),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_386),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_364),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_363),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_371),
.B(n_329),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_371),
.B(n_322),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_349),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_356),
.B(n_322),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_381),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_384),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_377),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_345),
.B(n_322),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_375),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_377),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_340),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_378),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_356),
.B(n_322),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_378),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_347),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_372),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_391),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_391),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_355),
.B(n_335),
.Y(n_447)
);

INVx3_ASAP7_75t_R g448 ( 
.A(n_344),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_387),
.B(n_361),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_358),
.B(n_335),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_379),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_358),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_365),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_353),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_365),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_367),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_L g457 ( 
.A(n_367),
.B(n_289),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_379),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_353),
.B(n_335),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_379),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_357),
.Y(n_461)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_351),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_380),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_352),
.B(n_327),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_382),
.B(n_335),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_340),
.B(n_318),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_370),
.B(n_338),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_462),
.B(n_313),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_418),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_468),
.B(n_313),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_402),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_468),
.B(n_318),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_405),
.B(n_326),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_405),
.B(n_416),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_396),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_411),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_439),
.B(n_452),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_326),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_418),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_419),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_454),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_459),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_428),
.B(n_331),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_406),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_431),
.A2(n_330),
.B(n_318),
.Y(n_488)
);

BUFx12f_ASAP7_75t_SL g489 ( 
.A(n_410),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_428),
.B(n_331),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_430),
.B(n_318),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_404),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_401),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_398),
.Y(n_494)
);

AND2x2_ASAP7_75t_SL g495 ( 
.A(n_467),
.B(n_318),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_430),
.B(n_330),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_445),
.B(n_330),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_406),
.Y(n_500)
);

BUFx4f_ASAP7_75t_L g501 ( 
.A(n_408),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_406),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_456),
.B(n_338),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_462),
.B(n_338),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_444),
.B(n_330),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_421),
.B(n_338),
.Y(n_508)
);

AND2x4_ASAP7_75t_SL g509 ( 
.A(n_454),
.B(n_330),
.Y(n_509)
);

NAND2x1p5_ASAP7_75t_L g510 ( 
.A(n_446),
.B(n_289),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_441),
.B(n_288),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_406),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_441),
.B(n_288),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_461),
.B(n_289),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_414),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_415),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_424),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_466),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_421),
.B(n_23),
.Y(n_520)
);

AND2x2_ASAP7_75t_SL g521 ( 
.A(n_434),
.B(n_305),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_427),
.B(n_288),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_453),
.A2(n_288),
.B1(n_307),
.B2(n_305),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_420),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_432),
.A2(n_288),
.B(n_292),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_422),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_437),
.B(n_25),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_423),
.Y(n_528)
);

BUFx4f_ASAP7_75t_L g529 ( 
.A(n_408),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_407),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_440),
.B(n_25),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_464),
.B(n_26),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_395),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_447),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_433),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_425),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g537 ( 
.A(n_427),
.B(n_403),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_399),
.B(n_305),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_412),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_435),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_464),
.A2(n_309),
.B1(n_307),
.B2(n_292),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_442),
.A2(n_309),
.B1(n_307),
.B2(n_292),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_436),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_457),
.B(n_289),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_417),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_429),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_409),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_410),
.B(n_26),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_443),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_410),
.B(n_307),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_403),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_463),
.B(n_27),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_399),
.B(n_309),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_545),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_479),
.B(n_469),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_479),
.B(n_410),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_540),
.B(n_426),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_537),
.B(n_532),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_482),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_545),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_518),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_518),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_486),
.B(n_438),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_482),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_550),
.B(n_451),
.Y(n_565)
);

NAND2x1p5_ASAP7_75t_L g566 ( 
.A(n_502),
.B(n_451),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_470),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_550),
.B(n_458),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_471),
.B(n_465),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_470),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_501),
.B(n_460),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_470),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_516),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_501),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_543),
.B(n_426),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_490),
.B(n_438),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_506),
.B(n_508),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_483),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_543),
.Y(n_579)
);

CKINVDCx6p67_ASAP7_75t_R g580 ( 
.A(n_484),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_508),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_471),
.B(n_449),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_550),
.B(n_448),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_484),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_483),
.B(n_27),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_483),
.B(n_28),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_505),
.B(n_28),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_475),
.B(n_478),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_516),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_502),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_475),
.B(n_29),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_478),
.B(n_29),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_505),
.B(n_30),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_550),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_489),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_502),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_545),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_536),
.B(n_535),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_549),
.B(n_30),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_474),
.B(n_31),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_549),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_474),
.B(n_32),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_535),
.B(n_32),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_536),
.B(n_33),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_501),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_494),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_494),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_520),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_520),
.B(n_552),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_480),
.B(n_33),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_498),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_514),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_497),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_480),
.B(n_34),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_527),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_498),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_514),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_510),
.B(n_309),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_514),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_510),
.B(n_36),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_605),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_579),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_578),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_606),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_605),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_557),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_555),
.B(n_527),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_582),
.A2(n_546),
.B1(n_539),
.B2(n_531),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_606),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_588),
.B(n_531),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_579),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_559),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_588),
.B(n_563),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_607),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_559),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_578),
.Y(n_636)
);

INVx3_ASAP7_75t_SL g637 ( 
.A(n_580),
.Y(n_637)
);

BUFx4_ASAP7_75t_SL g638 ( 
.A(n_584),
.Y(n_638)
);

INVx6_ASAP7_75t_L g639 ( 
.A(n_578),
.Y(n_639)
);

BUFx4_ASAP7_75t_SL g640 ( 
.A(n_584),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_564),
.Y(n_641)
);

BUFx8_ASAP7_75t_L g642 ( 
.A(n_595),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_580),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_585),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_595),
.Y(n_645)
);

BUFx4_ASAP7_75t_SL g646 ( 
.A(n_583),
.Y(n_646)
);

INVx6_ASAP7_75t_SL g647 ( 
.A(n_583),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_554),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_585),
.Y(n_649)
);

INVx8_ASAP7_75t_L g650 ( 
.A(n_565),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_554),
.Y(n_651)
);

CKINVDCx14_ASAP7_75t_R g652 ( 
.A(n_575),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_607),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_585),
.Y(n_654)
);

INVx3_ASAP7_75t_SL g655 ( 
.A(n_583),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_554),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_564),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_585),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_554),
.Y(n_659)
);

INVx5_ASAP7_75t_L g660 ( 
.A(n_612),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_554),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_613),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_613),
.Y(n_663)
);

CKINVDCx8_ASAP7_75t_R g664 ( 
.A(n_583),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_556),
.B(n_548),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_601),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_576),
.B(n_547),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_601),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_574),
.B(n_547),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_575),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_582),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_586),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_560),
.Y(n_673)
);

INVx3_ASAP7_75t_SL g674 ( 
.A(n_620),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_598),
.A2(n_547),
.B1(n_497),
.B2(n_495),
.Y(n_675)
);

BUFx5_ASAP7_75t_L g676 ( 
.A(n_586),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_611),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_676),
.B(n_577),
.Y(n_678)
);

INVx6_ASAP7_75t_L g679 ( 
.A(n_642),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_665),
.B(n_556),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_649),
.A2(n_609),
.B1(n_552),
.B2(n_620),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_671),
.A2(n_615),
.B1(n_539),
.B2(n_521),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_SL g683 ( 
.A1(n_676),
.A2(n_586),
.B1(n_548),
.B2(n_610),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_638),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_671),
.A2(n_521),
.B1(n_609),
.B2(n_569),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_624),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_629),
.Y(n_687)
);

INVx6_ASAP7_75t_L g688 ( 
.A(n_642),
.Y(n_688)
);

BUFx4f_ASAP7_75t_SL g689 ( 
.A(n_631),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_654),
.A2(n_586),
.B1(n_603),
.B2(n_599),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_SL g691 ( 
.A1(n_674),
.A2(n_620),
.B1(n_558),
.B2(n_614),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_634),
.Y(n_692)
);

CKINVDCx6p67_ASAP7_75t_R g693 ( 
.A(n_637),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_SL g694 ( 
.A1(n_676),
.A2(n_610),
.B1(n_495),
.B2(n_599),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_677),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_653),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_SL g697 ( 
.A1(n_676),
.A2(n_599),
.B1(n_600),
.B2(n_602),
.Y(n_697)
);

BUFx10_ASAP7_75t_L g698 ( 
.A(n_669),
.Y(n_698)
);

CKINVDCx11_ASAP7_75t_R g699 ( 
.A(n_637),
.Y(n_699)
);

INVx6_ASAP7_75t_L g700 ( 
.A(n_642),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_662),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_SL g702 ( 
.A1(n_676),
.A2(n_599),
.B1(n_600),
.B2(n_602),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_670),
.A2(n_569),
.B1(n_481),
.B2(n_493),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_654),
.A2(n_561),
.B1(n_562),
.B2(n_608),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_663),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_654),
.A2(n_561),
.B1(n_562),
.B2(n_604),
.Y(n_706)
);

INVx8_ASAP7_75t_L g707 ( 
.A(n_650),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_666),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_631),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_668),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_649),
.A2(n_620),
.B1(n_581),
.B2(n_485),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_652),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_632),
.Y(n_713)
);

AOI22x1_ASAP7_75t_SL g714 ( 
.A1(n_622),
.A2(n_530),
.B1(n_472),
.B2(n_477),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_632),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_635),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_628),
.A2(n_546),
.B1(n_472),
.B2(n_573),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_627),
.A2(n_589),
.B1(n_573),
.B2(n_489),
.Y(n_718)
);

OAI21xp5_ASAP7_75t_SL g719 ( 
.A1(n_672),
.A2(n_592),
.B(n_591),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_635),
.Y(n_720)
);

CKINVDCx11_ASAP7_75t_R g721 ( 
.A(n_626),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_641),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_650),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_SL g724 ( 
.A1(n_652),
.A2(n_530),
.B1(n_476),
.B2(n_574),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_641),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_657),
.Y(n_726)
);

INVxp67_ASAP7_75t_SL g727 ( 
.A(n_644),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_658),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_657),
.Y(n_729)
);

INVx6_ASAP7_75t_L g730 ( 
.A(n_643),
.Y(n_730)
);

BUFx8_ASAP7_75t_SL g731 ( 
.A(n_643),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_633),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_690),
.A2(n_658),
.B1(n_672),
.B2(n_630),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_686),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_684),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_690),
.A2(n_658),
.B1(n_674),
.B2(n_667),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_687),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_685),
.A2(n_665),
.B1(n_545),
.B2(n_589),
.Y(n_738)
);

CKINVDCx11_ASAP7_75t_R g739 ( 
.A(n_699),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_692),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_SL g741 ( 
.A1(n_679),
.A2(n_664),
.B1(n_655),
.B2(n_645),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_683),
.A2(n_545),
.B1(n_534),
.B2(n_515),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_721),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_696),
.Y(n_744)
);

AOI222xp33_ASAP7_75t_L g745 ( 
.A1(n_681),
.A2(n_592),
.B1(n_591),
.B2(n_529),
.C1(n_519),
.C2(n_593),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_731),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_683),
.A2(n_534),
.B1(n_485),
.B2(n_676),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_682),
.A2(n_534),
.B1(n_676),
.B2(n_616),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_724),
.A2(n_626),
.B1(n_669),
.B2(n_655),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_732),
.B(n_626),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_715),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_694),
.A2(n_534),
.B1(n_616),
.B2(n_611),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_SL g753 ( 
.A1(n_679),
.A2(n_664),
.B1(n_645),
.B2(n_646),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_701),
.Y(n_754)
);

AOI222xp33_ASAP7_75t_L g755 ( 
.A1(n_719),
.A2(n_529),
.B1(n_587),
.B2(n_533),
.C1(n_492),
.C2(n_509),
.Y(n_755)
);

BUFx4f_ASAP7_75t_SL g756 ( 
.A(n_709),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_689),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_697),
.A2(n_534),
.B1(n_551),
.B2(n_647),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_702),
.A2(n_551),
.B1(n_647),
.B2(n_517),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_705),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_718),
.A2(n_647),
.B1(n_517),
.B2(n_492),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_SL g762 ( 
.A1(n_714),
.A2(n_675),
.B1(n_650),
.B2(n_594),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_708),
.Y(n_763)
);

OAI222xp33_ASAP7_75t_L g764 ( 
.A1(n_703),
.A2(n_717),
.B1(n_704),
.B2(n_711),
.C1(n_565),
.C2(n_568),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_719),
.A2(n_639),
.B1(n_669),
.B2(n_636),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_704),
.A2(n_680),
.B1(n_691),
.B2(n_695),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_727),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_730),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_691),
.A2(n_533),
.B1(n_529),
.B2(n_650),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_706),
.A2(n_528),
.B1(n_524),
.B2(n_526),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_710),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_SL g772 ( 
.A1(n_706),
.A2(n_594),
.B1(n_509),
.B2(n_565),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_678),
.B(n_651),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_712),
.B(n_621),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_713),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_720),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_707),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_716),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_688),
.A2(n_568),
.B1(n_565),
.B2(n_594),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_688),
.Y(n_780)
);

NOR2x1p5_ASAP7_75t_L g781 ( 
.A(n_693),
.B(n_621),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_730),
.B(n_625),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_698),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_728),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_722),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_725),
.A2(n_528),
.B1(n_524),
.B2(n_526),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_726),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_729),
.A2(n_678),
.B1(n_568),
.B2(n_544),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_SL g789 ( 
.A1(n_700),
.A2(n_568),
.B1(n_625),
.B2(n_491),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_698),
.B(n_651),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_723),
.A2(n_496),
.B1(n_597),
.B2(n_560),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_723),
.A2(n_560),
.B1(n_597),
.B2(n_473),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_774),
.B(n_780),
.C(n_736),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_773),
.B(n_656),
.Y(n_794)
);

OAI222xp33_ASAP7_75t_L g795 ( 
.A1(n_766),
.A2(n_618),
.B1(n_541),
.B2(n_510),
.C1(n_542),
.C2(n_566),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_785),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_745),
.A2(n_560),
.B1(n_597),
.B2(n_700),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_773),
.B(n_656),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_738),
.A2(n_597),
.B1(n_560),
.B2(n_618),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_755),
.A2(n_597),
.B1(n_618),
.B2(n_567),
.Y(n_800)
);

AOI221xp5_ASAP7_75t_SL g801 ( 
.A1(n_733),
.A2(n_571),
.B1(n_37),
.B2(n_38),
.C(n_36),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_SL g802 ( 
.A1(n_765),
.A2(n_707),
.B1(n_723),
.B2(n_673),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_734),
.B(n_659),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_785),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_748),
.A2(n_618),
.B1(n_567),
.B2(n_570),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_761),
.A2(n_572),
.B1(n_570),
.B2(n_639),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_759),
.A2(n_639),
.B1(n_728),
.B2(n_636),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_737),
.B(n_659),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_740),
.B(n_661),
.Y(n_809)
);

OAI221xp5_ASAP7_75t_SL g810 ( 
.A1(n_749),
.A2(n_640),
.B1(n_538),
.B2(n_553),
.C(n_523),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_768),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_SL g812 ( 
.A1(n_764),
.A2(n_566),
.B(n_623),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_769),
.A2(n_572),
.B1(n_639),
.B2(n_707),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_752),
.A2(n_623),
.B1(n_473),
.B2(n_661),
.Y(n_814)
);

OAI21xp33_ASAP7_75t_L g815 ( 
.A1(n_767),
.A2(n_673),
.B(n_566),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_751),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_742),
.A2(n_623),
.B1(n_473),
.B2(n_522),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_762),
.A2(n_623),
.B1(n_507),
.B2(n_499),
.Y(n_818)
);

OAI211xp5_ASAP7_75t_L g819 ( 
.A1(n_771),
.A2(n_488),
.B(n_648),
.C(n_660),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_780),
.B(n_512),
.C(n_511),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_772),
.A2(n_499),
.B1(n_507),
.B2(n_487),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_750),
.A2(n_499),
.B1(n_507),
.B2(n_487),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_744),
.B(n_754),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_758),
.A2(n_500),
.B1(n_503),
.B2(n_504),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_741),
.A2(n_648),
.B1(n_660),
.B2(n_513),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_779),
.A2(n_500),
.B1(n_503),
.B2(n_504),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_788),
.A2(n_648),
.B1(n_512),
.B2(n_525),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_775),
.A2(n_776),
.B1(n_787),
.B2(n_751),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_760),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_763),
.B(n_648),
.Y(n_830)
);

OAI222xp33_ASAP7_75t_L g831 ( 
.A1(n_789),
.A2(n_660),
.B1(n_596),
.B2(n_38),
.C1(n_612),
.C2(n_512),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_790),
.B(n_660),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_753),
.A2(n_660),
.B1(n_619),
.B2(n_617),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_778),
.A2(n_619),
.B1(n_617),
.B2(n_590),
.Y(n_834)
);

AOI222xp33_ASAP7_75t_L g835 ( 
.A1(n_747),
.A2(n_292),
.B1(n_596),
.B2(n_617),
.C1(n_590),
.C2(n_619),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_778),
.A2(n_590),
.B1(n_612),
.B2(n_596),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_SL g837 ( 
.A1(n_777),
.A2(n_45),
.B(n_47),
.Y(n_837)
);

OAI22xp33_ASAP7_75t_L g838 ( 
.A1(n_780),
.A2(n_596),
.B1(n_49),
.B2(n_50),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_790),
.B(n_596),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_SL g840 ( 
.A1(n_777),
.A2(n_596),
.B1(n_51),
.B2(n_52),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_SL g841 ( 
.A1(n_777),
.A2(n_48),
.B(n_55),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_770),
.B(n_57),
.C(n_58),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_786),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_843)
);

OAI221xp5_ASAP7_75t_L g844 ( 
.A1(n_801),
.A2(n_782),
.B1(n_768),
.B2(n_783),
.C(n_791),
.Y(n_844)
);

NAND3xp33_ASAP7_75t_L g845 ( 
.A(n_793),
.B(n_783),
.C(n_743),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_823),
.B(n_784),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_823),
.B(n_829),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_815),
.B(n_784),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_829),
.B(n_781),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_796),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_803),
.B(n_784),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_803),
.B(n_743),
.Y(n_852)
);

OAI221xp5_ASAP7_75t_L g853 ( 
.A1(n_837),
.A2(n_792),
.B1(n_735),
.B2(n_746),
.C(n_777),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_810),
.B(n_777),
.C(n_739),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_798),
.B(n_739),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_L g856 ( 
.A(n_830),
.B(n_735),
.C(n_746),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_808),
.B(n_757),
.Y(n_857)
);

OAI221xp5_ASAP7_75t_L g858 ( 
.A1(n_841),
.A2(n_756),
.B1(n_757),
.B2(n_70),
.C(n_71),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_842),
.A2(n_831),
.B(n_819),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_808),
.B(n_809),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_SL g861 ( 
.A1(n_802),
.A2(n_195),
.B1(n_68),
.B2(n_72),
.Y(n_861)
);

AND4x1_ASAP7_75t_L g862 ( 
.A(n_833),
.B(n_65),
.C(n_79),
.D(n_80),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_809),
.B(n_194),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_797),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_798),
.B(n_193),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_815),
.B(n_833),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_794),
.B(n_87),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_SL g868 ( 
.A1(n_811),
.A2(n_190),
.B1(n_90),
.B2(n_91),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_818),
.A2(n_89),
.B1(n_92),
.B2(n_96),
.Y(n_869)
);

OAI221xp5_ASAP7_75t_L g870 ( 
.A1(n_818),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.C(n_100),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_794),
.B(n_189),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_794),
.B(n_102),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_L g873 ( 
.A(n_842),
.B(n_828),
.C(n_825),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_796),
.B(n_103),
.Y(n_874)
);

AOI221xp5_ASAP7_75t_L g875 ( 
.A1(n_838),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.C(n_110),
.Y(n_875)
);

OA21x2_ASAP7_75t_L g876 ( 
.A1(n_812),
.A2(n_111),
.B(n_113),
.Y(n_876)
);

NAND3xp33_ASAP7_75t_L g877 ( 
.A(n_820),
.B(n_114),
.C(n_119),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_832),
.B(n_120),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_804),
.B(n_121),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_804),
.B(n_122),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_807),
.B(n_839),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_816),
.B(n_187),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_SL g883 ( 
.A1(n_816),
.A2(n_123),
.B1(n_124),
.B2(n_126),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_850),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_846),
.B(n_800),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_873),
.A2(n_799),
.B1(n_813),
.B2(n_814),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_847),
.B(n_860),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_846),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_851),
.B(n_835),
.Y(n_889)
);

AND4x1_ASAP7_75t_L g890 ( 
.A(n_854),
.B(n_859),
.C(n_845),
.D(n_875),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_881),
.B(n_834),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_876),
.Y(n_892)
);

NAND3xp33_ASAP7_75t_L g893 ( 
.A(n_862),
.B(n_840),
.C(n_806),
.Y(n_893)
);

NOR3xp33_ASAP7_75t_L g894 ( 
.A(n_858),
.B(n_795),
.C(n_843),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_881),
.B(n_855),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_849),
.B(n_805),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_856),
.B(n_128),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_848),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_866),
.B(n_817),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_848),
.B(n_827),
.Y(n_900)
);

AO21x2_ASAP7_75t_L g901 ( 
.A1(n_866),
.A2(n_826),
.B(n_824),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_852),
.B(n_836),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_857),
.B(n_821),
.Y(n_903)
);

NOR3xp33_ASAP7_75t_L g904 ( 
.A(n_844),
.B(n_853),
.C(n_868),
.Y(n_904)
);

AOI221xp5_ASAP7_75t_L g905 ( 
.A1(n_870),
.A2(n_861),
.B1(n_869),
.B2(n_864),
.C(n_877),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_863),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_865),
.B(n_822),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_884),
.Y(n_908)
);

AO22x2_ASAP7_75t_L g909 ( 
.A1(n_892),
.A2(n_878),
.B1(n_872),
.B2(n_871),
.Y(n_909)
);

NOR2x1_ASAP7_75t_L g910 ( 
.A(n_898),
.B(n_876),
.Y(n_910)
);

NAND4xp75_ASAP7_75t_L g911 ( 
.A(n_905),
.B(n_876),
.C(n_867),
.D(n_879),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_884),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_895),
.Y(n_913)
);

INVxp67_ASAP7_75t_SL g914 ( 
.A(n_892),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_906),
.Y(n_915)
);

XNOR2xp5_ASAP7_75t_L g916 ( 
.A(n_890),
.B(n_883),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_898),
.B(n_889),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_884),
.Y(n_918)
);

NAND4xp75_ASAP7_75t_L g919 ( 
.A(n_905),
.B(n_879),
.C(n_874),
.D(n_880),
.Y(n_919)
);

NAND2x1p5_ASAP7_75t_L g920 ( 
.A(n_892),
.B(n_890),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_888),
.B(n_874),
.Y(n_921)
);

NOR4xp75_ASAP7_75t_L g922 ( 
.A(n_895),
.B(n_882),
.C(n_130),
.D(n_132),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_917),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_908),
.Y(n_924)
);

XOR2x2_ASAP7_75t_L g925 ( 
.A(n_916),
.B(n_904),
.Y(n_925)
);

OA22x2_ASAP7_75t_L g926 ( 
.A1(n_916),
.A2(n_892),
.B1(n_891),
.B2(n_902),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_912),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_915),
.Y(n_928)
);

XNOR2xp5_ASAP7_75t_L g929 ( 
.A(n_919),
.B(n_891),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_918),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_915),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_913),
.Y(n_932)
);

OA22x2_ASAP7_75t_L g933 ( 
.A1(n_929),
.A2(n_920),
.B1(n_914),
.B2(n_911),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_931),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_923),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_924),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_928),
.Y(n_937)
);

OA22x2_ASAP7_75t_L g938 ( 
.A1(n_925),
.A2(n_920),
.B1(n_914),
.B2(n_902),
.Y(n_938)
);

OA22x2_ASAP7_75t_L g939 ( 
.A1(n_925),
.A2(n_900),
.B1(n_921),
.B2(n_896),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_928),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_926),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_935),
.Y(n_942)
);

XNOR2xp5_ASAP7_75t_L g943 ( 
.A(n_933),
.B(n_926),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_936),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_934),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_940),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_940),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_946),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_943),
.A2(n_933),
.B1(n_938),
.B2(n_939),
.Y(n_949)
);

NAND2xp33_ASAP7_75t_L g950 ( 
.A(n_943),
.B(n_937),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_SL g951 ( 
.A1(n_947),
.A2(n_941),
.B1(n_942),
.B2(n_944),
.Y(n_951)
);

AOI221xp5_ASAP7_75t_L g952 ( 
.A1(n_949),
.A2(n_941),
.B1(n_945),
.B2(n_909),
.C(n_938),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_948),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_951),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_950),
.A2(n_939),
.B1(n_932),
.B2(n_909),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_954),
.A2(n_909),
.B1(n_910),
.B2(n_897),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_952),
.A2(n_894),
.B1(n_893),
.B2(n_896),
.Y(n_957)
);

XNOR2xp5_ASAP7_75t_L g958 ( 
.A(n_955),
.B(n_922),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_SL g959 ( 
.A1(n_953),
.A2(n_893),
.B1(n_899),
.B2(n_886),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_953),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_953),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_961),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_957),
.A2(n_900),
.B1(n_899),
.B2(n_889),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_960),
.B(n_930),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_959),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_956),
.B(n_927),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_958),
.Y(n_967)
);

AO22x2_ASAP7_75t_L g968 ( 
.A1(n_965),
.A2(n_903),
.B1(n_907),
.B2(n_887),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_962),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_963),
.A2(n_903),
.B1(n_907),
.B2(n_885),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_964),
.Y(n_971)
);

NAND4xp75_ASAP7_75t_L g972 ( 
.A(n_966),
.B(n_921),
.C(n_885),
.D(n_888),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_968),
.A2(n_967),
.B1(n_901),
.B2(n_887),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_972),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_969),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_971),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_970),
.A2(n_901),
.B1(n_133),
.B2(n_134),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_974),
.A2(n_901),
.B1(n_135),
.B2(n_138),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_973),
.A2(n_129),
.B1(n_139),
.B2(n_140),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_975),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_976),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_977),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_981),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_980),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_979),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_SL g986 ( 
.A1(n_983),
.A2(n_978),
.B1(n_982),
.B2(n_155),
.Y(n_986)
);

OAI22xp33_ASAP7_75t_L g987 ( 
.A1(n_984),
.A2(n_985),
.B1(n_154),
.B2(n_158),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_987),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_986),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_989),
.A2(n_988),
.B1(n_159),
.B2(n_164),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_989),
.A2(n_149),
.B1(n_165),
.B2(n_167),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_988),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_992)
);

OR2x6_ASAP7_75t_L g993 ( 
.A(n_990),
.B(n_171),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_992),
.Y(n_994)
);

AOI221xp5_ASAP7_75t_L g995 ( 
.A1(n_994),
.A2(n_991),
.B1(n_175),
.B2(n_177),
.C(n_181),
.Y(n_995)
);

AOI211xp5_ASAP7_75t_L g996 ( 
.A1(n_995),
.A2(n_993),
.B(n_182),
.C(n_183),
.Y(n_996)
);


endmodule