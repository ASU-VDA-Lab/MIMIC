module real_jpeg_15609_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_572;
wire n_155;
wire n_405;
wire n_412;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_313;
wire n_42;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_324;
wire n_86;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_572),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_0),
.B(n_573),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_1),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_1),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_1),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_1),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_1),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_1),
.B(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_1),
.A2(n_3),
.B1(n_301),
.B2(n_303),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_1),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_2),
.Y(n_178)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_2),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_3),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_3),
.B(n_241),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_3),
.B(n_369),
.Y(n_368)
);

AOI31xp33_ASAP7_75t_SL g401 ( 
.A1(n_3),
.A2(n_300),
.A3(n_402),
.B(n_404),
.Y(n_401)
);

NAND2x1_ASAP7_75t_SL g443 ( 
.A(n_3),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_3),
.B(n_109),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_3),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_3),
.B(n_516),
.Y(n_515)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_4),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_4),
.Y(n_206)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_4),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_5),
.Y(n_573)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_6),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_6),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_6),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_7),
.Y(n_180)
);

NAND2x1_ASAP7_75t_SL g182 ( 
.A(n_7),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_7),
.B(n_249),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_7),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g319 ( 
.A(n_7),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_7),
.B(n_109),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_7),
.B(n_409),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_7),
.B(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_8),
.B(n_66),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_8),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_8),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_8),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_8),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_8),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_SL g366 ( 
.A(n_8),
.B(n_257),
.Y(n_366)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_9),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g225 ( 
.A(n_9),
.Y(n_225)
);

BUFx4f_ASAP7_75t_L g411 ( 
.A(n_9),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_9),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_10),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_10),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_10),
.B(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_10),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_10),
.B(n_507),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_10),
.B(n_521),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_10),
.B(n_527),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_11),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_11),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_11),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_11),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_11),
.B(n_566),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_12),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_12),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_12),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_13),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_13),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_13),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_13),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_13),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_13),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_13),
.B(n_257),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_14),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_14),
.Y(n_145)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_14),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_14),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_15),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_15),
.B(n_68),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_15),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_15),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_15),
.B(n_374),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_15),
.B(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_15),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_15),
.B(n_324),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_16),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_16),
.B(n_94),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_16),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_16),
.B(n_85),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_16),
.B(n_245),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_16),
.B(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_16),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_16),
.B(n_413),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g183 ( 
.A(n_18),
.Y(n_183)
);

XOR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_560),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_117),
.B(n_559),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2x1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_73),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_24),
.B(n_73),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_55),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_26),
.B(n_41),
.C(n_55),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.C(n_36),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_27),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_27),
.A2(n_33),
.B1(n_48),
.B2(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_SL g563 ( 
.A(n_27),
.B(n_43),
.C(n_50),
.Y(n_563)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_31),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_32),
.Y(n_162)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_32),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_33),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_65),
.C(n_70),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_33),
.A2(n_59),
.B1(n_70),
.B2(n_71),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_35),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_50),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_43),
.A2(n_49),
.B1(n_565),
.B2(n_569),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_46),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_47),
.B(n_108),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_47),
.B(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.C(n_64),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_56),
.A2(n_57),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_63),
.Y(n_221)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_63),
.Y(n_322)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

XOR2x1_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_69),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_70),
.A2(n_71),
.B1(n_107),
.B2(n_164),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_SL g103 ( 
.A(n_71),
.B(n_104),
.C(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_112),
.C(n_113),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_103),
.C(n_110),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_75),
.B(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_92),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_93),
.C(n_97),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.C(n_88),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_77),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_172)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_80),
.Y(n_335)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_81),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_82),
.Y(n_305)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2x1_ASAP7_75t_L g171 ( 
.A(n_88),
.B(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_103),
.B(n_110),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_104),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_107),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_107),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_107),
.B(n_157),
.C(n_165),
.Y(n_189)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21x1_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_290),
.B(n_554),
.Y(n_117)
);

NOR3x1_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_194),
.C(n_284),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_119),
.A2(n_555),
.B(n_558),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_120),
.B(n_122),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_186),
.C(n_191),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_123),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_171),
.C(n_173),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_125),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_139),
.C(n_156),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_126),
.B(n_139),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_129),
.C(n_134),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_138),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.C(n_151),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_140),
.B(n_151),
.Y(n_217)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_144),
.Y(n_445)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_146),
.B(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_150),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_155),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_156),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_161),
.Y(n_268)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_165),
.A2(n_166),
.B1(n_176),
.B2(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_176),
.C(n_179),
.Y(n_175)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_169),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_171),
.B(n_173),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_182),
.C(n_184),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_175),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_219),
.C(n_222),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_176),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_176),
.A2(n_222),
.B1(n_230),
.B2(n_238),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_178),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_179),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_179),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_179),
.A2(n_227),
.B1(n_312),
.B2(n_361),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_182),
.B(n_184),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_182),
.B(n_256),
.C(n_260),
.Y(n_255)
);

XNOR2x2_ASAP7_75t_SL g297 ( 
.A(n_182),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_184),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_184),
.A2(n_213),
.B1(n_214),
.B2(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_186),
.A2(n_191),
.B1(n_192),
.B2(n_288),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g288 ( 
.A(n_186),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.C(n_190),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_187),
.B(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_189),
.B(n_190),
.Y(n_279)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_273),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_195),
.B(n_273),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_231),
.C(n_234),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_196),
.B(n_231),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_215),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_198),
.Y(n_276)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_201),
.B(n_275),
.C(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_213),
.C(n_214),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_202),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_207),
.C(n_212),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_203),
.B(n_212),
.Y(n_253)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_213),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_215),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.C(n_226),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_216),
.B(n_218),
.Y(n_344)
);

XNOR2x1_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_225),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_226),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_227),
.B(n_307),
.C(n_312),
.Y(n_306)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_234),
.B(n_384),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_254),
.C(n_269),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_235),
.B(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.C(n_252),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_236),
.B(n_239),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.C(n_247),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_240),
.A2(n_247),
.B1(n_248),
.B2(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_240),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_244),
.B(n_380),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_246),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_247),
.B(n_439),
.C(n_443),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_247),
.A2(n_248),
.B1(n_439),
.B2(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g353 ( 
.A(n_252),
.B(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_254),
.B(n_270),
.Y(n_341)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_263),
.C(n_266),
.Y(n_254)
);

XNOR2x1_ASAP7_75t_L g337 ( 
.A(n_255),
.B(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_260),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_259),
.Y(n_415)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_263),
.B(n_267),
.Y(n_338)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_264),
.Y(n_522)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_266),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_266),
.A2(n_267),
.B1(n_417),
.B2(n_418),
.Y(n_538)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_278),
.C(n_283),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_277)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_280),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_285),
.A2(n_556),
.B(n_557),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_286),
.B(n_289),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_388),
.B(n_551),
.Y(n_290)
);

NOR2xp67_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_382),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_347),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_293),
.B(n_347),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_339),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_294),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_316),
.C(n_336),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_296),
.B(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.C(n_306),
.Y(n_296)
);

XNOR2x1_ASAP7_75t_L g423 ( 
.A(n_297),
.B(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_299),
.A2(n_300),
.B1(n_306),
.B2(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_302),
.B(n_405),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_306),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_311),
.Y(n_463)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_317),
.A2(n_336),
.B1(n_337),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_317),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_327),
.C(n_334),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_318),
.B(n_377),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_321),
.C(n_323),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_319),
.B(n_323),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_319),
.B(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_319),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_321),
.B(n_400),
.Y(n_399)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx6_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_327),
.A2(n_328),
.B1(n_334),
.B2(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_340),
.A2(n_342),
.B1(n_345),
.B2(n_346),
.Y(n_339)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_340),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_342),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_342),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_386),
.C(n_387),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.C(n_355),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_349),
.A2(n_350),
.B1(n_353),
.B2(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_392),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_376),
.C(n_379),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_357),
.B(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_362),
.C(n_367),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_SL g448 ( 
.A(n_359),
.B(n_449),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_362),
.B(n_367),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_363),
.B(n_366),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_365),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_372),
.C(n_373),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_368),
.A2(n_372),
.B1(n_435),
.B2(n_436),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_372),
.B(n_503),
.C(n_505),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_372),
.A2(n_436),
.B1(n_505),
.B2(n_506),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_373),
.B(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_375),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_379),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_382),
.A2(n_552),
.B(n_553),
.Y(n_551)
);

AND2x2_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_385),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_383),
.B(n_385),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_450),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_394),
.C(n_426),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_391),
.B(n_395),
.Y(n_452)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_398),
.C(n_423),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_398),
.B(n_423),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_401),
.C(n_406),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_401),
.Y(n_431)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_431),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_416),
.C(n_417),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g537 ( 
.A(n_407),
.B(n_538),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_412),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_408),
.B(n_412),
.Y(n_489)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_408),
.A2(n_514),
.B1(n_515),
.B2(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_415),
.Y(n_473)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NOR2x1_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_429),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_429),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_432),
.C(n_448),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_430),
.B(n_549),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_432),
.B(n_448),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_437),
.C(n_446),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_433),
.B(n_543),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_438),
.B(n_447),
.Y(n_543)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_439),
.Y(n_496)
);

INVx8_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

XOR2x2_ASAP7_75t_L g494 ( 
.A(n_443),
.B(n_495),
.Y(n_494)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

NAND3xp33_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_452),
.C(n_453),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_454),
.A2(n_546),
.B(n_550),
.Y(n_453)
);

AOI21x1_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_532),
.B(n_545),
.Y(n_454)
);

OAI21x1_ASAP7_75t_SL g455 ( 
.A1(n_456),
.A2(n_497),
.B(n_531),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_485),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_457),
.B(n_485),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_465),
.C(n_474),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_458),
.B(n_500),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_464),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_464),
.C(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_465),
.A2(n_466),
.B1(n_474),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_471),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_467),
.B(n_471),
.Y(n_504)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_470),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

AO22x1_ASAP7_75t_SL g474 ( 
.A1(n_475),
.A2(n_480),
.B1(n_483),
.B2(n_484),
.Y(n_474)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_475),
.Y(n_483)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_480),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_480),
.B(n_483),
.Y(n_487)
);

INVx6_ASAP7_75t_L g517 ( 
.A(n_481),
.Y(n_517)
);

INVx5_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_484),
.B(n_526),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_491),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_486),
.B(n_492),
.C(n_494),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

MAJx2_ASAP7_75t_L g540 ( 
.A(n_487),
.B(n_489),
.C(n_490),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_494),
.Y(n_491)
);

AOI21x1_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_508),
.B(n_530),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_502),
.Y(n_498)
);

NOR2x1_ASAP7_75t_L g530 ( 
.A(n_499),
.B(n_502),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_503),
.A2(n_504),
.B1(n_511),
.B2(n_512),
.Y(n_510)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_509),
.A2(n_518),
.B(n_529),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_SL g509 ( 
.A(n_510),
.B(n_513),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_510),
.B(n_513),
.Y(n_529)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_515),
.Y(n_524)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_525),
.B(n_528),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_523),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_520),
.B(n_523),
.Y(n_528)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_533),
.B(n_544),
.Y(n_532)
);

NOR2x1p5_ASAP7_75t_L g545 ( 
.A(n_533),
.B(n_544),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_534),
.A2(n_535),
.B1(n_541),
.B2(n_542),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_535),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_536),
.A2(n_537),
.B1(n_539),
.B2(n_540),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_536),
.B(n_540),
.C(n_541),
.Y(n_547)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

NOR2xp67_ASAP7_75t_SL g546 ( 
.A(n_547),
.B(n_548),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_547),
.B(n_548),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_R g560 ( 
.A(n_561),
.B(n_571),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_562),
.B(n_570),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_570),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_564),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_565),
.Y(n_569)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);


endmodule