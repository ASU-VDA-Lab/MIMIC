module real_jpeg_31471_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_290;
wire n_239;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_487;
wire n_493;
wire n_93;
wire n_242;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_0),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_0),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_0),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_0),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_1),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_2),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_3),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_3),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_4),
.Y(n_91)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_4),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_4),
.Y(n_225)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_4),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_5),
.A2(n_195),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_5),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_5),
.A2(n_198),
.B1(n_285),
.B2(n_290),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_5),
.A2(n_198),
.B1(n_342),
.B2(n_346),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_5),
.A2(n_198),
.B1(n_364),
.B2(n_370),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_6),
.Y(n_111)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_6),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_6),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_8),
.A2(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_8),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_8),
.A2(n_150),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_L g440 ( 
.A1(n_8),
.A2(n_108),
.B1(n_150),
.B2(n_441),
.Y(n_440)
);

OAI22xp33_ASAP7_75t_SL g513 ( 
.A1(n_8),
.A2(n_150),
.B1(n_514),
.B2(n_516),
.Y(n_513)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

OAI22x1_ASAP7_75t_SL g65 ( 
.A1(n_10),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_10),
.Y(n_69)
);

AO22x2_ASAP7_75t_SL g114 ( 
.A1(n_10),
.A2(n_69),
.B1(n_115),
.B2(n_118),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_10),
.A2(n_69),
.B1(n_211),
.B2(n_214),
.Y(n_210)
);

OAI22x1_ASAP7_75t_L g243 ( 
.A1(n_10),
.A2(n_69),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_11),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_11),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_12),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_12),
.A2(n_54),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

AO22x1_ASAP7_75t_SL g222 ( 
.A1(n_12),
.A2(n_54),
.B1(n_223),
.B2(n_226),
.Y(n_222)
);

AOI22x1_ASAP7_75t_SL g262 ( 
.A1(n_12),
.A2(n_54),
.B1(n_263),
.B2(n_266),
.Y(n_262)
);

NAND2xp33_ASAP7_75t_SL g455 ( 
.A(n_12),
.B(n_456),
.Y(n_455)
);

OAI32xp33_ASAP7_75t_L g480 ( 
.A1(n_12),
.A2(n_481),
.A3(n_487),
.B1(n_489),
.B2(n_493),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_12),
.B(n_157),
.Y(n_507)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp67_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_21),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_20),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_73),
.B(n_553),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_57),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_23),
.A2(n_316),
.B(n_354),
.Y(n_407)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_24),
.A2(n_398),
.B(n_428),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_25),
.A2(n_317),
.B1(n_320),
.B2(n_353),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_25),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_48),
.B(n_49),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_26),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_26),
.B(n_49),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_26),
.B(n_161),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_26),
.Y(n_373)
);

NOR2x1p5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_38),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_29),
.Y(n_167)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_32),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_32),
.Y(n_185)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_35),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_35),
.Y(n_180)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_38),
.B(n_161),
.Y(n_160)
);

AO22x2_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_41),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_41),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g345 ( 
.A(n_41),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_44),
.Y(n_187)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_60),
.Y(n_59)
);

OAI21x1_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_54),
.B(n_55),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_53),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_56),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_54),
.B(n_61),
.Y(n_219)
);

AOI32xp33_ASAP7_75t_L g445 ( 
.A1(n_54),
.A2(n_446),
.A3(n_449),
.B1(n_454),
.B2(n_455),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_54),
.B(n_490),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_54),
.B(n_529),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_54),
.B(n_204),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_55),
.Y(n_188)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_57),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_59),
.B(n_258),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_60),
.B(n_65),
.Y(n_257)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_61),
.Y(n_378)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OA21x2_ASAP7_75t_SL g377 ( 
.A1(n_63),
.A2(n_363),
.B(n_378),
.Y(n_377)
);

OA21x2_ASAP7_75t_SL g386 ( 
.A1(n_63),
.A2(n_363),
.B(n_378),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_64),
.B(n_160),
.Y(n_301)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_422),
.C(n_429),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_359),
.C(n_400),
.Y(n_74)
);

INVxp33_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_328),
.B(n_330),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_303),
.B(n_306),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_269),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_235),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_80),
.B(n_235),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_168),
.C(n_216),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_81),
.B(n_459),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_158),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_112),
.Y(n_82)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_83),
.B(n_112),
.C(n_158),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_83),
.B(n_377),
.C(n_379),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_83),
.A2(n_380),
.B(n_388),
.Y(n_387)
);

NOR3xp33_ASAP7_75t_L g388 ( 
.A(n_83),
.B(n_348),
.C(n_382),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_83),
.Y(n_395)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_83),
.Y(n_412)
);

OA21x2_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_95),
.B(n_105),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_84),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_84),
.B(n_284),
.Y(n_283)
);

AO22x2_ASAP7_75t_L g319 ( 
.A1(n_84),
.A2(n_95),
.B1(n_243),
.B2(n_284),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_84),
.B(n_105),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_84),
.B(n_440),
.Y(n_474)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_84),
.Y(n_529)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_96),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B1(n_92),
.B2(n_94),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_88),
.Y(n_501)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_90),
.Y(n_201)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_90),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_90),
.Y(n_492)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_91),
.Y(n_209)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_95),
.B(n_105),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_95),
.B(n_243),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_95),
.B(n_440),
.Y(n_439)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_99),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_99),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_104),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_107),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_110),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_111),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_148),
.Y(n_112)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_113),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_114),
.B(n_157),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_L g394 ( 
.A(n_114),
.B(n_157),
.Y(n_394)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_122),
.B(n_149),
.Y(n_231)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_123),
.Y(n_300)
);

NOR2x1_ASAP7_75t_L g326 ( 
.A(n_123),
.B(n_262),
.Y(n_326)
);

AO21x2_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_132),
.B(n_140),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g454 ( 
.A(n_124),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_127),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_141),
.B1(n_143),
.B2(n_145),
.Y(n_140)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_141),
.Y(n_496)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_142),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_148),
.B(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_157),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_157),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_157),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_157),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_159),
.B(n_257),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_168),
.B(n_217),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_189),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_169),
.B(n_189),
.Y(n_253)
);

OAI31xp33_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_173),
.A3(n_177),
.B(n_181),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_186),
.B(n_188),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_186),
.Y(n_346)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_194),
.B(n_202),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_210),
.Y(n_229)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g238 ( 
.A1(n_194),
.A2(n_229),
.B(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_196),
.Y(n_515)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_202),
.B(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_202),
.B(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_210),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_203),
.B(n_513),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_230),
.B(n_234),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_218),
.A2(n_219),
.B(n_220),
.Y(n_437)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_219),
.B(n_220),
.Y(n_234)
);

NOR2x1p5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_228),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_221),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_222),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_222),
.Y(n_318)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp33_ASAP7_75t_SL g530 ( 
.A(n_229),
.B(n_512),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_230),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2x1p5_ASAP7_75t_SL g325 ( 
.A(n_233),
.B(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_251),
.Y(n_235)
);

XOR2x1_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_250),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_250),
.C(n_251),
.Y(n_270)
);

XOR2x2_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_238),
.B(n_240),
.Y(n_302)
);

AO21x2_ASAP7_75t_L g317 ( 
.A1(n_239),
.A2(n_280),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_241),
.B(n_474),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_242),
.B(n_439),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_268),
.C(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_268),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_257),
.A2(n_363),
.B(n_373),
.Y(n_362)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_260),
.Y(n_382)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_262),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_269),
.B(n_551),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_270),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_295),
.B2(n_296),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_277),
.A2(n_283),
.B(n_294),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_278),
.B(n_512),
.Y(n_511)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_294),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_294),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_294),
.B(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_308),
.C(n_310),
.Y(n_307)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_302),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_300),
.A2(n_341),
.B(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_302),
.C(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR3xp33_ASAP7_75t_L g549 ( 
.A(n_306),
.B(n_331),
.C(n_550),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_311),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_311),
.Y(n_329)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_313),
.A2(n_362),
.B1(n_374),
.B2(n_375),
.Y(n_361)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_322),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_333),
.C(n_334),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_SL g444 ( 
.A(n_317),
.B(n_445),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_317),
.A2(n_320),
.B1(n_445),
.B2(n_468),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_320),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_322),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g357 ( 
.A(n_323),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_325),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_326),
.Y(n_471)
);

INVxp33_ASAP7_75t_SL g356 ( 
.A(n_327),
.Y(n_356)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_332),
.B(n_335),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_355),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_351),
.Y(n_336)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_337),
.Y(n_404)
);

XNOR2x1_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_349),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_338),
.B(n_349),
.Y(n_415)
);

NAND2x1_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_347),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_347),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_350),
.B(n_439),
.Y(n_438)
);

INVxp33_ASAP7_75t_SL g403 ( 
.A(n_351),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.C(n_358),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_359),
.A2(n_423),
.B(n_426),
.Y(n_422)
);

NAND3xp33_ASAP7_75t_L g429 ( 
.A(n_359),
.B(n_400),
.C(n_430),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_383),
.B(n_397),
.Y(n_359)
);

OAI31xp33_ASAP7_75t_SL g426 ( 
.A1(n_360),
.A2(n_383),
.A3(n_397),
.B(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_376),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_362),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_362),
.B(n_374),
.C(n_376),
.Y(n_399)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx6_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_389),
.C(n_390),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_385),
.A2(n_389),
.B1(n_396),
.B2(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_385),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_389),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_389),
.A2(n_396),
.B1(n_411),
.B2(n_413),
.Y(n_410)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_391),
.B(n_420),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.C(n_396),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_412),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_398),
.B(n_399),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_416),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_406),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_406),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.C(n_405),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_407),
.B(n_414),
.C(n_418),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_409),
.A2(n_410),
.B1(n_414),
.B2(n_415),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_410),
.Y(n_418)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_411),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_416),
.A2(n_424),
.B(n_425),
.Y(n_423)
);

NOR2x1_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_419),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_549),
.B(n_552),
.Y(n_431)
);

AO21x1_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_460),
.B(n_548),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_458),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_434),
.B(n_458),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_438),
.C(n_444),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_435),
.A2(n_436),
.B1(n_463),
.B2(n_464),
.Y(n_462)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_444),
.Y(n_464)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_445),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx8_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

BUFx6f_ASAP7_75t_SL g456 ( 
.A(n_457),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_461),
.A2(n_475),
.B(n_547),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_465),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_462),
.B(n_465),
.Y(n_547)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.C(n_472),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_467),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_467),
.B(n_543),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_469),
.A2(n_470),
.B1(n_472),
.B2(n_473),
.Y(n_543)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_541),
.B(n_546),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_477),
.A2(n_519),
.B(n_540),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_504),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_478),
.B(n_504),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_502),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_479),
.A2(n_480),
.B1(n_502),
.B2(n_503),
.Y(n_525)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_486),
.Y(n_518)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_497),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_510),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_507),
.B1(n_508),
.B2(n_509),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_506),
.B(n_511),
.C(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_509),
.Y(n_545)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_513),
.B(n_523),
.Y(n_522)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_516),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

AOI21x1_ASAP7_75t_L g519 ( 
.A1(n_520),
.A2(n_526),
.B(n_539),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_525),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_L g539 ( 
.A(n_521),
.B(n_525),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_522),
.B(n_533),
.Y(n_532)
);

BUFx4f_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_531),
.B(n_538),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_530),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_530),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_532),
.B(n_534),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_537),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_544),
.Y(n_541)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_542),
.B(n_544),
.Y(n_546)
);


endmodule