module fake_jpeg_30136_n_539 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_539);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_6),
.B(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_12),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_55),
.B(n_56),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_66),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_58),
.B(n_71),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_1),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_20),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_76),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_78),
.B(n_81),
.Y(n_165)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_19),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g166 ( 
.A(n_82),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_83),
.B(n_87),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_18),
.B(n_1),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g158 ( 
.A(n_92),
.Y(n_158)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_93),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_95),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_21),
.Y(n_99)
);

OR2x4_ASAP7_75t_SL g146 ( 
.A(n_99),
.B(n_49),
.Y(n_146)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_18),
.B(n_1),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_105),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_44),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_54),
.A2(n_49),
.B1(n_51),
.B2(n_48),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_123),
.A2(n_138),
.B1(n_148),
.B2(n_70),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_80),
.A2(n_49),
.B1(n_44),
.B2(n_48),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_56),
.B(n_29),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_38),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g177 ( 
.A(n_146),
.B(n_103),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_73),
.A2(n_53),
.B1(n_45),
.B2(n_41),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_59),
.A2(n_53),
.B1(n_45),
.B2(n_41),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_108),
.B1(n_96),
.B2(n_94),
.Y(n_204)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_64),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_171),
.B(n_178),
.C(n_185),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_173),
.B(n_187),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_175),
.Y(n_259)
);

BUFx8_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_177),
.A2(n_190),
.B(n_210),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_68),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_118),
.A2(n_84),
.B1(n_77),
.B2(n_74),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_180),
.A2(n_204),
.B1(n_121),
.B2(n_132),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_166),
.A2(n_95),
.B1(n_88),
.B2(n_106),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_183),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_91),
.B1(n_92),
.B2(n_43),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_125),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_82),
.B(n_47),
.C(n_43),
.Y(n_187)
);

INVx6_ASAP7_75t_SL g188 ( 
.A(n_158),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_188),
.B(n_219),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_136),
.B(n_44),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_38),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_193),
.B(n_194),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_127),
.A2(n_37),
.B1(n_35),
.B2(n_46),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_37),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_221),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_35),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_199),
.B(n_211),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_139),
.A2(n_92),
.B1(n_46),
.B2(n_52),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_200),
.A2(n_202),
.B1(n_212),
.B2(n_217),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_147),
.A2(n_26),
.B1(n_52),
.B2(n_47),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_138),
.A2(n_60),
.B(n_78),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_203),
.A2(n_112),
.B(n_111),
.Y(n_268)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_134),
.Y(n_207)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_207),
.Y(n_262)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_128),
.Y(n_208)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_208),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_78),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_141),
.A2(n_48),
.B1(n_157),
.B2(n_85),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_111),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_213),
.Y(n_239)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_109),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_214),
.B(n_216),
.Y(n_267)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_215),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_60),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_114),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_218),
.B(n_222),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_122),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_222),
.B1(n_178),
.B2(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_137),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_123),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_155),
.A2(n_48),
.B1(n_63),
.B2(n_62),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_159),
.Y(n_258)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_133),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_170),
.Y(n_263)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_129),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_114),
.A2(n_48),
.B1(n_4),
.B2(n_5),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_227),
.A2(n_243),
.B1(n_251),
.B2(n_244),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_126),
.B1(n_161),
.B2(n_113),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_231),
.A2(n_245),
.B1(n_250),
.B2(n_252),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_174),
.B(n_133),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_237),
.B(n_265),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_171),
.A2(n_113),
.B1(n_161),
.B2(n_126),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_185),
.A2(n_129),
.B1(n_115),
.B2(n_140),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_178),
.A2(n_158),
.B(n_132),
.C(n_159),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_247),
.A2(n_188),
.B(n_197),
.C(n_176),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_185),
.A2(n_140),
.B1(n_116),
.B2(n_119),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_201),
.A2(n_119),
.B1(n_116),
.B2(n_221),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_263),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_173),
.B(n_170),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_195),
.B(n_121),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_269),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_190),
.B(n_17),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_203),
.B1(n_208),
.B2(n_191),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_273),
.A2(n_274),
.B1(n_280),
.B2(n_239),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_186),
.B1(n_196),
.B2(n_183),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_276),
.Y(n_316)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_228),
.Y(n_277)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_193),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_172),
.C(n_187),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_230),
.C(n_257),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_231),
.A2(n_225),
.B1(n_189),
.B2(n_215),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_227),
.A2(n_238),
.B1(n_268),
.B2(n_266),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_282),
.A2(n_285),
.B1(n_246),
.B2(n_235),
.Y(n_310)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_228),
.Y(n_283)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_236),
.B(n_194),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_284),
.Y(n_328)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_242),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_286),
.Y(n_331)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_205),
.CI(n_207),
.CON(n_287),
.SN(n_287)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_287),
.B(n_299),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_238),
.B(n_224),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_179),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_232),
.Y(n_291)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_291),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_237),
.B(n_210),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_294),
.Y(n_323)
);

OAI32xp33_ASAP7_75t_L g293 ( 
.A1(n_264),
.A2(n_197),
.A3(n_213),
.B1(n_218),
.B2(n_219),
.Y(n_293)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_175),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_242),
.Y(n_296)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_296),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_297),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_192),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_300),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_255),
.B(n_209),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_255),
.B(n_182),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_301),
.A2(n_304),
.B1(n_197),
.B2(n_239),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_243),
.B(n_176),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_239),
.B(n_253),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_254),
.B(n_206),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_303),
.B(n_305),
.Y(n_338)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_261),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_247),
.B(n_214),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_234),
.B(n_198),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_252),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_270),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_L g325 ( 
.A1(n_307),
.A2(n_230),
.B(n_262),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_308),
.B(n_281),
.Y(n_349)
);

OA22x2_ASAP7_75t_L g344 ( 
.A1(n_310),
.A2(n_340),
.B1(n_274),
.B2(n_280),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_246),
.B(n_235),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_311),
.Y(n_371)
);

INVx13_ASAP7_75t_L g358 ( 
.A(n_312),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_271),
.A2(n_289),
.B1(n_276),
.B2(n_273),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_317),
.B1(n_318),
.B2(n_302),
.Y(n_351)
);

AND2x2_ASAP7_75t_SL g314 ( 
.A(n_292),
.B(n_260),
.Y(n_314)
);

FAx1_ASAP7_75t_SL g363 ( 
.A(n_314),
.B(n_287),
.CI(n_293),
.CON(n_363),
.SN(n_363)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_329),
.C(n_337),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_271),
.A2(n_230),
.B1(n_260),
.B2(n_234),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_306),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_320),
.B(n_321),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_294),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_322),
.A2(n_335),
.B(n_297),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_L g370 ( 
.A1(n_325),
.A2(n_334),
.B(n_338),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_279),
.B(n_249),
.C(n_232),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_272),
.A2(n_233),
.B(n_241),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_281),
.B(n_249),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_290),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_291),
.Y(n_365)
);

AO22x1_ASAP7_75t_L g340 ( 
.A1(n_282),
.A2(n_259),
.B1(n_262),
.B2(n_257),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_342),
.Y(n_380)
);

OAI32xp33_ASAP7_75t_L g343 ( 
.A1(n_333),
.A2(n_298),
.A3(n_300),
.B1(n_305),
.B2(n_275),
.Y(n_343)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_343),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_351),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_319),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_350),
.Y(n_379)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_349),
.B(n_353),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_284),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_328),
.C(n_315),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_357),
.C(n_362),
.Y(n_378)
);

MAJx2_ASAP7_75t_L g353 ( 
.A(n_323),
.B(n_284),
.C(n_272),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_326),
.B(n_275),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_354),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_313),
.A2(n_272),
.B1(n_285),
.B2(n_302),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_356),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_331),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_288),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_327),
.Y(n_361)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_361),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_287),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_365),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_331),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_233),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_309),
.B(n_283),
.Y(n_367)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_316),
.Y(n_368)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_368),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_328),
.B(n_277),
.C(n_296),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_372),
.C(n_348),
.Y(n_387)
);

OAI21xp33_ASAP7_75t_L g385 ( 
.A1(n_370),
.A2(n_332),
.B(n_334),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_309),
.B(n_301),
.C(n_253),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_308),
.A2(n_295),
.B1(n_248),
.B2(n_304),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_373),
.A2(n_317),
.B1(n_340),
.B2(n_318),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_381),
.A2(n_402),
.B1(n_351),
.B2(n_373),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_342),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_383),
.B(n_397),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_363),
.Y(n_410)
);

A2O1A1O1Ixp25_ASAP7_75t_L g416 ( 
.A1(n_385),
.A2(n_405),
.B(n_379),
.C(n_374),
.D(n_395),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_371),
.A2(n_338),
.B(n_335),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_386),
.A2(n_403),
.B(n_356),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_389),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_321),
.Y(n_388)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_388),
.Y(n_430)
);

XNOR2x1_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_362),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_314),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_396),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_353),
.B(n_314),
.C(n_332),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_395),
.B(n_404),
.C(n_363),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_333),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_346),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_368),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_399),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_371),
.A2(n_340),
.B1(n_320),
.B2(n_339),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_359),
.A2(n_322),
.B(n_311),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_310),
.C(n_316),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_375),
.Y(n_406)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_406),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_407),
.B(n_401),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_386),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_409),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_402),
.Y(n_409)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_367),
.Y(n_411)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_411),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_356),
.Y(n_414)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_414),
.Y(n_456)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_375),
.Y(n_415)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_415),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_416),
.B(n_403),
.Y(n_439)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_417),
.B(n_418),
.Y(n_435)
);

BUFx5_ASAP7_75t_L g418 ( 
.A(n_382),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_419),
.A2(n_420),
.B1(n_427),
.B2(n_376),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_374),
.A2(n_330),
.B1(n_355),
.B2(n_358),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_405),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_421),
.B(n_423),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_376),
.A2(n_330),
.B1(n_344),
.B2(n_358),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_422),
.A2(n_426),
.B1(n_429),
.B2(n_401),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_372),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_349),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_424),
.B(n_433),
.Y(n_449)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_377),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_390),
.A2(n_361),
.B1(n_360),
.B2(n_347),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_400),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_434),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_387),
.B(n_389),
.C(n_378),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_392),
.C(n_391),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_380),
.B(n_241),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_364),
.Y(n_434)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_438),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_439),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_454),
.C(n_455),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_442),
.A2(n_410),
.B1(n_413),
.B2(n_429),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_425),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_445),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_425),
.B(n_391),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_446),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_390),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_450),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_381),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_394),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_451),
.B(n_452),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_393),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_407),
.B(n_344),
.C(n_400),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_419),
.B(n_344),
.C(n_341),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_452),
.B(n_414),
.C(n_422),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_464),
.C(n_471),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_430),
.Y(n_461)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_461),
.Y(n_480)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_463),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_435),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_450),
.B(n_413),
.C(n_411),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_465),
.A2(n_470),
.B1(n_457),
.B2(n_451),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_454),
.A2(n_416),
.B1(n_426),
.B2(n_415),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_417),
.C(n_406),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_440),
.A2(n_418),
.B1(n_428),
.B2(n_336),
.Y(n_472)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_472),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_341),
.Y(n_473)
);

CKINVDCx14_ASAP7_75t_R g488 ( 
.A(n_473),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_444),
.B(n_336),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_476),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_439),
.B(n_229),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_471),
.B(n_436),
.C(n_441),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_478),
.B(n_482),
.C(n_489),
.Y(n_503)
);

OAI321xp33_ASAP7_75t_L g479 ( 
.A1(n_465),
.A2(n_443),
.A3(n_453),
.B1(n_456),
.B2(n_455),
.C(n_446),
.Y(n_479)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_448),
.Y(n_482)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_483),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_460),
.B(n_445),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_8),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_459),
.A2(n_286),
.B(n_229),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_486),
.Y(n_505)
);

AOI31xp33_ASAP7_75t_L g487 ( 
.A1(n_469),
.A2(n_286),
.A3(n_259),
.B(n_240),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_487),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_248),
.C(n_240),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_217),
.C(n_4),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_493),
.C(n_8),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_469),
.A2(n_470),
.B1(n_475),
.B2(n_468),
.Y(n_491)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_491),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_458),
.B(n_17),
.C(n_4),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_485),
.A2(n_475),
.B1(n_466),
.B2(n_467),
.Y(n_494)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_494),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_480),
.A2(n_467),
.B1(n_458),
.B2(n_7),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_495),
.B(n_504),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_491),
.A2(n_17),
.B(n_5),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_496),
.A2(n_498),
.B(n_507),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_483),
.A2(n_3),
.B(n_5),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_477),
.A2(n_488),
.B1(n_490),
.B2(n_489),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_501),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_502),
.B(n_493),
.Y(n_513)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_481),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_8),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_507),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_508),
.B(n_9),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_506),
.B(n_477),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_511),
.A2(n_515),
.B(n_518),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_508),
.C(n_497),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_503),
.B(n_478),
.Y(n_515)
);

AOI21xp33_ASAP7_75t_L g522 ( 
.A1(n_516),
.A2(n_514),
.B(n_510),
.Y(n_522)
);

OAI221xp5_ASAP7_75t_L g521 ( 
.A1(n_517),
.A2(n_519),
.B1(n_498),
.B2(n_500),
.C(n_505),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_482),
.Y(n_518)
);

OA21x2_ASAP7_75t_SL g519 ( 
.A1(n_499),
.A2(n_484),
.B(n_10),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_511),
.A2(n_500),
.B(n_496),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_520),
.B(n_523),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_521),
.B(n_522),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_494),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_524),
.B(n_526),
.Y(n_527)
);

AOI322xp5_ASAP7_75t_L g526 ( 
.A1(n_509),
.A2(n_497),
.A3(n_501),
.B1(n_11),
.B2(n_12),
.C1(n_9),
.C2(n_15),
.Y(n_526)
);

A2O1A1O1Ixp25_ASAP7_75t_L g530 ( 
.A1(n_525),
.A2(n_509),
.B(n_524),
.C(n_510),
.D(n_15),
.Y(n_530)
);

NOR3xp33_ASAP7_75t_L g532 ( 
.A(n_530),
.B(n_11),
.C(n_14),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_529),
.B(n_10),
.C(n_11),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_533),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_532),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_527),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_528),
.B(n_16),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_534),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_537),
.B(n_16),
.Y(n_538)
);

AO21x1_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_16),
.B(n_536),
.Y(n_539)
);


endmodule