module fake_jpeg_17910_n_360 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_360);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_17),
.Y(n_82)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_0),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_54),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_63),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_21),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_59),
.B1(n_39),
.B2(n_57),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_68),
.A2(n_105),
.B1(n_112),
.B2(n_10),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_18),
.B1(n_35),
.B2(n_30),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_70),
.A2(n_76),
.B1(n_83),
.B2(n_90),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_18),
.B1(n_35),
.B2(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_44),
.B(n_27),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_80),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_81),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_13),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_60),
.B1(n_29),
.B2(n_35),
.Y(n_83)
);

NAND2x1_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_15),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_85),
.A2(n_87),
.B(n_12),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_26),
.B(n_29),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_19),
.B1(n_27),
.B2(n_25),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_92),
.B1(n_10),
.B2(n_11),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_37),
.A2(n_20),
.B1(n_23),
.B2(n_30),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_94),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_36),
.B1(n_25),
.B2(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_34),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_41),
.A2(n_23),
.B1(n_20),
.B2(n_26),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_97),
.A2(n_98),
.B1(n_108),
.B2(n_109),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_52),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_34),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_104),
.Y(n_122)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_58),
.B(n_34),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_61),
.A2(n_34),
.B1(n_21),
.B2(n_3),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_53),
.A2(n_34),
.B1(n_21),
.B2(n_3),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_53),
.A2(n_21),
.B1(n_2),
.B2(n_4),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_44),
.B(n_1),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_8),
.B(n_10),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_53),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_53),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_87),
.B1(n_106),
.B2(n_81),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_117),
.A2(n_123),
.B1(n_146),
.B2(n_128),
.Y(n_174)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_66),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_68),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_126),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_8),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_127),
.B(n_164),
.Y(n_199)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_130),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_131),
.A2(n_148),
.B1(n_79),
.B2(n_114),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_13),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_133),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_105),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_93),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_135),
.B(n_138),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_110),
.B1(n_99),
.B2(n_84),
.Y(n_180)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_66),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_85),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_141),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_146),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_93),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_12),
.B(n_13),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_72),
.C(n_102),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_74),
.B(n_12),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_144),
.B(n_149),
.Y(n_205)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_71),
.B(n_104),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_159),
.Y(n_207)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_161),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_82),
.B(n_111),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_158),
.Y(n_167)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_95),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_88),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_160),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_88),
.B(n_101),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_75),
.B(n_106),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_69),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_88),
.B(n_101),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx4_ASAP7_75t_SL g164 ( 
.A(n_79),
.Y(n_164)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_170),
.B(n_174),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_171),
.A2(n_180),
.B1(n_200),
.B2(n_188),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_182),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_134),
.B(n_69),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_175),
.B(n_190),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_183),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_72),
.C(n_102),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_186),
.C(n_199),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_84),
.Y(n_182)
);

AOI32xp33_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_99),
.A3(n_110),
.B1(n_114),
.B2(n_122),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_125),
.B(n_134),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_185),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_156),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_162),
.C(n_121),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_136),
.A2(n_152),
.B1(n_141),
.B2(n_124),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_197),
.B1(n_175),
.B2(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_135),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_164),
.A2(n_150),
.B1(n_127),
.B2(n_133),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_204),
.B(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_149),
.A2(n_129),
.B1(n_137),
.B2(n_130),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_167),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_157),
.A2(n_120),
.B1(n_138),
.B2(n_150),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_143),
.B(n_159),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_165),
.A2(n_145),
.B1(n_118),
.B2(n_143),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_129),
.B(n_160),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_209),
.A2(n_232),
.B(n_241),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_160),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_215),
.Y(n_246)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_151),
.C(n_170),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_151),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_218),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_217),
.A2(n_221),
.B1(n_225),
.B2(n_172),
.Y(n_255)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_208),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_222),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_231),
.C(n_188),
.Y(n_253)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_226),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_183),
.B1(n_182),
.B2(n_179),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_166),
.A2(n_198),
.B1(n_202),
.B2(n_180),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_228),
.A2(n_237),
.B1(n_240),
.B2(n_233),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_205),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_229),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_168),
.A2(n_201),
.B(n_178),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_233),
.Y(n_268)
);

AO22x1_ASAP7_75t_L g234 ( 
.A1(n_201),
.A2(n_192),
.B1(n_184),
.B2(n_190),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_172),
.B(n_211),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_237),
.B(n_239),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_178),
.A2(n_185),
.B1(n_167),
.B2(n_186),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_238),
.A2(n_244),
.B1(n_245),
.B2(n_170),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_202),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_206),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_178),
.A2(n_187),
.B(n_169),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_174),
.A2(n_169),
.B1(n_176),
.B2(n_166),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_176),
.A2(n_181),
.B1(n_203),
.B2(n_188),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_247),
.B(n_266),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_250),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_265),
.C(n_270),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_172),
.B1(n_235),
.B2(n_244),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_259),
.B1(n_263),
.B2(n_247),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_255),
.A2(n_276),
.B1(n_269),
.B2(n_271),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_272),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_211),
.A2(n_214),
.B1(n_221),
.B2(n_224),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_242),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_261),
.B(n_267),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_242),
.B(n_234),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_273),
.B(n_256),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_220),
.B(n_231),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_212),
.B(n_218),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_234),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_225),
.B(n_217),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_269),
.B(n_271),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_223),
.C(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_223),
.B(n_226),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_209),
.B(n_245),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_255),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_219),
.A2(n_239),
.B(n_222),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_213),
.B(n_227),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_274),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_278),
.A2(n_297),
.B(n_289),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_279),
.A2(n_277),
.B1(n_297),
.B2(n_283),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_246),
.B1(n_249),
.B2(n_267),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_280),
.A2(n_288),
.B1(n_290),
.B2(n_282),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_270),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_286),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_282),
.A2(n_251),
.B(n_262),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_268),
.B1(n_254),
.B2(n_272),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_283),
.A2(n_273),
.B1(n_256),
.B2(n_250),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_293),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_252),
.Y(n_285)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_285),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_252),
.Y(n_287)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_246),
.B1(n_259),
.B2(n_257),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_253),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_295),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_248),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_258),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_249),
.B(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_251),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_258),
.B(n_261),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_291),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_SL g322 ( 
.A1(n_302),
.A2(n_309),
.B(n_314),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_275),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_305),
.A2(n_308),
.B(n_311),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_306),
.B(n_317),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_266),
.Y(n_307)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_307),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_286),
.A2(n_262),
.B1(n_292),
.B2(n_300),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_299),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_301),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_301),
.C(n_295),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_278),
.B1(n_298),
.B2(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_315),
.B1(n_302),
.B2(n_314),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_330),
.C(n_304),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_327),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_289),
.Y(n_325)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_325),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_333),
.Y(n_337)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_307),
.B(n_306),
.CI(n_309),
.CON(n_327),
.SN(n_327)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_329),
.B(n_334),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_312),
.C(n_303),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_332),
.A2(n_317),
.B(n_311),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_303),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_318),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_341),
.Y(n_345)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_338),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_332),
.A2(n_319),
.B(n_305),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_340),
.B(n_331),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_329),
.A2(n_308),
.B(n_323),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_327),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_344),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_324),
.B(n_327),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_331),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_348),
.Y(n_354)
);

XOR2x1_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_328),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_349),
.A2(n_322),
.B1(n_340),
.B2(n_342),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_352),
.C(n_353),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_345),
.B(n_333),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_336),
.C(n_330),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_343),
.B(n_347),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_355),
.A2(n_350),
.B(n_339),
.Y(n_357)
);

FAx1_ASAP7_75t_SL g358 ( 
.A(n_357),
.B(n_356),
.CI(n_352),
.CON(n_358),
.SN(n_358)
);

OAI211xp5_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_353),
.B(n_337),
.C(n_341),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_359),
.Y(n_360)
);


endmodule