module fake_netlist_6_623_n_875 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_875);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_875;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_680;
wire n_465;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_772;
wire n_656;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_624;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_652;
wire n_553;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g186 ( 
.A(n_27),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_158),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_17),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_106),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_18),
.Y(n_194)
);

BUFx2_ASAP7_75t_SL g195 ( 
.A(n_84),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_86),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_150),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_95),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_61),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_98),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_102),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_93),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_64),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_139),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_80),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_101),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_136),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_79),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_39),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_125),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_168),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_156),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_177),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_14),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_20),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_46),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_59),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_45),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_17),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_121),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_20),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_99),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_31),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_103),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_67),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_171),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_176),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_52),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_92),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_130),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_107),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_122),
.Y(n_239)
);

BUFx8_ASAP7_75t_SL g240 ( 
.A(n_183),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_153),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_129),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_128),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_26),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_78),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_43),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_71),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_35),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_105),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_21),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_97),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_175),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_90),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_41),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_179),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_42),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_22),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_167),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_56),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_66),
.Y(n_261)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_203),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_189),
.B(n_0),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_199),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_199),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_189),
.B(n_0),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_194),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_228),
.B(n_1),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

AND2x4_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_261),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_188),
.B(n_190),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_224),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_188),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_1),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_211),
.B(n_225),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_199),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_186),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g283 ( 
.A(n_218),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_219),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_191),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_234),
.B(n_2),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_248),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_243),
.B(n_2),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_250),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_187),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_196),
.B(n_3),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_198),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_200),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_205),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_206),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_246),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_208),
.B(n_3),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_212),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_214),
.Y(n_300)
);

AND2x4_ASAP7_75t_L g301 ( 
.A(n_223),
.B(n_4),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_233),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_241),
.B(n_4),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_193),
.Y(n_305)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_248),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_256),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_260),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_264),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_197),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g315 ( 
.A1(n_263),
.A2(n_259),
.B1(n_210),
.B2(n_235),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_263),
.A2(n_238),
.B1(n_254),
.B2(n_253),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_297),
.A2(n_229),
.B1(n_251),
.B2(n_249),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_268),
.A2(n_257),
.B1(n_247),
.B2(n_245),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_276),
.B(n_201),
.Y(n_319)
);

CKINVDCx6p67_ASAP7_75t_R g320 ( 
.A(n_282),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_276),
.A2(n_244),
.B1(n_242),
.B2(n_239),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_293),
.Y(n_322)
);

BUFx6f_ASAP7_75t_SL g323 ( 
.A(n_272),
.Y(n_323)
);

OR2x6_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_195),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_L g326 ( 
.A1(n_268),
.A2(n_237),
.B1(n_236),
.B2(n_232),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_202),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_284),
.A2(n_231),
.B1(n_230),
.B2(n_227),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_L g331 ( 
.A1(n_267),
.A2(n_222),
.B1(n_220),
.B2(n_217),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_L g332 ( 
.A1(n_267),
.A2(n_216),
.B1(n_215),
.B2(n_213),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_204),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_262),
.A2(n_209),
.B1(n_207),
.B2(n_7),
.Y(n_334)
);

AO22x2_ASAP7_75t_L g335 ( 
.A1(n_270),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_L g336 ( 
.A1(n_292),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_L g338 ( 
.A1(n_292),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_304),
.B(n_9),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_290),
.B(n_10),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_262),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_341)
);

AO22x2_ASAP7_75t_L g342 ( 
.A1(n_270),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_291),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_291),
.B(n_14),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_262),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_274),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_286),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_290),
.A2(n_19),
.B1(n_21),
.B2(n_23),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_269),
.B(n_24),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_287),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_R g352 ( 
.A1(n_271),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_305),
.B(n_34),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_280),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_305),
.B(n_36),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_277),
.B(n_185),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_279),
.Y(n_357)
);

AO22x2_ASAP7_75t_L g358 ( 
.A1(n_301),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_287),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_280),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_279),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g362 ( 
.A1(n_298),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_362)
);

NOR2x1p5_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_53),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_279),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_278),
.B(n_54),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_322),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_343),
.Y(n_369)
);

NAND2x1p5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_301),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_313),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_273),
.Y(n_372)
);

XOR2x2_ASAP7_75t_L g373 ( 
.A(n_340),
.B(n_295),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_330),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_337),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_327),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_316),
.B(n_295),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_275),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_360),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_323),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_333),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_308),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_319),
.B(n_278),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_339),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

XNOR2x1_ASAP7_75t_L g395 ( 
.A(n_335),
.B(n_308),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_353),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_355),
.B(n_281),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_288),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_320),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_321),
.B(n_274),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_349),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_331),
.B(n_289),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_317),
.B(n_271),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_314),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_326),
.A2(n_303),
.B(n_307),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_358),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_335),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_324),
.Y(n_410)
);

INVx4_ASAP7_75t_SL g411 ( 
.A(n_341),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_324),
.B(n_275),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_342),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_348),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_318),
.A2(n_303),
.B(n_289),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_315),
.B(n_280),
.Y(n_417)
);

NAND2x1p5_ASAP7_75t_L g418 ( 
.A(n_352),
.B(n_285),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_334),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_362),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_332),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

NAND2x1p5_ASAP7_75t_L g424 ( 
.A(n_338),
.B(n_285),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_322),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_327),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_322),
.Y(n_427)
);

AND2x4_ASAP7_75t_SL g428 ( 
.A(n_320),
.B(n_285),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_322),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_322),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_322),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_319),
.B(n_294),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_327),
.B(n_294),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_325),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_320),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_347),
.B(n_265),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_374),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_419),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_388),
.B(n_55),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_366),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_294),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_428),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_414),
.B(n_400),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_436),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_396),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_399),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_390),
.Y(n_449)
);

AND2x2_ASAP7_75t_SL g450 ( 
.A(n_421),
.B(n_296),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_433),
.Y(n_452)
);

AND2x2_ASAP7_75t_SL g453 ( 
.A(n_402),
.B(n_400),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_367),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_392),
.B(n_296),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_368),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_389),
.B(n_296),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_433),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_416),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_383),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_R g462 ( 
.A(n_435),
.B(n_57),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_401),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_412),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_434),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_432),
.B(n_299),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_416),
.B(n_382),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_436),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_382),
.B(n_299),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_372),
.B(n_299),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_369),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_380),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_425),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_424),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_378),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_427),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_381),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_429),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_372),
.B(n_310),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_373),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_430),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_431),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_397),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_404),
.B(n_310),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_397),
.B(n_398),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_393),
.B(n_394),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_424),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_370),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_370),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_426),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_398),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_415),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_420),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_423),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_403),
.B(n_310),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_405),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_422),
.B(n_311),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_406),
.B(n_58),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_408),
.B(n_311),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_418),
.B(n_409),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_407),
.A2(n_266),
.B(n_265),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_413),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_418),
.B(n_311),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_395),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_379),
.B(n_312),
.Y(n_507)
);

BUFx4f_ASAP7_75t_L g508 ( 
.A(n_386),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_387),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_483),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_483),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_476),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_493),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_507),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g515 ( 
.A(n_488),
.B(n_411),
.Y(n_515)
);

NOR2x1_ASAP7_75t_L g516 ( 
.A(n_491),
.B(n_444),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_476),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_452),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_312),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_504),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_459),
.B(n_452),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_481),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_459),
.B(n_410),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_481),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_482),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_492),
.B(n_312),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_452),
.B(n_411),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_482),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_453),
.B(n_375),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_437),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_484),
.B(n_411),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_504),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_452),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_501),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_484),
.B(n_486),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_453),
.B(n_444),
.Y(n_536)
);

AO21x2_ASAP7_75t_L g537 ( 
.A1(n_497),
.A2(n_60),
.B(n_62),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_453),
.B(n_306),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_437),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_438),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_463),
.B(n_63),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_447),
.B(n_306),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_442),
.B(n_306),
.Y(n_543)
);

NAND2x1p5_ASAP7_75t_L g544 ( 
.A(n_488),
.B(n_265),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_438),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_454),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_496),
.B(n_306),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_489),
.B(n_65),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_489),
.B(n_68),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_474),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_507),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_448),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_470),
.B(n_309),
.Y(n_553)
);

BUFx8_ASAP7_75t_SL g554 ( 
.A(n_447),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_497),
.B(n_309),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_498),
.B(n_309),
.Y(n_556)
);

AO21x2_ASAP7_75t_L g557 ( 
.A1(n_498),
.A2(n_69),
.B(n_70),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_496),
.B(n_309),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_456),
.B(n_265),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_487),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_470),
.B(n_479),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_449),
.B(n_72),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_502),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_487),
.Y(n_564)
);

NAND2x1p5_ASAP7_75t_L g565 ( 
.A(n_500),
.B(n_266),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_448),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_501),
.B(n_73),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_490),
.B(n_74),
.Y(n_568)
);

BUFx12f_ASAP7_75t_L g569 ( 
.A(n_562),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_514),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_554),
.Y(n_571)
);

BUFx12f_ASAP7_75t_L g572 ( 
.A(n_551),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_532),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_536),
.B(n_487),
.Y(n_574)
);

INVx5_ASAP7_75t_L g575 ( 
.A(n_532),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_510),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_520),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_540),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_535),
.B(n_460),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_518),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_511),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_520),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_563),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_531),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_530),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_527),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_527),
.B(n_560),
.Y(n_588)
);

BUFx5_ASAP7_75t_L g589 ( 
.A(n_521),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_515),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_518),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g592 ( 
.A(n_531),
.Y(n_592)
);

CKINVDCx6p67_ASAP7_75t_R g593 ( 
.A(n_515),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_552),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_546),
.Y(n_595)
);

CKINVDCx16_ASAP7_75t_R g596 ( 
.A(n_542),
.Y(n_596)
);

BUFx12f_ASAP7_75t_L g597 ( 
.A(n_523),
.Y(n_597)
);

BUFx12f_ASAP7_75t_L g598 ( 
.A(n_523),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_532),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_546),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_548),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_566),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_539),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_545),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_550),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_512),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_542),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_535),
.B(n_460),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_564),
.Y(n_609)
);

BUFx8_ASAP7_75t_L g610 ( 
.A(n_515),
.Y(n_610)
);

BUFx2_ASAP7_75t_SL g611 ( 
.A(n_533),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_522),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_517),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_529),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_603),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_581),
.Y(n_616)
);

INVx6_ASAP7_75t_L g617 ( 
.A(n_572),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_603),
.Y(n_618)
);

CKINVDCx11_ASAP7_75t_R g619 ( 
.A(n_571),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_579),
.A2(n_536),
.B1(n_446),
.B2(n_516),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_574),
.A2(n_487),
.B1(n_467),
.B2(n_439),
.Y(n_621)
);

CKINVDCx14_ASAP7_75t_R g622 ( 
.A(n_571),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_575),
.Y(n_623)
);

BUFx12f_ASAP7_75t_L g624 ( 
.A(n_597),
.Y(n_624)
);

BUFx2_ASAP7_75t_SL g625 ( 
.A(n_583),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_572),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_573),
.Y(n_627)
);

INVx6_ASAP7_75t_L g628 ( 
.A(n_597),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_578),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_581),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_577),
.Y(n_631)
);

INVx6_ASAP7_75t_L g632 ( 
.A(n_598),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_576),
.Y(n_633)
);

OAI22xp33_ASAP7_75t_L g634 ( 
.A1(n_596),
.A2(n_513),
.B1(n_506),
.B2(n_480),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_578),
.Y(n_635)
);

OAI21xp33_ASAP7_75t_SL g636 ( 
.A1(n_608),
.A2(n_450),
.B(n_446),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_608),
.B(n_561),
.Y(n_637)
);

BUFx5_ASAP7_75t_L g638 ( 
.A(n_586),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_SL g639 ( 
.A1(n_614),
.A2(n_480),
.B1(n_506),
.B2(n_443),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_SL g640 ( 
.A1(n_607),
.A2(n_541),
.B1(n_450),
.B2(n_462),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_575),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_573),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_577),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_594),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_605),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_594),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_602),
.Y(n_647)
);

NAND2x1p5_ASAP7_75t_L g648 ( 
.A(n_577),
.B(n_533),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_614),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_583),
.Y(n_650)
);

INVx8_ASAP7_75t_L g651 ( 
.A(n_598),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_602),
.Y(n_652)
);

INVx6_ASAP7_75t_L g653 ( 
.A(n_569),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_613),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_613),
.Y(n_655)
);

CKINVDCx6p67_ASAP7_75t_R g656 ( 
.A(n_569),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_615),
.Y(n_657)
);

OAI21xp33_ASAP7_75t_L g658 ( 
.A1(n_621),
.A2(n_505),
.B(n_495),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_L g659 ( 
.A1(n_636),
.A2(n_467),
.B(n_538),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_650),
.B(n_588),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g661 ( 
.A1(n_640),
.A2(n_443),
.B(n_464),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_L g662 ( 
.A1(n_645),
.A2(n_585),
.B1(n_592),
.B2(n_495),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_616),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_SL g664 ( 
.A1(n_634),
.A2(n_505),
.B(n_509),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_637),
.B(n_570),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_616),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_630),
.Y(n_667)
);

INVx4_ASAP7_75t_SL g668 ( 
.A(n_627),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_633),
.B(n_570),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_SL g670 ( 
.A1(n_653),
.A2(n_450),
.B1(n_508),
.B2(n_601),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_639),
.A2(n_440),
.B1(n_601),
.B2(n_454),
.Y(n_671)
);

OAI222xp33_ASAP7_75t_L g672 ( 
.A1(n_649),
.A2(n_567),
.B1(n_609),
.B2(n_538),
.C1(n_524),
.C2(n_525),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_SL g673 ( 
.A1(n_626),
.A2(n_509),
.B(n_502),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_653),
.A2(n_440),
.B1(n_454),
.B2(n_446),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_618),
.Y(n_675)
);

BUFx12f_ASAP7_75t_L g676 ( 
.A(n_619),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_622),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_656),
.A2(n_588),
.B1(n_490),
.B2(n_469),
.Y(n_678)
);

AOI222xp33_ASAP7_75t_L g679 ( 
.A1(n_633),
.A2(n_494),
.B1(n_636),
.B2(n_441),
.C1(n_478),
.C2(n_473),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_620),
.A2(n_440),
.B1(n_454),
.B2(n_446),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_630),
.A2(n_494),
.B1(n_612),
.B2(n_606),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_625),
.B(n_609),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_646),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_628),
.A2(n_440),
.B1(n_454),
.B2(n_548),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_624),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_629),
.B(n_534),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_646),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_635),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_SL g689 ( 
.A1(n_648),
.A2(n_471),
.B(n_441),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_SL g690 ( 
.A1(n_617),
.A2(n_508),
.B1(n_610),
.B2(n_589),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_651),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_628),
.A2(n_568),
.B1(n_549),
.B2(n_500),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_644),
.B(n_588),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_651),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_632),
.A2(n_549),
.B1(n_568),
.B2(n_500),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_632),
.A2(n_491),
.B1(n_508),
.B2(n_565),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_SL g697 ( 
.A1(n_617),
.A2(n_610),
.B1(n_589),
.B2(n_500),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_SL g698 ( 
.A1(n_631),
.A2(n_473),
.B(n_471),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_631),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_627),
.Y(n_700)
);

BUFx4f_ASAP7_75t_SL g701 ( 
.A(n_627),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_652),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_652),
.Y(n_703)
);

OAI21xp33_ASAP7_75t_L g704 ( 
.A1(n_655),
.A2(n_456),
.B(n_499),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_647),
.B(n_587),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_655),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_658),
.A2(n_670),
.B1(n_671),
.B2(n_695),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_665),
.B(n_654),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_692),
.A2(n_458),
.B1(n_478),
.B2(n_485),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_663),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_664),
.A2(n_491),
.B1(n_593),
.B2(n_587),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_660),
.A2(n_684),
.B1(n_704),
.B2(n_693),
.Y(n_712)
);

OAI22xp33_ASAP7_75t_L g713 ( 
.A1(n_661),
.A2(n_491),
.B1(n_519),
.B2(n_526),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_673),
.A2(n_593),
.B1(n_590),
.B2(n_604),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_660),
.A2(n_458),
.B1(n_528),
.B2(n_479),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_678),
.A2(n_697),
.B1(n_682),
.B2(n_662),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_669),
.B(n_638),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_SL g718 ( 
.A1(n_696),
.A2(n_659),
.B1(n_537),
.B2(n_557),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_659),
.A2(n_451),
.B1(n_469),
.B2(n_638),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_705),
.B(n_686),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_674),
.A2(n_590),
.B1(n_565),
.B2(n_475),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_679),
.A2(n_451),
.B1(n_638),
.B2(n_515),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_SL g723 ( 
.A1(n_676),
.A2(n_537),
.B1(n_557),
.B2(n_638),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_679),
.A2(n_638),
.B1(n_455),
.B2(n_521),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_SL g725 ( 
.A1(n_681),
.A2(n_610),
.B1(n_589),
.B2(n_611),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_666),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_681),
.A2(n_589),
.B1(n_611),
.B2(n_643),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_698),
.A2(n_526),
.B1(n_519),
.B2(n_643),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_690),
.A2(n_643),
.B1(n_445),
.B2(n_468),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_SL g730 ( 
.A1(n_677),
.A2(n_504),
.B1(n_642),
.B2(n_623),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_688),
.B(n_642),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_680),
.A2(n_455),
.B1(n_558),
.B2(n_547),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_657),
.A2(n_472),
.B1(n_477),
.B2(n_589),
.Y(n_733)
);

OR3x1_ASAP7_75t_L g734 ( 
.A(n_667),
.B(n_642),
.C(n_573),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_689),
.A2(n_589),
.B1(n_559),
.B2(n_504),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_672),
.A2(n_589),
.B1(n_623),
.B2(n_641),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_SL g737 ( 
.A1(n_691),
.A2(n_694),
.B1(n_703),
.B2(n_702),
.Y(n_737)
);

AOI221xp5_ASAP7_75t_L g738 ( 
.A1(n_675),
.A2(n_504),
.B1(n_466),
.B2(n_503),
.C(n_477),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_685),
.A2(n_472),
.B1(n_477),
.B2(n_457),
.Y(n_739)
);

OA21x2_ASAP7_75t_L g740 ( 
.A1(n_683),
.A2(n_556),
.B(n_555),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_700),
.A2(n_457),
.B1(n_465),
.B2(n_461),
.Y(n_741)
);

AOI222xp33_ASAP7_75t_L g742 ( 
.A1(n_687),
.A2(n_461),
.B1(n_465),
.B2(n_553),
.C1(n_472),
.C2(n_556),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_706),
.B(n_699),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_699),
.A2(n_580),
.B1(n_591),
.B2(n_595),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_L g745 ( 
.A1(n_668),
.A2(n_543),
.B(n_544),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_708),
.B(n_668),
.Y(n_746)
);

OAI221xp5_ASAP7_75t_SL g747 ( 
.A1(n_707),
.A2(n_599),
.B1(n_555),
.B2(n_582),
.C(n_595),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_720),
.B(n_668),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_726),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_716),
.B(n_701),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_710),
.B(n_75),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_717),
.B(n_580),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_743),
.B(n_76),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_L g754 ( 
.A(n_723),
.B(n_573),
.C(n_599),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_736),
.B(n_77),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_737),
.A2(n_600),
.B1(n_595),
.B2(n_582),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_737),
.B(n_81),
.Y(n_757)
);

OAI221xp5_ASAP7_75t_L g758 ( 
.A1(n_736),
.A2(n_544),
.B1(n_600),
.B2(n_641),
.C(n_584),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_731),
.B(n_580),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_714),
.A2(n_600),
.B1(n_573),
.B2(n_575),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_713),
.B(n_575),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_735),
.A2(n_591),
.B1(n_575),
.B2(n_584),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_740),
.B(n_82),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_712),
.B(n_719),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_SL g765 ( 
.A(n_709),
.B(n_584),
.C(n_85),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_711),
.A2(n_591),
.B1(n_266),
.B2(n_88),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_718),
.B(n_83),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_725),
.B(n_87),
.Y(n_768)
);

NAND2xp33_ASAP7_75t_SL g769 ( 
.A(n_730),
.B(n_89),
.Y(n_769)
);

NAND3xp33_ASAP7_75t_L g770 ( 
.A(n_741),
.B(n_266),
.C(n_94),
.Y(n_770)
);

NAND3xp33_ASAP7_75t_L g771 ( 
.A(n_742),
.B(n_91),
.C(n_96),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_727),
.B(n_184),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_728),
.A2(n_100),
.B1(n_104),
.B2(n_108),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_727),
.B(n_722),
.Y(n_774)
);

OA211x2_ASAP7_75t_L g775 ( 
.A1(n_757),
.A2(n_745),
.B(n_724),
.C(n_738),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_749),
.B(n_748),
.Y(n_776)
);

NOR3xp33_ASAP7_75t_L g777 ( 
.A(n_765),
.B(n_729),
.C(n_721),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_752),
.B(n_740),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_771),
.A2(n_715),
.B1(n_732),
.B2(n_739),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_763),
.B(n_744),
.Y(n_780)
);

INVxp33_ASAP7_75t_L g781 ( 
.A(n_750),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_746),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_763),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_754),
.B(n_759),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_774),
.B(n_733),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_L g786 ( 
.A(n_757),
.B(n_734),
.C(n_111),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_751),
.Y(n_787)
);

NAND4xp25_ASAP7_75t_L g788 ( 
.A(n_750),
.B(n_110),
.C(n_112),
.D(n_113),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_751),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_764),
.B(n_116),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_753),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_753),
.B(n_755),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_768),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_L g794 ( 
.A(n_767),
.B(n_117),
.C(n_118),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_783),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_776),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_778),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_789),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_782),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_791),
.B(n_755),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_789),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_775),
.A2(n_777),
.B1(n_769),
.B2(n_788),
.Y(n_802)
);

XNOR2xp5_ASAP7_75t_L g803 ( 
.A(n_781),
.B(n_772),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_787),
.Y(n_804)
);

NAND4xp75_ASAP7_75t_SL g805 ( 
.A(n_785),
.B(n_769),
.C(n_747),
.D(n_760),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_784),
.Y(n_806)
);

XOR2xp5_ASAP7_75t_L g807 ( 
.A(n_803),
.B(n_781),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_799),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_795),
.Y(n_809)
);

XNOR2xp5_ASAP7_75t_L g810 ( 
.A(n_802),
.B(n_793),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_806),
.Y(n_811)
);

OAI22x1_ASAP7_75t_L g812 ( 
.A1(n_807),
.A2(n_806),
.B1(n_799),
.B2(n_800),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_811),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_809),
.Y(n_814)
);

XNOR2xp5_ASAP7_75t_L g815 ( 
.A(n_810),
.B(n_792),
.Y(n_815)
);

XOR2x2_ASAP7_75t_L g816 ( 
.A(n_810),
.B(n_805),
.Y(n_816)
);

AOI322xp5_ASAP7_75t_L g817 ( 
.A1(n_816),
.A2(n_808),
.A3(n_793),
.B1(n_785),
.B2(n_779),
.C1(n_797),
.C2(n_780),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_814),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_814),
.Y(n_819)
);

XOR2x2_ASAP7_75t_L g820 ( 
.A(n_815),
.B(n_805),
.Y(n_820)
);

AOI221xp5_ASAP7_75t_L g821 ( 
.A1(n_818),
.A2(n_812),
.B1(n_813),
.B2(n_794),
.C(n_786),
.Y(n_821)
);

OAI322xp33_ASAP7_75t_L g822 ( 
.A1(n_819),
.A2(n_790),
.A3(n_801),
.B1(n_798),
.B2(n_804),
.C1(n_761),
.C2(n_796),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_820),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_823),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_821),
.A2(n_784),
.B1(n_780),
.B2(n_817),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_822),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_823),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_824),
.Y(n_828)
);

AO22x2_ASAP7_75t_L g829 ( 
.A1(n_827),
.A2(n_826),
.B1(n_825),
.B2(n_804),
.Y(n_829)
);

AO22x2_ASAP7_75t_L g830 ( 
.A1(n_827),
.A2(n_770),
.B1(n_756),
.B2(n_784),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_826),
.A2(n_773),
.B1(n_761),
.B2(n_779),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_825),
.B(n_762),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_824),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_827),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_828),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_829),
.A2(n_766),
.B1(n_758),
.B2(n_123),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_833),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_834),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_832),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_830),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_830),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_835),
.Y(n_842)
);

NOR4xp25_ASAP7_75t_L g843 ( 
.A(n_837),
.B(n_831),
.C(n_120),
.D(n_124),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_838),
.B(n_119),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_841),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_839),
.B(n_126),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_840),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_836),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_847),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_845),
.A2(n_836),
.B1(n_135),
.B2(n_137),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_842),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_846),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_844),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_848),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_843),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_845),
.Y(n_856)
);

OAI22x1_ASAP7_75t_L g857 ( 
.A1(n_856),
.A2(n_133),
.B1(n_138),
.B2(n_141),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_855),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_853),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_849),
.Y(n_860)
);

AO22x2_ASAP7_75t_L g861 ( 
.A1(n_851),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_854),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_862)
);

OAI22x1_ASAP7_75t_L g863 ( 
.A1(n_852),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_860),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_861),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_861),
.Y(n_866)
);

INVxp67_ASAP7_75t_SL g867 ( 
.A(n_857),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_863),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_867),
.A2(n_850),
.B1(n_858),
.B2(n_862),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_868),
.A2(n_859),
.B1(n_163),
.B2(n_164),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_869),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_871),
.A2(n_866),
.B1(n_865),
.B2(n_864),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_872),
.Y(n_873)
);

AOI221xp5_ASAP7_75t_L g874 ( 
.A1(n_873),
.A2(n_870),
.B1(n_165),
.B2(n_166),
.C(n_169),
.Y(n_874)
);

AOI211xp5_ASAP7_75t_L g875 ( 
.A1(n_874),
.A2(n_162),
.B(n_170),
.C(n_172),
.Y(n_875)
);


endmodule