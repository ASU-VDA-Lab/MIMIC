module fake_jpeg_22107_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_16),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_28),
.Y(n_53)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_28),
.Y(n_46)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_55),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_25),
.B1(n_21),
.B2(n_26),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_51),
.B1(n_54),
.B2(n_63),
.Y(n_74)
);

FAx1_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_42),
.CI(n_41),
.CON(n_48),
.SN(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_32),
.B(n_1),
.C(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_25),
.B1(n_21),
.B2(n_31),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_39),
.B1(n_44),
.B2(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_60),
.B(n_0),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_30),
.B1(n_27),
.B2(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_31),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_72),
.B(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_76),
.Y(n_98)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_79),
.Y(n_100)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_87),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_83)
);

OA21x2_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_61),
.B(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_0),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_91),
.Y(n_110)
);

NAND2x1p5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_48),
.Y(n_101)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_32),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_55),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_106),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_1),
.C(n_2),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_32),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_52),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_61),
.B1(n_59),
.B2(n_64),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_98),
.B(n_119),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_7),
.C(n_14),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_86),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_92),
.B1(n_76),
.B2(n_91),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_125),
.B1(n_128),
.B2(n_132),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_116),
.B(n_70),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_126),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_118),
.B1(n_97),
.B2(n_114),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_99),
.B(n_85),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_109),
.B1(n_117),
.B2(n_106),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_77),
.C(n_93),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_108),
.C(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_138),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_116),
.B(n_104),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_102),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_112),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_144),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_105),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_136),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_104),
.C(n_103),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_154),
.A2(n_129),
.B1(n_127),
.B2(n_132),
.Y(n_167)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_127),
.B1(n_133),
.B2(n_124),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_166),
.B1(n_143),
.B2(n_141),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_159),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_155),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_154),
.B(n_153),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_175),
.B1(n_170),
.B2(n_174),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_159),
.B(n_152),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_177),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_138),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_144),
.C(n_157),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_176),
.C(n_140),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_143),
.B1(n_156),
.B2(n_165),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_145),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_169),
.A2(n_164),
.B1(n_134),
.B2(n_137),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_184),
.B1(n_79),
.B2(n_107),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_11),
.C(n_13),
.Y(n_189)
);

OAI321xp33_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_158),
.A3(n_148),
.B1(n_126),
.B2(n_150),
.C(n_140),
.Y(n_180)
);

XOR2x2_ASAP7_75t_SL g187 ( 
.A(n_180),
.B(n_182),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_171),
.B1(n_177),
.B2(n_176),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_173),
.A2(n_139),
.B(n_123),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_178),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_189),
.B(n_179),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_183),
.C(n_187),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_183),
.B(n_8),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_193),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_8),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.C(n_15),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_12),
.Y(n_195)
);

INVxp33_ASAP7_75t_SL g197 ( 
.A(n_196),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_198),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_199),
.B(n_6),
.Y(n_200)
);


endmodule