module fake_jpeg_4449_n_313 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_2),
.B(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_39),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_43),
.B(n_12),
.Y(n_92)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_51),
.Y(n_74)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_0),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_18),
.B1(n_17),
.B2(n_35),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_18),
.B1(n_17),
.B2(n_35),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_54),
.A2(n_62),
.B1(n_64),
.B2(n_10),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_17),
.B1(n_18),
.B2(n_35),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_81),
.B1(n_83),
.B2(n_11),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_15),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_56),
.A2(n_70),
.B(n_11),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_60),
.B(n_86),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_20),
.B1(n_29),
.B2(n_30),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_61),
.A2(n_63),
.B1(n_69),
.B2(n_87),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_21),
.B1(n_31),
.B2(n_22),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_30),
.B1(n_29),
.B2(n_16),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_24),
.B1(n_31),
.B2(n_21),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_77),
.Y(n_104)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_16),
.B1(n_24),
.B2(n_22),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_19),
.C(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_73),
.Y(n_116)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_28),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_16),
.Y(n_76)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_34),
.Y(n_78)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_34),
.C(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_27),
.Y(n_84)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_26),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_44),
.A2(n_32),
.B1(n_15),
.B2(n_13),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_32),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_94),
.Y(n_110)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_43),
.B(n_32),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_43),
.B(n_32),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_10),
.Y(n_120)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_101),
.A2(n_125),
.B1(n_80),
.B2(n_65),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_122),
.B(n_80),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g112 ( 
.A1(n_60),
.A2(n_11),
.A3(n_10),
.B1(n_9),
.B2(n_7),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_74),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_74),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_77),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_8),
.B1(n_4),
.B2(n_6),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_92),
.B1(n_70),
.B2(n_97),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_56),
.A2(n_1),
.B1(n_4),
.B2(n_7),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_132),
.B(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_141),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_86),
.C(n_98),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_160),
.C(n_121),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_58),
.B1(n_72),
.B2(n_73),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_67),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_110),
.B1(n_128),
.B2(n_115),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_94),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_146),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_64),
.Y(n_142)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_88),
.Y(n_143)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_62),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_155),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_53),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_154),
.Y(n_180)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_149),
.B(n_126),
.CI(n_112),
.CON(n_176),
.SN(n_176)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_82),
.Y(n_150)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_140),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_153),
.B(n_114),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_SL g153 ( 
.A(n_101),
.B(n_65),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_105),
.A2(n_97),
.B1(n_91),
.B2(n_58),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_156),
.A2(n_159),
.B1(n_124),
.B2(n_117),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_161),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_105),
.A2(n_91),
.B1(n_99),
.B2(n_93),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_89),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_79),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_121),
.A2(n_68),
.B1(n_89),
.B2(n_57),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_161),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_173),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_175),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_135),
.C(n_149),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_188),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_158),
.A2(n_126),
.B1(n_103),
.B2(n_115),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_144),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_128),
.B1(n_103),
.B2(n_113),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_192),
.B1(n_66),
.B2(n_107),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_151),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_131),
.B(n_113),
.Y(n_188)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

INVxp33_ASAP7_75t_SL g207 ( 
.A(n_190),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_100),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_191),
.A2(n_152),
.B(n_148),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_142),
.A2(n_124),
.B1(n_100),
.B2(n_66),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_143),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_199),
.B(n_202),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_200),
.A2(n_167),
.B(n_191),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_186),
.B(n_133),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_165),
.A2(n_169),
.B1(n_164),
.B2(n_193),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_209),
.B1(n_224),
.B2(n_175),
.Y(n_230)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_204),
.B(n_210),
.Y(n_241)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_151),
.B(n_138),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_206),
.A2(n_176),
.B1(n_192),
.B2(n_187),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_157),
.B(n_155),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_221),
.B(n_170),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_165),
.A2(n_164),
.B1(n_179),
.B2(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_185),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_215),
.C(n_222),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_151),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_217),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_154),
.Y(n_219)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_147),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_225),
.B(n_180),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_180),
.A2(n_153),
.B(n_146),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_134),
.C(n_129),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_1),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_207),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_247),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_228),
.B(n_237),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_235),
.B1(n_246),
.B2(n_201),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_238),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_171),
.Y(n_234)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_223),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_166),
.B(n_170),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_245),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_174),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_225),
.B1(n_216),
.B2(n_219),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_191),
.C(n_189),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_244),
.C(n_212),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_243),
.B(n_203),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_200),
.B(n_174),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_184),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_209),
.A2(n_194),
.B1(n_177),
.B2(n_187),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_199),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_248),
.B(n_249),
.CI(n_246),
.CON(n_275),
.SN(n_275)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_260),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_256),
.C(n_258),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_224),
.B1(n_223),
.B2(n_194),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_242),
.C(n_233),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_244),
.C(n_239),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_264),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_221),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_198),
.C(n_222),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_263),
.C(n_228),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_214),
.C(n_208),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_257),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_265),
.B(n_266),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_236),
.Y(n_270)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_277),
.C(n_250),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_243),
.B(n_214),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_253),
.B1(n_218),
.B2(n_231),
.Y(n_287)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_274),
.B(n_278),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_240),
.C(n_227),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_268),
.A2(n_240),
.B1(n_236),
.B2(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_226),
.B1(n_220),
.B2(n_252),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_285),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_217),
.B1(n_230),
.B2(n_213),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_288),
.C(n_269),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_271),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_250),
.C(n_213),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_290),
.B(n_273),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_275),
.A2(n_206),
.B1(n_176),
.B2(n_202),
.Y(n_290)
);

NOR2x1_ASAP7_75t_SL g291 ( 
.A(n_281),
.B(n_275),
.Y(n_291)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_283),
.B(n_272),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_293),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_269),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_288),
.C(n_282),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_295),
.C(n_289),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_300),
.A2(n_301),
.B(n_302),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_241),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_210),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_304),
.B(n_303),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_306),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_279),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_282),
.B1(n_278),
.B2(n_293),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_308),
.B(n_310),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_296),
.Y(n_313)
);


endmodule