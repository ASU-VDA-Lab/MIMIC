module real_jpeg_5816_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_1),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_1),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_1),
.B(n_186),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_1),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_1),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_1),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_1),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_2),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_2),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_2),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_2),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_2),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_2),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_3),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_3),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_3),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_3),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_3),
.B(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_4),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_5),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_5),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_5),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_5),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_5),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_5),
.B(n_348),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_5),
.B(n_389),
.Y(n_388)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_7),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_7),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_7),
.B(n_14),
.Y(n_295)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_8),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_8),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_8),
.Y(n_230)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_10),
.B(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_10),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_10),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_10),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_10),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_10),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_10),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_10),
.B(n_391),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_11),
.Y(n_153)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_11),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_12),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_12),
.B(n_81),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_12),
.B(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_12),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_12),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_12),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_12),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_12),
.B(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_13),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_14),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_14),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_14),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_15),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_15),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_15),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_15),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_15),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_15),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_196),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_194),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_161),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_19),
.B(n_161),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_95),
.C(n_125),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_20),
.B(n_95),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_61),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_22),
.B(n_43),
.C(n_61),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.C(n_40),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_23),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.C(n_30),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_24),
.B(n_53),
.C(n_57),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_24),
.A2(n_57),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_24),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_24),
.A2(n_30),
.B1(n_91),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_24),
.A2(n_91),
.B1(n_361),
.B2(n_366),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_24),
.B(n_366),
.Y(n_408)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_26),
.Y(n_359)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_26),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_27),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_27),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_27),
.A2(n_128),
.B1(n_190),
.B2(n_193),
.Y(n_189)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_29),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_30),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_30),
.B(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_30),
.A2(n_131),
.B1(n_255),
.B2(n_256),
.Y(n_327)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_32),
.Y(n_365)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g356 ( 
.A(n_33),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_34),
.A2(n_40),
.B1(n_51),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_34),
.Y(n_160)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_38),
.Y(n_252)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_39),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_45),
.B1(n_46),
.B2(n_51),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_46),
.B(n_51),
.C(n_60),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_49),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_49),
.Y(n_317)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_50),
.Y(n_192)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_53),
.B(n_221),
.C(n_224),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_53),
.A2(n_93),
.B1(n_221),
.B2(n_285),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_55),
.Y(n_371)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_55),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_57),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_79),
.C(n_89),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_62),
.B(n_79),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_70),
.C(n_74),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_63),
.A2(n_64),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_63),
.B(n_119),
.C(n_124),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_63),
.A2(n_64),
.B1(n_142),
.B2(n_143),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_64),
.B(n_143),
.Y(n_293)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_65),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_66),
.Y(n_383)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_74),
.B2(n_78),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_73),
.Y(n_345)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_73),
.Y(n_376)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.C(n_86),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_86),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_85),
.Y(n_237)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_89),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_116),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_97),
.B(n_98),
.C(n_116),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_111),
.B2(n_112),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_104),
.B1(n_109),
.B2(n_110),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_104),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_104),
.B(n_109),
.C(n_112),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_104),
.B(n_134),
.Y(n_205)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_108),
.Y(n_250)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_108),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_133),
.C(n_135),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_124),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_119),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_122),
.A2(n_124),
.B1(n_174),
.B2(n_177),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_122),
.B(n_249),
.C(n_251),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_122),
.A2(n_124),
.B1(n_251),
.B2(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_125),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_140),
.C(n_158),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_126),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.C(n_138),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_127),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_132),
.B(n_138),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_135),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_140),
.B(n_158),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_154),
.C(n_156),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_141),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.C(n_152),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_142),
.A2(n_143),
.B1(n_152),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_146),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_146),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_151),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_152),
.Y(n_263)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_154),
.A2(n_156),
.B1(n_157),
.B2(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_154),
.Y(n_241)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g442 ( 
.A(n_161),
.Y(n_442)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.CI(n_178),
.CON(n_161),
.SN(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_207),
.C(n_212),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_168),
.A2(n_169),
.B1(n_207),
.B2(n_208),
.Y(n_247)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_174),
.Y(n_177)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.Y(n_184)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_188),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_188),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_190),
.Y(n_193)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI221xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_333),
.B1(n_433),
.B2(n_438),
.C(n_439),
.Y(n_197)
);

NOR3xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_273),
.C(n_277),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_199),
.A2(n_434),
.B(n_437),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_266),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_200),
.B(n_266),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_242),
.C(n_244),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_201),
.B(n_242),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_227),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_202),
.B(n_228),
.C(n_239),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.C(n_219),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_204),
.B(n_220),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_206),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_211),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_212),
.B(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_221),
.Y(n_285)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_224),
.B(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_239),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_235),
.C(n_238),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_265),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_229),
.A2(n_231),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_238),
.Y(n_265)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_244),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_259),
.C(n_264),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.C(n_253),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_246),
.B(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_248),
.A2(n_253),
.B1(n_254),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_248),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_249),
.B(n_310),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_264),
.Y(n_281)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_270),
.C(n_272),
.Y(n_274)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_273),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_274),
.B(n_275),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_304),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_278),
.A2(n_435),
.B(n_436),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_302),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_279),
.B(n_302),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.C(n_300),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_280),
.B(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_282),
.B(n_300),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.C(n_291),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_286),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_288),
.B(n_370),
.Y(n_369)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.C(n_296),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_292),
.A2(n_293),
.B1(n_421),
.B2(n_422),
.Y(n_420)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_331),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_305),
.B(n_331),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.C(n_328),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_306),
.B(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_308),
.B(n_328),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.C(n_326),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_309),
.B(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_312),
.A2(n_326),
.B1(n_327),
.B2(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_312),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_318),
.C(n_323),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_313),
.A2(n_314),
.B1(n_323),
.B2(n_324),
.Y(n_412)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_318),
.B(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_428),
.B(n_432),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_414),
.B(n_427),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_401),
.B(n_413),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_377),
.B(n_400),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_367),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_338),
.B(n_367),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_352),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_339),
.B(n_353),
.C(n_360),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_346),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_340),
.B(n_347),
.C(n_349),
.Y(n_410)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_360),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_357),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_355),
.Y(n_389)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_361),
.Y(n_366)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.C(n_372),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_369),
.A2(n_372),
.B1(n_373),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_369),
.Y(n_398)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_394),
.B(n_399),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_387),
.B(n_393),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_386),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_386),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_384),
.Y(n_395)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_385),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_390),
.Y(n_387)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_396),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_403),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_409),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_410),
.C(n_411),
.Y(n_426)
);

BUFx24_ASAP7_75t_SL g441 ( 
.A(n_404),
.Y(n_441)
);

FAx1_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_407),
.CI(n_408),
.CON(n_404),
.SN(n_404)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_407),
.C(n_408),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_426),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_426),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_423),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_419),
.B2(n_420),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_420),
.C(n_423),
.Y(n_429)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_421),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_429),
.B(n_430),
.Y(n_432)
);


endmodule