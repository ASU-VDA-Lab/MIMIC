module fake_jpeg_9990_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_41),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_43),
.Y(n_55)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_46),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_30),
.B1(n_35),
.B2(n_23),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_49),
.A2(n_53),
.B(n_54),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_51),
.B(n_59),
.Y(n_108)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_66),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_30),
.B1(n_35),
.B2(n_23),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_30),
.B1(n_35),
.B2(n_23),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_22),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_30),
.B1(n_23),
.B2(n_34),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_62),
.A2(n_65),
.B1(n_67),
.B2(n_20),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_18),
.B1(n_22),
.B2(n_28),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_17),
.B1(n_24),
.B2(n_27),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_18),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_14),
.B(n_11),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_17),
.B1(n_20),
.B2(n_24),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_77),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_20),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_97),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_85),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_90),
.Y(n_125)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

CKINVDCx12_ASAP7_75t_R g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_87),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_61),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_89),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_19),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_39),
.Y(n_90)
);

CKINVDCx11_ASAP7_75t_R g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_100),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_92),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_60),
.B(n_0),
.Y(n_95)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_97),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_46),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_36),
.C(n_40),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_45),
.C(n_56),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_33),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_107),
.B1(n_111),
.B2(n_71),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_42),
.B(n_36),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_106),
.B1(n_47),
.B2(n_71),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_110),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_43),
.B1(n_33),
.B2(n_29),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_55),
.A2(n_17),
.B1(n_27),
.B2(n_29),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_25),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_48),
.A2(n_27),
.B1(n_26),
.B2(n_29),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_108),
.B(n_28),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_88),
.B1(n_77),
.B2(n_104),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_109),
.C(n_75),
.Y(n_159)
);

HAxp5_ASAP7_75t_SL g164 ( 
.A(n_118),
.B(n_80),
.CON(n_164),
.SN(n_164)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_127),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_122),
.A2(n_36),
.B(n_26),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_0),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_0),
.Y(n_170)
);

CKINVDCx12_ASAP7_75t_R g127 ( 
.A(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_140),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_28),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_36),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_26),
.Y(n_165)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_142),
.B1(n_168),
.B2(n_131),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_104),
.B1(n_84),
.B2(n_90),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_103),
.B1(n_97),
.B2(n_101),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_147),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_149),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_132),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_155),
.Y(n_194)
);

AO21x2_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_104),
.B(n_97),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_154),
.A2(n_117),
.B1(n_70),
.B2(n_72),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_112),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_103),
.B1(n_101),
.B2(n_88),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_165),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_99),
.B1(n_81),
.B2(n_78),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_160),
.C(n_172),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_87),
.C(n_79),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_106),
.B1(n_79),
.B2(n_95),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_68),
.B1(n_80),
.B2(n_111),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_133),
.B(n_124),
.Y(n_185)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_167),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_112),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_114),
.A2(n_72),
.B1(n_85),
.B2(n_70),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_169),
.B(n_126),
.Y(n_174)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_70),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_86),
.C(n_37),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_174),
.B(n_182),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_116),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_187),
.C(n_193),
.Y(n_214)
);

A2O1A1O1Ixp25_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_122),
.B(n_119),
.C(n_126),
.D(n_133),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_154),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_177),
.A2(n_196),
.B1(n_201),
.B2(n_143),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_116),
.C(n_119),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_180),
.B(n_195),
.C(n_206),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_161),
.B(n_119),
.Y(n_182)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_139),
.A3(n_119),
.B1(n_122),
.B2(n_126),
.Y(n_183)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_143),
.B(n_130),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_184),
.B(n_186),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_198),
.B1(n_146),
.B2(n_173),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_124),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_200),
.B(n_162),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_155),
.B(n_113),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_167),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_120),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_117),
.C(n_127),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_120),
.B1(n_129),
.B2(n_85),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_154),
.B1(n_153),
.B2(n_147),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_199),
.A2(n_170),
.B1(n_37),
.B2(n_26),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_144),
.A2(n_129),
.B(n_31),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_154),
.A2(n_142),
.B1(n_141),
.B2(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_154),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_37),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_210),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_191),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_149),
.Y(n_211)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_211),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_216),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_165),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_219),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_181),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_196),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_221),
.B1(n_225),
.B2(n_227),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_166),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_157),
.C(n_145),
.Y(n_222)
);

OA21x2_ASAP7_75t_SL g249 ( 
.A1(n_222),
.A2(n_66),
.B(n_45),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_178),
.B1(n_182),
.B2(n_201),
.Y(n_237)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_151),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_230),
.B1(n_98),
.B2(n_45),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_170),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_187),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_98),
.B1(n_31),
.B2(n_94),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_231),
.A2(n_98),
.B1(n_94),
.B2(n_66),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_179),
.C(n_175),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_235),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_179),
.C(n_180),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_4),
.Y(n_273)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_183),
.B1(n_174),
.B2(n_176),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_238),
.A2(n_242),
.B1(n_247),
.B2(n_250),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_206),
.C(n_195),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

OAI22x1_ASAP7_75t_SL g247 ( 
.A1(n_226),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_94),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_223),
.Y(n_263)
);

OAI321xp33_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_229),
.A3(n_225),
.B1(n_217),
.B2(n_230),
.C(n_212),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_213),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_66),
.C(n_2),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_213),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_253)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_209),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_210),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_4),
.C(n_5),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_229),
.Y(n_262)
);

AOI31xp33_ASAP7_75t_L g289 ( 
.A1(n_257),
.A2(n_270),
.A3(n_9),
.B(n_14),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_252),
.B(n_215),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_271),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_207),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_264),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_245),
.Y(n_265)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

INVxp33_ASAP7_75t_SL g282 ( 
.A(n_266),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_241),
.A2(n_208),
.B1(n_220),
.B2(n_219),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_267),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_287)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_242),
.B1(n_253),
.B2(n_240),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_224),
.Y(n_270)
);

A2O1A1O1Ixp25_ASAP7_75t_L g271 ( 
.A1(n_238),
.A2(n_218),
.B(n_224),
.C(n_231),
.D(n_12),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_254),
.Y(n_285)
);

BUFx12_ASAP7_75t_L g275 ( 
.A(n_234),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_235),
.C(n_239),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_283),
.C(n_260),
.Y(n_298)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_278),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_258),
.A2(n_237),
.B1(n_244),
.B2(n_236),
.Y(n_279)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_251),
.C(n_248),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_236),
.Y(n_284)
);

OAI221xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_289),
.B1(n_274),
.B2(n_272),
.C(n_273),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_286),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_244),
.B1(n_250),
.B2(n_256),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_285),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_269),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_298),
.C(n_288),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_267),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_297),
.Y(n_305)
);

OAI321xp33_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_294),
.A3(n_295),
.B1(n_286),
.B2(n_281),
.C(n_263),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_273),
.B(n_261),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_274),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_11),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_301),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_281),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_300),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_275),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_302),
.B(n_278),
.Y(n_304)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

AOI31xp67_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_303),
.A3(n_8),
.B(n_11),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_283),
.B1(n_275),
.B2(n_277),
.Y(n_309)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_310),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_312),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_9),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_16),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_13),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_13),
.C(n_8),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_310),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_320),
.C(n_315),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_323),
.B(n_324),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g325 ( 
.A1(n_321),
.A2(n_308),
.A3(n_319),
.B1(n_305),
.B2(n_7),
.C1(n_5),
.C2(n_6),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_6),
.C(n_326),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_328),
.Y(n_329)
);


endmodule