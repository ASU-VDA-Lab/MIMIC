module fake_jpeg_7766_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_26),
.B1(n_32),
.B2(n_27),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_59),
.B1(n_66),
.B2(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_53),
.Y(n_85)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_65),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_32),
.B1(n_26),
.B2(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_39),
.A2(n_26),
.B1(n_32),
.B2(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_69),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_71),
.A2(n_107),
.B1(n_23),
.B2(n_29),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_72),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_75),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_26),
.B(n_22),
.C(n_20),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_102),
.B1(n_106),
.B2(n_109),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_22),
.B(n_20),
.C(n_36),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_82),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_42),
.B1(n_43),
.B2(n_37),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_105),
.B1(n_108),
.B2(n_33),
.Y(n_111)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_86),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_92),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_36),
.C(n_45),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_100),
.Y(n_128)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_21),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_52),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_17),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_17),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_49),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_57),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_98),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_55),
.B(n_22),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_18),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_18),
.B1(n_21),
.B2(n_19),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_63),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_49),
.A2(n_23),
.B(n_21),
.C(n_29),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_58),
.A2(n_43),
.B1(n_37),
.B2(n_46),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_111),
.A2(n_134),
.B1(n_29),
.B2(n_23),
.Y(n_166)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_132),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_43),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_100),
.B(n_77),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_41),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_124),
.C(n_120),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_156),
.C(n_159),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_141),
.B(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_145),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_83),
.B1(n_102),
.B2(n_90),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_150),
.B1(n_164),
.B2(n_166),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_112),
.B(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_147),
.B(n_148),
.Y(n_198)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_72),
.B1(n_73),
.B2(n_103),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_149),
.A2(n_154),
.B1(n_160),
.B2(n_114),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_85),
.B1(n_75),
.B2(n_79),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_155),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_76),
.B1(n_107),
.B2(n_82),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_88),
.C(n_100),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_36),
.B(n_108),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_172),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_108),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_111),
.A2(n_95),
.B1(n_43),
.B2(n_108),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_122),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_162),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_17),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_16),
.B(n_131),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_109),
.B1(n_104),
.B2(n_49),
.Y(n_164)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_167),
.B1(n_121),
.B2(n_101),
.Y(n_201)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_113),
.C(n_119),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_139),
.C(n_33),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_95),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_117),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_119),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_179),
.C(n_180),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_113),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_46),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_186),
.C(n_200),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_182),
.A2(n_191),
.B(n_35),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_188),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_193),
.B1(n_194),
.B2(n_167),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_41),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_196),
.Y(n_227)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_155),
.B(n_41),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_149),
.A2(n_131),
.B1(n_123),
.B2(n_81),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_144),
.A2(n_131),
.B1(n_137),
.B2(n_70),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_126),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_202),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_46),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_151),
.B(n_46),
.C(n_45),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_160),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_154),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_210),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_208),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_214),
.A2(n_191),
.B1(n_200),
.B2(n_195),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_16),
.B1(n_87),
.B2(n_98),
.Y(n_215)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_177),
.A2(n_84),
.B1(n_16),
.B2(n_45),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_225),
.B1(n_30),
.B2(n_31),
.Y(n_240)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_217),
.B(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_178),
.B(n_28),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_219),
.B(n_226),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_189),
.A2(n_28),
.B1(n_30),
.B2(n_25),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_222),
.B(n_224),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g222 ( 
.A1(n_176),
.A2(n_30),
.B(n_25),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_190),
.A2(n_0),
.B(n_1),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_175),
.A2(n_45),
.B1(n_31),
.B2(n_24),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_195),
.B(n_34),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_228),
.B(n_181),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_191),
.B(n_174),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_185),
.A2(n_184),
.B1(n_193),
.B2(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_183),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_255),
.B1(n_221),
.B2(n_216),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_236),
.B(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_239),
.A2(n_246),
.B(n_0),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_240),
.A2(n_245),
.B1(n_249),
.B2(n_221),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_174),
.B(n_12),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_229),
.B(n_210),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_24),
.B1(n_31),
.B2(n_30),
.Y(n_245)
);

AO22x1_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_35),
.B1(n_24),
.B2(n_31),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_35),
.C(n_7),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_253),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_212),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_249)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_224),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_212),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_217),
.Y(n_260)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_230),
.C(n_231),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_264),
.C(n_268),
.Y(n_291)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_231),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_263),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_208),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_230),
.C(n_211),
.Y(n_264)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_269),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_207),
.C(n_213),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_249),
.A2(n_225),
.B1(n_220),
.B2(n_222),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_250),
.C(n_244),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_272),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_251),
.B(n_12),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_275),
.B(n_246),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_35),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_240),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_192),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_7),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_3),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_255),
.Y(n_279)
);

OAI321xp33_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_288),
.A3(n_6),
.B1(n_12),
.B2(n_13),
.C(n_15),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_235),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_284),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_235),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_245),
.Y(n_285)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_247),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_266),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_289),
.A2(n_264),
.B1(n_8),
.B2(n_6),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_274),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_258),
.B(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_261),
.B(n_259),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_294),
.A2(n_3),
.B(n_4),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_303),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_300),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_298),
.B(n_299),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_280),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_6),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_301),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_287),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_305),
.C(n_289),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_277),
.A2(n_13),
.B(n_15),
.Y(n_305)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_291),
.C(n_282),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_309),
.B(n_298),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_291),
.C(n_282),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_295),
.A2(n_283),
.B1(n_284),
.B2(n_286),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_302),
.Y(n_317)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_315),
.B(n_299),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_322),
.B(n_308),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_317),
.B(n_312),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_320),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_314),
.A2(n_296),
.B(n_303),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_306),
.B(n_313),
.Y(n_322)
);

AOI21xp33_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_324),
.B(n_326),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_311),
.Y(n_326)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_325),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_318),
.B(n_321),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_327),
.B(n_309),
.C(n_312),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_5),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_5),
.Y(n_332)
);


endmodule