module fake_jpeg_5115_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx11_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_43),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_18),
.B1(n_20),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_68),
.B1(n_20),
.B2(n_22),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_31),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_58),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_21),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_26),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_35),
.A2(n_30),
.B1(n_18),
.B2(n_32),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_36),
.C(n_42),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_89),
.C(n_94),
.Y(n_122)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_74),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_43),
.Y(n_77)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_77),
.B(n_41),
.CI(n_34),
.CON(n_119),
.SN(n_119)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_18),
.B1(n_20),
.B2(n_43),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_63),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_32),
.B(n_44),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_18),
.B1(n_44),
.B2(n_32),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_93),
.B1(n_66),
.B2(n_50),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_20),
.B1(n_25),
.B2(n_43),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_58),
.A2(n_25),
.B1(n_36),
.B2(n_29),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_46),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_100),
.Y(n_132)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_82),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_112),
.B1(n_36),
.B2(n_65),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_57),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_105),
.A2(n_107),
.B(n_120),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_21),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_110),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_62),
.B1(n_60),
.B2(n_56),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_113),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_69),
.B1(n_82),
.B2(n_94),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_116),
.Y(n_139)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_72),
.B(n_63),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_90),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_33),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_92),
.Y(n_123)
);

BUFx4f_ASAP7_75t_SL g154 ( 
.A(n_123),
.Y(n_154)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_128),
.Y(n_150)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_142),
.Y(n_162)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_133),
.Y(n_166)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_53),
.C(n_72),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_119),
.C(n_105),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_53),
.B(n_81),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_40),
.B(n_88),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_103),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_104),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_112),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_152),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_95),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_157),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_120),
.A3(n_105),
.B1(n_115),
.B2(n_119),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_120),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_164),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_115),
.B1(n_102),
.B2(n_65),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_174),
.B1(n_56),
.B2(n_91),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_140),
.A2(n_102),
.B(n_107),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_163),
.A2(n_160),
.B(n_156),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_107),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_42),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_176),
.B(n_101),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_81),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_173),
.B(n_175),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_36),
.B1(n_56),
.B2(n_80),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_164),
.C(n_168),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_171),
.B(n_127),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_179),
.B(n_187),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_145),
.B1(n_143),
.B2(n_138),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_183),
.B1(n_152),
.B2(n_173),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_146),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_186),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_138),
.B1(n_142),
.B2(n_146),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_146),
.B(n_131),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_189),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_130),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_162),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_147),
.Y(n_192)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

NAND2x1_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_42),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_193),
.A2(n_202),
.B(n_110),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_SL g228 ( 
.A1(n_194),
.A2(n_198),
.B(n_41),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_130),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_48),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_74),
.Y(n_219)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_201),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_169),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_155),
.B(n_133),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_203),
.B(n_125),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_163),
.B(n_158),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_211),
.B1(n_198),
.B2(n_180),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_213),
.B1(n_193),
.B2(n_184),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_197),
.A2(n_153),
.B1(n_157),
.B2(n_159),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_214),
.C(n_215),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_151),
.B1(n_167),
.B2(n_172),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_151),
.C(n_67),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_67),
.C(n_48),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_185),
.B(n_169),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_223),
.C(n_225),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_185),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_108),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_228),
.B(n_189),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_101),
.C(n_42),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_129),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_91),
.C(n_134),
.Y(n_225)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_236),
.B1(n_244),
.B2(n_246),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_238),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_248),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_202),
.C(n_193),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_237),
.C(n_234),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_191),
.B1(n_199),
.B2(n_179),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_194),
.C(n_187),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_188),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_249),
.Y(n_251)
);

AOI211xp5_ASAP7_75t_SL g266 ( 
.A1(n_240),
.A2(n_220),
.B(n_33),
.C(n_34),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_148),
.Y(n_241)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_204),
.A2(n_201),
.B1(n_177),
.B2(n_25),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_205),
.A2(n_76),
.B1(n_87),
.B2(n_31),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_245),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_148),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_144),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_210),
.A2(n_76),
.B1(n_19),
.B2(n_24),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_222),
.A2(n_33),
.B(n_31),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_216),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_255),
.B1(n_266),
.B2(n_265),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_205),
.B1(n_219),
.B2(n_207),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_256),
.B(n_264),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_214),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_260),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_263),
.C(n_264),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_229),
.B(n_207),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_223),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_262),
.B(n_268),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_212),
.C(n_215),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_221),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_144),
.C(n_45),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_45),
.C(n_23),
.Y(n_279)
);

OAI321xp33_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_236),
.A3(n_250),
.B1(n_244),
.B2(n_238),
.C(n_240),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_273),
.B(n_277),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_237),
.B1(n_243),
.B2(n_230),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_275),
.B1(n_282),
.B2(n_283),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_252),
.B1(n_28),
.B2(n_13),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_251),
.A2(n_24),
.B1(n_26),
.B2(n_19),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_252),
.B(n_17),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_16),
.Y(n_296)
);

OA21x2_ASAP7_75t_SL g277 ( 
.A1(n_256),
.A2(n_41),
.B(n_34),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_281),
.C(n_257),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_15),
.C(n_14),
.Y(n_280)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_45),
.C(n_71),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_87),
.B1(n_26),
.B2(n_71),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_263),
.A2(n_71),
.B1(n_23),
.B2(n_28),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_267),
.B(n_253),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_287),
.A2(n_40),
.B1(n_8),
.B2(n_12),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_292),
.C(n_293),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_12),
.B1(n_10),
.B2(n_8),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_34),
.B1(n_41),
.B2(n_13),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_290),
.A2(n_11),
.B1(n_14),
.B2(n_12),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_294),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_71),
.C(n_61),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_61),
.C(n_47),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_271),
.B(n_283),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g295 ( 
.A1(n_274),
.A2(n_10),
.B(n_15),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_295),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_271),
.Y(n_301)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_299),
.B(n_300),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_275),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_303),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_47),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_306),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_28),
.C(n_1),
.Y(n_306)
);

AOI321xp33_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_286),
.A3(n_296),
.B1(n_295),
.B2(n_292),
.C(n_293),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_305),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_313),
.B(n_314),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_28),
.B1(n_10),
.B2(n_2),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_310),
.B(n_312),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_305),
.A3(n_303),
.B1(n_16),
.B2(n_4),
.C1(n_0),
.C2(n_6),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_319),
.B(n_0),
.Y(n_320)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_314),
.A2(n_311),
.A3(n_1),
.B1(n_3),
.B2(n_5),
.C1(n_6),
.C2(n_0),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_315),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_321),
.B(n_5),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_3),
.B(n_5),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_5),
.Y(n_326)
);

AO21x1_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_6),
.B(n_247),
.Y(n_327)
);


endmodule