module real_jpeg_17756_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_370, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_370;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_0),
.A2(n_14),
.B(n_367),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_0),
.B(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_1),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_2),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_2),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_2),
.Y(n_198)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_3),
.Y(n_368)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_4),
.Y(n_244)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_5),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_5),
.Y(n_151)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_5),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_5),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_6),
.A2(n_246),
.B1(n_249),
.B2(n_250),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_6),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_6),
.A2(n_249),
.B1(n_272),
.B2(n_275),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_6),
.A2(n_249),
.B1(n_356),
.B2(n_358),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_7),
.Y(n_95)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_7),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_8),
.A2(n_257),
.B1(n_261),
.B2(n_262),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_8),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_8),
.A2(n_261),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_10),
.Y(n_144)
);

BUFx4f_ASAP7_75t_L g248 ( 
.A(n_10),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_11),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_11),
.A2(n_48),
.B1(n_68),
.B2(n_72),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_11),
.A2(n_48),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_11),
.B(n_24),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_11),
.B(n_196),
.C(n_199),
.Y(n_195)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_12),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g121 ( 
.A(n_12),
.Y(n_121)
);

XOR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_339),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

AO221x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_228),
.B1(n_331),
.B2(n_337),
.C(n_338),
.Y(n_16)
);

AO21x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_178),
.B(n_227),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_154),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_19),
.B(n_154),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_115),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_21),
.B(n_82),
.C(n_115),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_55),
.C(n_64),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_22),
.A2(n_130),
.B1(n_152),
.B2(n_153),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_22),
.A2(n_152),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_22),
.A2(n_153),
.B(n_183),
.C(n_185),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_22),
.A2(n_297),
.B(n_302),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_22),
.B(n_297),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_23),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_23),
.B(n_130),
.Y(n_185)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_23),
.B(n_117),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_23),
.B(n_117),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_23),
.B(n_117),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_34),
.B(n_47),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_24),
.A2(n_34),
.B1(n_47),
.B2(n_355),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_35),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_29),
.Y(n_133)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_30),
.Y(n_136)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_40),
.Y(n_357)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_44),
.Y(n_359)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B(n_51),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_48),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_48),
.B(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_48),
.A2(n_111),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_48),
.B(n_138),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_48),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_51),
.A2(n_162),
.A3(n_164),
.B1(n_167),
.B2(n_173),
.Y(n_161)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_55),
.A2(n_65),
.B1(n_66),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_57),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_124),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_65),
.B1(n_83),
.B2(n_114),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_64),
.B(n_161),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_64),
.B(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_64),
.B(n_153),
.C(n_192),
.Y(n_222)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_65),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_65),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_65),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_65),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_65),
.B(n_83),
.Y(n_312)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_77),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_67),
.A2(n_237),
.B1(n_245),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_71),
.A2(n_139),
.B1(n_141),
.B2(n_143),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_71),
.Y(n_199)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_71),
.Y(n_240)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_71),
.Y(n_251)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_75),
.Y(n_212)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_77),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_79),
.Y(n_254)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_79),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_81),
.Y(n_216)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_90),
.B(n_100),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B(n_110),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_129),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_116),
.A2(n_265),
.B1(n_278),
.B2(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_116),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_116),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_117),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_117),
.B(n_130),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_121),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_129),
.A2(n_183),
.B1(n_184),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_129),
.Y(n_224)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_130),
.A2(n_153),
.B1(n_159),
.B2(n_160),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_130),
.A2(n_153),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_130),
.A2(n_153),
.B1(n_194),
.B2(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_130),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_130),
.B(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_130),
.A2(n_153),
.B1(n_236),
.B2(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_130),
.A2(n_153),
.B1(n_282),
.B2(n_322),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_131),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_268)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_133),
.Y(n_299)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g352 ( 
.A(n_137),
.B(n_298),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_145),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_138),
.Y(n_270)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_145),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_147),
.Y(n_301)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.C(n_177),
.Y(n_154)
);

XOR2x2_ASAP7_75t_SL g180 ( 
.A(n_155),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

OAI21x1_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_186),
.B(n_226),
.Y(n_178)
);

NOR2xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_182),
.Y(n_226)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AND3x1_ASAP7_75t_L g324 ( 
.A(n_185),
.B(n_286),
.C(n_325),
.Y(n_324)
);

AOI21x1_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_221),
.B(n_225),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_202),
.B(n_220),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_193),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_200),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_217),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_315),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_303),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_230),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_287),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_231),
.B(n_287),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_264),
.C(n_279),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_232),
.B(n_264),
.Y(n_314)
);

OAI22x1_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_263),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_233),
.B(n_312),
.Y(n_318)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_234),
.A2(n_281),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_234),
.Y(n_307)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_235),
.A2(n_280),
.B(n_284),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_236),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_245),
.B1(n_252),
.B2(n_255),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_267),
.B1(n_268),
.B2(n_278),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_R g292 ( 
.A(n_265),
.B(n_268),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_298),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_278),
.A2(n_348),
.B1(n_363),
.B2(n_370),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B(n_284),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_280),
.A2(n_284),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_295),
.B2(n_296),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_291),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_292),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_295),
.B(n_342),
.C(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_302),
.A2(n_346),
.B1(n_347),
.B2(n_360),
.Y(n_345)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_302),
.Y(n_360)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_303),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_313),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_313),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.C(n_311),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_309),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_327),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_326),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_326),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_321),
.C(n_323),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_323),
.B2(n_324),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_329),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_334),
.B(n_335),
.C(n_336),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_365),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.Y(n_340)
);

NOR2xp67_ASAP7_75t_SL g366 ( 
.A(n_341),
.B(n_344),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_361),
.B1(n_362),
.B2(n_364),
.Y(n_344)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_345),
.Y(n_364)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);


endmodule