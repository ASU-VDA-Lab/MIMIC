module fake_jpeg_5454_n_187 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_38),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_16),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_57),
.Y(n_72)
);

NAND2x1_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_25),
.Y(n_44)
);

AO22x1_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_50),
.B1(n_25),
.B2(n_39),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_27),
.B1(n_18),
.B2(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_54),
.B1(n_60),
.B2(n_15),
.Y(n_73)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_24),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_18),
.B1(n_27),
.B2(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_33),
.A2(n_27),
.B1(n_18),
.B2(n_17),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_62),
.Y(n_88)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_78),
.Y(n_83)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_68),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_19),
.B1(n_31),
.B2(n_15),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_22),
.Y(n_87)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_39),
.B1(n_32),
.B2(n_24),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_58),
.B1(n_53),
.B2(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_75),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_21),
.B1(n_23),
.B2(n_20),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_85),
.B1(n_86),
.B2(n_91),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_28),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_81),
.B(n_25),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_75),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_56),
.B1(n_48),
.B2(n_53),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_22),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g89 ( 
.A(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_80),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_55),
.B1(n_52),
.B2(n_43),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_59),
.B1(n_19),
.B2(n_21),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_77),
.B(n_76),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_21),
.B1(n_23),
.B2(n_20),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_26),
.B1(n_78),
.B2(n_94),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_99),
.B1(n_90),
.B2(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_64),
.B(n_20),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_70),
.B1(n_62),
.B2(n_61),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_81),
.B1(n_80),
.B2(n_65),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_70),
.C(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_103),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_106),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_24),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_25),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_24),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_24),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_81),
.B1(n_99),
.B2(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_114),
.A2(n_116),
.B1(n_94),
.B2(n_95),
.Y(n_118)
);

NOR2x1_ASAP7_75t_R g129 ( 
.A(n_115),
.B(n_49),
.Y(n_129)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_119),
.B(n_129),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_120),
.B1(n_127),
.B2(n_104),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_91),
.B(n_86),
.Y(n_119)
);

XOR2x2_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_32),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_125),
.C(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_100),
.Y(n_139)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_39),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_95),
.B1(n_30),
.B2(n_24),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_128),
.B(n_132),
.Y(n_134)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_49),
.Y(n_146)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_138),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_111),
.C(n_106),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_142),
.C(n_147),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_131),
.C(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_105),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_0),
.Y(n_157)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_101),
.C(n_116),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_143),
.B(n_148),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_146),
.B1(n_129),
.B2(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_0),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_49),
.C(n_1),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_156),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_125),
.B1(n_132),
.B2(n_122),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_145),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_124),
.B1(n_119),
.B2(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_160),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_139),
.B1(n_138),
.B2(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_13),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_164),
.C(n_167),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_151),
.B(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_136),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_160),
.C(n_13),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_150),
.B1(n_156),
.B2(n_153),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_157),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_153),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_173),
.B(n_174),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_161),
.Y(n_175)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_166),
.Y(n_176)
);

AOI31xp67_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_175),
.A3(n_172),
.B(n_165),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_8),
.B(n_10),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_170),
.C(n_176),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_181),
.B(n_182),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_173),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_184),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_186),
.Y(n_187)
);


endmodule