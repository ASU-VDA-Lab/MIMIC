module real_jpeg_26308_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_1),
.B(n_54),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_4),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_4),
.B(n_27),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_54),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_4),
.B(n_51),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_4),
.B(n_33),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_4),
.B(n_17),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_4),
.B(n_49),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_4),
.B(n_69),
.Y(n_271)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_6),
.B(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_6),
.B(n_49),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_6),
.B(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_6),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_6),
.B(n_33),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_6),
.B(n_54),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_6),
.B(n_51),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_7),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_7),
.B(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_7),
.B(n_54),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_7),
.B(n_69),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_7),
.B(n_270),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_9),
.B(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_9),
.B(n_51),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_9),
.B(n_49),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_9),
.B(n_54),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_9),
.B(n_33),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_9),
.B(n_37),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_9),
.B(n_69),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_9),
.B(n_27),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_10),
.B(n_49),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_10),
.B(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_10),
.B(n_17),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_10),
.B(n_33),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_10),
.B(n_54),
.Y(n_292)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_13),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_13),
.B(n_33),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_13),
.B(n_54),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_13),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_13),
.B(n_51),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_13),
.B(n_49),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_13),
.B(n_69),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_14),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_14),
.B(n_27),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_14),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_14),
.B(n_174),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_14),
.B(n_33),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_14),
.B(n_54),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_15),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_15),
.B(n_51),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_15),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_15),
.B(n_49),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_16),
.B(n_49),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_16),
.B(n_69),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_16),
.B(n_51),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_16),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_16),
.B(n_33),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_16),
.B(n_27),
.Y(n_242)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_17),
.Y(n_115)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_17),
.Y(n_175)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_17),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_149),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_119),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.C(n_92),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_21),
.B(n_80),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_56),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_22),
.B(n_57),
.C(n_74),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.C(n_47),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_23),
.B(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_30),
.C(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_26),
.B(n_63),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_30),
.A2(n_40),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_30),
.B(n_82),
.C(n_85),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_31),
.B(n_64),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_32),
.B(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_35),
.A2(n_39),
.B1(n_42),
.B2(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_42),
.C(n_43),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_41),
.B(n_47),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_42),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_43),
.A2(n_44),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_46),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_47),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_50),
.CI(n_53),
.CON(n_47),
.SN(n_47)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_50),
.C(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_54),
.Y(n_216)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_74),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_68),
.C(n_72),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_58),
.A2(n_59),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.C(n_65),
.Y(n_59)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_62),
.CI(n_65),
.CON(n_94),
.SN(n_94)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_72),
.B1(n_78),
.B2(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_68),
.B(n_77),
.C(n_79),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_72),
.Y(n_107)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_73),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_76),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_87),
.C(n_88),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_85),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_88),
.Y(n_331)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_90),
.CI(n_91),
.CON(n_88),
.SN(n_88)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_90),
.C(n_91),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_92),
.B(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_105),
.C(n_109),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_93),
.B(n_105),
.CI(n_109),
.CON(n_324),
.SN(n_324)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.C(n_101),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_94),
.B(n_308),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_94),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_95),
.B(n_101),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.C(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_98),
.B(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_117),
.C(n_118),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_110),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_110),
.B(n_314),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.CI(n_116),
.CON(n_110),
.SN(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_117),
.B(n_118),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_134),
.B2(n_135),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_130),
.B2(n_131),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_128),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_147),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_326),
.C(n_327),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_317),
.C(n_318),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_303),
.C(n_304),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_281),
.C(n_282),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_249),
.C(n_250),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_224),
.C(n_225),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_185),
.C(n_198),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_170),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_165),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_158),
.B(n_165),
.C(n_170),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_160),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_168),
.C(n_169),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_171),
.B(n_179),
.C(n_180),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_175),
.Y(n_270)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_182),
.B(n_184),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_197),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_190),
.B1(n_197),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_220),
.C(n_221),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_207),
.C(n_212),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_205),
.C(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.C(n_217),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_215),
.B(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_238),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_239),
.C(n_248),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_233),
.C(n_234),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_229),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_232),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_234),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.CI(n_237),
.CON(n_234),
.SN(n_234)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_236),
.C(n_237),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_248),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_242),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_245),
.C(n_247),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_246),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_265),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_254),
.C(n_265),
.Y(n_281)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_260),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_261),
.C(n_264),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_256),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_258),
.CI(n_259),
.CON(n_256),
.SN(n_256)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_258),
.C(n_259),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_273),
.C(n_279),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_273),
.B1(n_279),
.B2(n_280),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_268),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_271),
.B(n_272),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_271),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_300),
.C(n_301),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_273),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_277),
.C(n_278),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_296),
.B2(n_302),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_297),
.C(n_298),
.Y(n_303)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_287),
.C(n_289),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_295),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_294),
.C(n_295),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_293),
.Y(n_294)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_296),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_315),
.B2(n_316),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_305),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_309),
.C(n_315),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_321),
.C(n_325),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_324),
.Y(n_333)
);


endmodule