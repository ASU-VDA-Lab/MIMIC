module fake_netlist_5_482_n_1847 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1847);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1847;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_798;
wire n_350;
wire n_196;
wire n_215;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_61),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_89),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_172),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_99),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_136),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_20),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_160),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_124),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_84),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_110),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_42),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_92),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_14),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_61),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_1),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_63),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_101),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_96),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_40),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_164),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_30),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_142),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_73),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_122),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_137),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_100),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_62),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_55),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_9),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_95),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_104),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_79),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_5),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_106),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_93),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_55),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_147),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_28),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_111),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_94),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_105),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_156),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_13),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_46),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_120),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_49),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_116),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_150),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_3),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_65),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_14),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_40),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_149),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_21),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_135),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_50),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_26),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_62),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_109),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_102),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_157),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_66),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_16),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_2),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_117),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_43),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_27),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_41),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_71),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_143),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_125),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_127),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_166),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_34),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_107),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_67),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_129),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_145),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_97),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_28),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_151),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_76),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_159),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_123),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_50),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_91),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_141),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_19),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_15),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_90),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_60),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_10),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_128),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_167),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_45),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_8),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_132),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_56),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_31),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_130),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_77),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_49),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_25),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_8),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_12),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_48),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_4),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_72),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_33),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_15),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_51),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_85),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_30),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_58),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_114),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_48),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_78),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_17),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_87),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_53),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_12),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_18),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_5),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_45),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_83),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_51),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_108),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_162),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_47),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_139),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_60),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_148),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_68),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_16),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_56),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_18),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_81),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_7),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_17),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_25),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_46),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_7),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_70),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_26),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_113),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_98),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_59),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_38),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_115),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_6),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_20),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_41),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_121),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_0),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_112),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_176),
.Y(n_343)
);

BUFx2_ASAP7_75t_SL g344 ( 
.A(n_193),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_178),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_243),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_279),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_243),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_180),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_182),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_243),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_243),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_282),
.B(n_0),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_184),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_243),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_185),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_243),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_176),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_186),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_232),
.B(n_1),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_175),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_188),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_279),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_179),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_243),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_243),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_243),
.Y(n_367)
);

XNOR2x1_ASAP7_75t_L g368 ( 
.A(n_173),
.B(n_2),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_292),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_200),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_292),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_203),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_211),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_205),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_292),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_211),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_309),
.B(n_193),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_292),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_292),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_206),
.Y(n_380)
);

NOR2xp67_ASAP7_75t_L g381 ( 
.A(n_282),
.B(n_4),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_L g382 ( 
.A(n_282),
.B(n_6),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_246),
.B(n_9),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_292),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_208),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_207),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_221),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_282),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_228),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_246),
.B(n_11),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_204),
.B(n_11),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_298),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_298),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_209),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_204),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_218),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_222),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_224),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_285),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_237),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_217),
.A2(n_19),
.B(n_21),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_212),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_212),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_223),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_223),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_230),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_230),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_231),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_231),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_174),
.B(n_22),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_260),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_240),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_285),
.B(n_22),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_229),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_189),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_235),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_236),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_236),
.Y(n_420)
);

CKINVDCx14_ASAP7_75t_R g421 ( 
.A(n_276),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_238),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_238),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_239),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_239),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_198),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_242),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_262),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_250),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_250),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_369),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_383),
.B(n_247),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_344),
.B(n_252),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_346),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_382),
.B(n_210),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_347),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_371),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_348),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_368),
.A2(n_286),
.B1(n_283),
.B2(n_322),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_351),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_344),
.B(n_198),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_375),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_351),
.Y(n_448)
);

INVx6_ASAP7_75t_L g449 ( 
.A(n_414),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_391),
.B(n_210),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_426),
.B(n_306),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_377),
.B(n_390),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_352),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_363),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_378),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_378),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_L g458 ( 
.A(n_391),
.B(n_241),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_415),
.B(n_210),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_352),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_415),
.B(n_219),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_395),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_414),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_368),
.B(n_417),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_382),
.B(n_219),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_388),
.B(n_219),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_355),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_355),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_384),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_388),
.B(n_274),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_357),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_357),
.Y(n_474)
);

OR2x6_ASAP7_75t_L g475 ( 
.A(n_403),
.B(n_274),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_365),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_404),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_395),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_365),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_404),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_400),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_353),
.B(n_274),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_366),
.B(n_259),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_366),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_367),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_403),
.A2(n_226),
.B(n_217),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_367),
.Y(n_487)
);

INVx6_ASAP7_75t_L g488 ( 
.A(n_426),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_400),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_343),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_421),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_392),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_381),
.B(n_342),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_392),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_393),
.B(n_342),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_360),
.B(n_306),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_393),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_396),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_396),
.B(n_342),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_405),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_402),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_345),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_405),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_349),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_406),
.B(n_240),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_406),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_435),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_435),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_432),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_435),
.Y(n_511)
);

INVx8_ASAP7_75t_L g512 ( 
.A(n_475),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_432),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_432),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_487),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_442),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_478),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_445),
.B(n_350),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_435),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_487),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_435),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_434),
.B(n_354),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_SL g524 ( 
.A(n_451),
.B(n_241),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_435),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_445),
.B(n_356),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_442),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_452),
.B(n_483),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_442),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_434),
.B(n_359),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_435),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_452),
.B(n_407),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_449),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_491),
.B(n_362),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_442),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_444),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_485),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_491),
.B(n_370),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_435),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_449),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_505),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_438),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_471),
.B(n_407),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_444),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_485),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_438),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_491),
.B(n_372),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_438),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_444),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_438),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_475),
.A2(n_412),
.B1(n_310),
.B2(n_291),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_496),
.B(n_374),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_443),
.B(n_361),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_444),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_496),
.B(n_380),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_503),
.B(n_386),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_453),
.Y(n_558)
);

CKINVDCx6p67_ASAP7_75t_R g559 ( 
.A(n_451),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_471),
.B(n_450),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_478),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_453),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_433),
.B(n_394),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_453),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_485),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_449),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_483),
.B(n_433),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_449),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_L g569 ( 
.A1(n_462),
.A2(n_311),
.B1(n_358),
.B2(n_422),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_471),
.B(n_408),
.Y(n_570)
);

AOI21x1_ASAP7_75t_L g571 ( 
.A1(n_431),
.A2(n_455),
.B(n_436),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_482),
.B(n_397),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_481),
.B(n_398),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_450),
.B(n_408),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_485),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_453),
.Y(n_576)
);

NAND3xp33_ASAP7_75t_L g577 ( 
.A(n_462),
.B(n_416),
.C(n_399),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_482),
.B(n_418),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_503),
.B(n_427),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_468),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_438),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_503),
.B(n_201),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_482),
.B(n_249),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_468),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_468),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_450),
.B(n_409),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_482),
.B(n_249),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_468),
.Y(n_588)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_481),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_449),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_489),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_459),
.B(n_409),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_438),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_464),
.B(n_364),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_482),
.B(n_183),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_469),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

XOR2x2_ASAP7_75t_SL g598 ( 
.A(n_443),
.B(n_310),
.Y(n_598)
);

OAI22x1_ASAP7_75t_L g599 ( 
.A1(n_464),
.A2(n_291),
.B1(n_303),
.B2(n_316),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_469),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_503),
.B(n_201),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_459),
.B(n_410),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_469),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_469),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_438),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_472),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_472),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_472),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_449),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_488),
.B(n_503),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_475),
.A2(n_316),
.B1(n_303),
.B2(n_325),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_472),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_449),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_476),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_505),
.Y(n_615)
);

BUFx8_ASAP7_75t_SL g616 ( 
.A(n_439),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_454),
.B(n_385),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_475),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_454),
.B(n_387),
.Y(n_619)
);

AND2x6_ASAP7_75t_L g620 ( 
.A(n_437),
.B(n_226),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_476),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_476),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_475),
.A2(n_325),
.B1(n_337),
.B2(n_253),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_476),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_484),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_458),
.A2(n_225),
.B1(n_251),
.B2(n_267),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_484),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_484),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_489),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_484),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_439),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_440),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_459),
.B(n_410),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_448),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_490),
.B(n_389),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_448),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_463),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_440),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_439),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_482),
.B(n_263),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_490),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_441),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_488),
.A2(n_315),
.B1(n_271),
.B2(n_299),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_448),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_467),
.B(n_174),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_441),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_448),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_448),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_448),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_488),
.Y(n_650)
);

XNOR2x2_ASAP7_75t_R g651 ( 
.A(n_464),
.B(n_401),
.Y(n_651)
);

AND2x6_ASAP7_75t_L g652 ( 
.A(n_437),
.B(n_227),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_446),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_448),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_461),
.B(n_411),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_458),
.B(n_376),
.C(n_373),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_463),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_475),
.A2(n_253),
.B1(n_337),
.B2(n_287),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_493),
.B(n_266),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_493),
.B(n_268),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_528),
.B(n_488),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_567),
.B(n_461),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_563),
.B(n_461),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_560),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_523),
.B(n_437),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_530),
.B(n_437),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_516),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_516),
.Y(n_668)
);

NAND3xp33_ASAP7_75t_L g669 ( 
.A(n_556),
.B(n_506),
.C(n_493),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_560),
.B(n_437),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_533),
.B(n_437),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_574),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_519),
.B(n_488),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_533),
.B(n_466),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_526),
.B(n_488),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_573),
.B(n_488),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_618),
.B(n_466),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_521),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_574),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_571),
.Y(n_680)
);

CKINVDCx16_ASAP7_75t_R g681 ( 
.A(n_589),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_631),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_521),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_573),
.B(n_413),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_658),
.B(n_466),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_586),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_531),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_571),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_586),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_611),
.B(n_466),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_592),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_650),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_592),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_602),
.Y(n_694)
);

AND2x2_ASAP7_75t_SL g695 ( 
.A(n_552),
.B(n_227),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_602),
.B(n_467),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_623),
.B(n_466),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_531),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_645),
.A2(n_475),
.B1(n_466),
.B2(n_493),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_618),
.B(n_650),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_633),
.B(n_467),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_639),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_538),
.B(n_493),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_633),
.B(n_467),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_655),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_655),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_538),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_544),
.B(n_467),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_518),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_546),
.B(n_493),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_546),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_565),
.B(n_448),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_512),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_565),
.B(n_460),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_575),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_618),
.B(n_463),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_577),
.B(n_553),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_575),
.B(n_460),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_632),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_595),
.B(n_460),
.Y(n_720)
);

AND2x2_ASAP7_75t_SL g721 ( 
.A(n_645),
.B(n_257),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_632),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_544),
.B(n_467),
.Y(n_723)
);

INVx8_ASAP7_75t_L g724 ( 
.A(n_512),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_570),
.B(n_460),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_638),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_520),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_638),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_570),
.B(n_642),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_618),
.B(n_257),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_642),
.B(n_460),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_646),
.B(n_460),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_646),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_520),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_653),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_653),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_583),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_618),
.B(n_645),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_645),
.B(n_572),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_578),
.B(n_460),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_579),
.B(n_460),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_524),
.A2(n_428),
.B1(n_317),
.B2(n_195),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_587),
.B(n_474),
.Y(n_743)
);

OAI22xp33_ASAP7_75t_SL g744 ( 
.A1(n_582),
.A2(n_284),
.B1(n_288),
.B2(n_281),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_620),
.A2(n_486),
.B1(n_287),
.B2(n_312),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_618),
.B(n_463),
.Y(n_746)
);

NOR2xp67_ASAP7_75t_L g747 ( 
.A(n_643),
.B(n_463),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_641),
.B(n_265),
.Y(n_748)
);

OAI221xp5_ASAP7_75t_L g749 ( 
.A1(n_626),
.A2(n_477),
.B1(n_480),
.B2(n_500),
.C(n_258),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_576),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_L g751 ( 
.A(n_512),
.B(n_177),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_640),
.B(n_474),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_L g753 ( 
.A(n_512),
.B(n_177),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_589),
.B(n_506),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_635),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_659),
.B(n_474),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_660),
.B(n_508),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_518),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_SL g759 ( 
.A1(n_598),
.A2(n_326),
.B1(n_334),
.B2(n_201),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_508),
.B(n_474),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_542),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_508),
.B(n_474),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_512),
.B(n_463),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_576),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_580),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_580),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_641),
.B(n_495),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_508),
.B(n_474),
.Y(n_768)
);

BUFx5_ASAP7_75t_L g769 ( 
.A(n_620),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_617),
.B(n_506),
.C(n_499),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_561),
.B(n_181),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_511),
.B(n_474),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_585),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_511),
.B(n_474),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_647),
.B(n_463),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_620),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_561),
.B(n_187),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_510),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_511),
.B(n_479),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_647),
.B(n_463),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_522),
.B(n_479),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_610),
.A2(n_559),
.B1(n_557),
.B2(n_591),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_620),
.B(n_191),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_510),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_534),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_656),
.A2(n_486),
.B(n_507),
.C(n_281),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_559),
.A2(n_269),
.B1(n_270),
.B2(n_302),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_585),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_591),
.B(n_190),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_596),
.Y(n_790)
);

NAND2x1p5_ASAP7_75t_L g791 ( 
.A(n_534),
.B(n_486),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_513),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_522),
.B(n_479),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_596),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_513),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_647),
.B(n_463),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_513),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_639),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_514),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_629),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_649),
.B(n_479),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_514),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_626),
.A2(n_507),
.B(n_284),
.C(n_312),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_649),
.B(n_479),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_514),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_522),
.B(n_479),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_620),
.A2(n_652),
.B1(n_604),
.B2(n_606),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_603),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_601),
.B(n_192),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_620),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_603),
.A2(n_507),
.B(n_436),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_515),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_543),
.B(n_507),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_543),
.B(n_507),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_543),
.B(n_446),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_604),
.Y(n_816)
);

AOI221xp5_ASAP7_75t_L g817 ( 
.A1(n_569),
.A2(n_278),
.B1(n_294),
.B2(n_293),
.C(n_290),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_607),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_649),
.B(n_273),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_543),
.B(n_447),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_515),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_620),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_515),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_527),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_535),
.B(n_539),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_612),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_654),
.B(n_295),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_786),
.A2(n_614),
.B(n_612),
.Y(n_828)
);

OAI321xp33_ASAP7_75t_L g829 ( 
.A1(n_749),
.A2(n_619),
.A3(n_598),
.B1(n_548),
.B2(n_234),
.C(n_194),
.Y(n_829)
);

O2A1O1Ixp5_ASAP7_75t_L g830 ( 
.A1(n_661),
.A2(n_654),
.B(n_581),
.C(n_593),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_663),
.B(n_610),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_723),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_755),
.B(n_599),
.Y(n_833)
);

BUFx12f_ASAP7_75t_L g834 ( 
.A(n_761),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_662),
.B(n_615),
.Y(n_835)
);

OAI21xp33_ASAP7_75t_L g836 ( 
.A1(n_759),
.A2(n_599),
.B(n_202),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_667),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_671),
.B(n_610),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_707),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_769),
.B(n_615),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_674),
.B(n_610),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_665),
.A2(n_541),
.B(n_534),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_798),
.B(n_615),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_798),
.Y(n_844)
);

O2A1O1Ixp5_ASAP7_75t_L g845 ( 
.A1(n_819),
.A2(n_654),
.B(n_593),
.C(n_605),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_664),
.A2(n_258),
.B(n_304),
.C(n_288),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_666),
.A2(n_566),
.B(n_541),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_707),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_754),
.B(n_615),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_717),
.A2(n_610),
.B1(n_652),
.B2(n_620),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_767),
.B(n_554),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_691),
.B(n_652),
.Y(n_852)
);

O2A1O1Ixp5_ASAP7_75t_L g853 ( 
.A1(n_819),
.A2(n_593),
.B(n_549),
.C(n_634),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_740),
.A2(n_566),
.B(n_541),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_786),
.A2(n_624),
.B(n_621),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_691),
.B(n_652),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_702),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_667),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_803),
.A2(n_214),
.B(n_304),
.C(n_216),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_670),
.A2(n_628),
.B(n_627),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_705),
.B(n_652),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_725),
.A2(n_628),
.B(n_627),
.Y(n_862)
);

AOI21x1_ASAP7_75t_L g863 ( 
.A1(n_677),
.A2(n_630),
.B(n_545),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_721),
.A2(n_652),
.B1(n_581),
.B2(n_593),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_705),
.B(n_652),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_707),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_769),
.B(n_549),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_713),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_754),
.B(n_709),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_709),
.B(n_554),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_739),
.A2(n_568),
.B(n_566),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_720),
.A2(n_590),
.B(n_568),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_682),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_743),
.A2(n_590),
.B(n_568),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_695),
.A2(n_256),
.B(n_277),
.C(n_264),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_758),
.B(n_549),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_723),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_758),
.B(n_748),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_677),
.A2(n_609),
.B(n_590),
.Y(n_879)
);

O2A1O1Ixp5_ASAP7_75t_L g880 ( 
.A1(n_827),
.A2(n_549),
.B(n_581),
.C(n_605),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_825),
.B(n_581),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_713),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_696),
.B(n_605),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_729),
.A2(n_608),
.B(n_527),
.C(n_529),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_752),
.A2(n_613),
.B(n_609),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_668),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_756),
.A2(n_757),
.B(n_688),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_680),
.A2(n_613),
.B(n_609),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_701),
.B(n_605),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_701),
.B(n_634),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_769),
.B(n_634),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_680),
.A2(n_613),
.B(n_532),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_668),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_688),
.A2(n_532),
.B(n_509),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_704),
.B(n_634),
.Y(n_895)
);

NOR2x1_ASAP7_75t_L g896 ( 
.A(n_692),
.B(n_191),
.Y(n_896)
);

O2A1O1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_672),
.A2(n_584),
.B(n_527),
.C(n_529),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_678),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_678),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_685),
.A2(n_532),
.B(n_509),
.Y(n_900)
);

O2A1O1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_679),
.A2(n_529),
.B(n_537),
.C(n_536),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_723),
.Y(n_902)
);

NOR3xp33_ASAP7_75t_L g903 ( 
.A(n_684),
.B(n_499),
.C(n_495),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_713),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_683),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_704),
.B(n_517),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_737),
.A2(n_669),
.B(n_708),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_695),
.A2(n_277),
.B(n_196),
.C(n_197),
.Y(n_908)
);

OAI321xp33_ASAP7_75t_L g909 ( 
.A1(n_817),
.A2(n_809),
.A3(n_742),
.B1(n_771),
.B2(n_789),
.C(n_777),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_676),
.B(n_509),
.Y(n_910)
);

INVx4_ASAP7_75t_L g911 ( 
.A(n_713),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_683),
.Y(n_912)
);

AOI21x1_ASAP7_75t_L g913 ( 
.A1(n_801),
.A2(n_600),
.B(n_517),
.Y(n_913)
);

AOI21x1_ASAP7_75t_L g914 ( 
.A1(n_804),
.A2(n_600),
.B(n_537),
.Y(n_914)
);

NOR2x1_ASAP7_75t_R g915 ( 
.A(n_761),
.B(n_651),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_741),
.A2(n_532),
.B(n_509),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_687),
.Y(n_917)
);

NOR2x1p5_ASAP7_75t_SL g918 ( 
.A(n_769),
.B(n_536),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_708),
.B(n_536),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_767),
.B(n_594),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_686),
.A2(n_689),
.B(n_694),
.C(n_693),
.Y(n_921)
);

NOR3xp33_ASAP7_75t_L g922 ( 
.A(n_800),
.B(n_499),
.C(n_495),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_800),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_706),
.A2(n_550),
.B(n_555),
.C(n_625),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_713),
.B(n_692),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_698),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_719),
.B(n_477),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_703),
.A2(n_555),
.B(n_550),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_698),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_769),
.B(n_520),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_770),
.B(n_594),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_710),
.A2(n_551),
.B(n_540),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_681),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_699),
.A2(n_197),
.B1(n_256),
.B2(n_248),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_722),
.A2(n_234),
.B(n_214),
.C(n_264),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_733),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_745),
.A2(n_551),
.B(n_540),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_726),
.B(n_480),
.Y(n_938)
);

AOI21xp33_ASAP7_75t_L g939 ( 
.A1(n_673),
.A2(n_196),
.B(n_194),
.Y(n_939)
);

AO21x2_ASAP7_75t_L g940 ( 
.A1(n_747),
.A2(n_248),
.B(n_216),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_738),
.A2(n_551),
.B(n_540),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_733),
.Y(n_942)
);

AOI21xp33_ASAP7_75t_L g943 ( 
.A1(n_675),
.A2(n_213),
.B(n_199),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_728),
.B(n_550),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_736),
.B(n_555),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_738),
.A2(n_551),
.B(n_540),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_700),
.A2(n_597),
.B(n_637),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_735),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_700),
.A2(n_597),
.B(n_637),
.Y(n_949)
);

NAND3xp33_ASAP7_75t_L g950 ( 
.A(n_787),
.B(n_220),
.C(n_215),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_735),
.B(n_558),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_721),
.B(n_711),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_690),
.A2(n_562),
.B(n_558),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_715),
.B(n_562),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_697),
.A2(n_622),
.B1(n_564),
.B2(n_584),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_782),
.B(n_597),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_765),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_804),
.A2(n_625),
.B(n_584),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_765),
.B(n_564),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_766),
.B(n_564),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_766),
.B(n_597),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_807),
.A2(n_657),
.B(n_637),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_811),
.A2(n_657),
.B(n_648),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_763),
.A2(n_657),
.B(n_648),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_785),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_750),
.B(n_764),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_773),
.B(n_588),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_744),
.A2(n_625),
.B(n_622),
.C(n_608),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_776),
.A2(n_608),
.B1(n_588),
.B2(n_622),
.Y(n_969)
);

OAI21xp33_ASAP7_75t_L g970 ( 
.A1(n_788),
.A2(n_301),
.B(n_323),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_751),
.A2(n_588),
.B1(n_340),
.B2(n_320),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_810),
.A2(n_648),
.B(n_644),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_769),
.B(n_810),
.Y(n_973)
);

AOI21x1_ASAP7_75t_L g974 ( 
.A1(n_716),
.A2(n_465),
.B(n_431),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_730),
.A2(n_648),
.B(n_644),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_790),
.B(n_520),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_769),
.B(n_520),
.Y(n_977)
);

NOR2xp67_ASAP7_75t_L g978 ( 
.A(n_731),
.B(n_732),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_794),
.B(n_525),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_785),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_724),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_808),
.B(n_816),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_818),
.B(n_500),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_712),
.A2(n_431),
.B(n_455),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_751),
.A2(n_456),
.B(n_470),
.C(n_473),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_SL g986 ( 
.A1(n_813),
.A2(n_425),
.B(n_430),
.C(n_411),
.Y(n_986)
);

NOR2x1_ASAP7_75t_L g987 ( 
.A(n_776),
.B(n_447),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_822),
.A2(n_644),
.B1(n_636),
.B2(n_547),
.Y(n_988)
);

CKINVDCx10_ASAP7_75t_R g989 ( 
.A(n_753),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_791),
.A2(n_636),
.B(n_547),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_826),
.B(n_616),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_724),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_822),
.B(n_276),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_SL g994 ( 
.A1(n_814),
.A2(n_425),
.B(n_430),
.C(n_419),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_778),
.B(n_525),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_714),
.B(n_419),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_784),
.B(n_525),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_784),
.B(n_276),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_792),
.B(n_525),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_724),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_795),
.B(n_525),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_795),
.B(n_276),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_753),
.A2(n_420),
.B(n_423),
.C(n_424),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_724),
.A2(n_783),
.B(n_718),
.C(n_821),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_791),
.A2(n_636),
.B(n_547),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_909),
.A2(n_783),
.B(n_815),
.C(n_820),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_838),
.A2(n_785),
.B(n_734),
.Y(n_1007)
);

INVx6_ASAP7_75t_L g1008 ( 
.A(n_834),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_878),
.B(n_797),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_878),
.B(n_835),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_835),
.B(n_799),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_841),
.A2(n_785),
.B(n_734),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_873),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_937),
.A2(n_785),
.B(n_734),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_881),
.B(n_799),
.Y(n_1015)
);

NOR2x1_ASAP7_75t_R g1016 ( 
.A(n_933),
.B(n_851),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_952),
.A2(n_727),
.B1(n_779),
.B2(n_760),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_857),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_957),
.Y(n_1019)
);

OR2x6_ASAP7_75t_SL g1020 ( 
.A(n_950),
.B(n_233),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_843),
.B(n_727),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_920),
.B(n_420),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_829),
.A2(n_921),
.B(n_939),
.C(n_956),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_843),
.B(n_727),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_905),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_870),
.B(n_423),
.Y(n_1026)
);

O2A1O1Ixp5_ASAP7_75t_SL g1027 ( 
.A1(n_943),
.A2(n_429),
.B(n_424),
.C(n_473),
.Y(n_1027)
);

OAI21xp33_ASAP7_75t_SL g1028 ( 
.A1(n_850),
.A2(n_746),
.B(n_716),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_956),
.A2(n_881),
.B(n_907),
.C(n_903),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_938),
.B(n_802),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_870),
.B(n_429),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_857),
.Y(n_1032)
);

OAI21xp33_ASAP7_75t_L g1033 ( 
.A1(n_869),
.A2(n_305),
.B(n_341),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_844),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_903),
.A2(n_746),
.B1(n_775),
.B2(n_780),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_869),
.B(n_244),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_849),
.A2(n_775),
.B1(n_780),
.B2(n_796),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_910),
.B(n_802),
.Y(n_1038)
);

O2A1O1Ixp5_ASAP7_75t_L g1039 ( 
.A1(n_910),
.A2(n_768),
.B(n_762),
.C(n_772),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_868),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_831),
.A2(n_806),
.B(n_781),
.Y(n_1041)
);

AO32x1_ASAP7_75t_L g1042 ( 
.A1(n_934),
.A2(n_824),
.A3(n_823),
.B1(n_821),
.B2(n_812),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_844),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_858),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_SL g1045 ( 
.A(n_915),
.B(n_201),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_948),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_R g1047 ( 
.A(n_989),
.B(n_774),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_849),
.A2(n_793),
.B(n_823),
.C(n_812),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_922),
.B(n_805),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_887),
.A2(n_796),
.B(n_636),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_923),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_931),
.B(n_833),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_942),
.Y(n_1053)
);

INVx6_ASAP7_75t_L g1054 ( 
.A(n_868),
.Y(n_1054)
);

NOR2x1_ASAP7_75t_SL g1055 ( 
.A(n_868),
.B(n_824),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_961),
.A2(n_547),
.B(n_504),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_922),
.B(n_504),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_927),
.B(n_245),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_832),
.B(n_314),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_832),
.B(n_319),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_877),
.A2(n_324),
.B1(n_330),
.B2(n_332),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_877),
.B(n_333),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_902),
.B(n_336),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_875),
.A2(n_498),
.B(n_254),
.C(n_328),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_842),
.A2(n_436),
.B(n_455),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_993),
.B(n_280),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_836),
.A2(n_280),
.B1(n_498),
.B2(n_255),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_991),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_847),
.A2(n_916),
.B(n_973),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_875),
.A2(n_498),
.B(n_261),
.C(n_329),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_868),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_SL g1072 ( 
.A(n_991),
.B(n_275),
.C(n_272),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_973),
.A2(n_465),
.B(n_457),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_896),
.B(n_280),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_925),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_942),
.B(n_498),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_894),
.A2(n_465),
.B(n_457),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_936),
.B(n_470),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_858),
.A2(n_280),
.B1(n_321),
.B2(n_318),
.Y(n_1079)
);

BUFx12f_ASAP7_75t_L g1080 ( 
.A(n_925),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_839),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_998),
.B(n_335),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_882),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_837),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_930),
.A2(n_456),
.B(n_501),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_908),
.A2(n_331),
.B(n_296),
.C(n_297),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_882),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_893),
.A2(n_338),
.B1(n_300),
.B2(n_307),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1002),
.B(n_502),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_966),
.A2(n_289),
.B1(n_308),
.B2(n_313),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_930),
.A2(n_501),
.B(n_497),
.Y(n_1091)
);

AOI21x1_ASAP7_75t_L g1092 ( 
.A1(n_990),
.A2(n_502),
.B(n_501),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_908),
.A2(n_339),
.B(n_501),
.C(n_497),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_983),
.B(n_23),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_882),
.B(n_494),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_882),
.B(n_494),
.Y(n_1096)
);

NOR2xp67_ASAP7_75t_L g1097 ( 
.A(n_970),
.B(n_170),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_899),
.B(n_502),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_912),
.B(n_502),
.Y(n_1099)
);

NOR2xp67_ASAP7_75t_L g1100 ( 
.A(n_996),
.B(n_155),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_982),
.B(n_23),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_852),
.B(n_494),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_886),
.B(n_497),
.Y(n_1103)
);

INVxp67_ASAP7_75t_SL g1104 ( 
.A(n_904),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_828),
.A2(n_497),
.B(n_492),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_977),
.A2(n_1005),
.B(n_892),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_926),
.B(n_492),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_864),
.A2(n_492),
.B1(n_494),
.B2(n_154),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_883),
.B(n_24),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_898),
.B(n_492),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_856),
.B(n_494),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_977),
.A2(n_494),
.B(n_153),
.Y(n_1112)
);

CKINVDCx8_ASAP7_75t_R g1113 ( 
.A(n_904),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_871),
.A2(n_494),
.B(n_152),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_846),
.A2(n_24),
.B(n_27),
.C(n_29),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_917),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_848),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_932),
.A2(n_494),
.B(n_144),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_SL g1119 ( 
.A(n_911),
.B(n_992),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_R g1120 ( 
.A(n_981),
.B(n_1000),
.Y(n_1120)
);

INVx8_ASAP7_75t_L g1121 ( 
.A(n_904),
.Y(n_1121)
);

AO32x1_ASAP7_75t_L g1122 ( 
.A1(n_955),
.A2(n_29),
.A3(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_929),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_900),
.A2(n_133),
.B(n_126),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_861),
.B(n_119),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_889),
.B(n_32),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_846),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_866),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_944),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_904),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_945),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_865),
.A2(n_919),
.B1(n_906),
.B2(n_840),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_987),
.A2(n_118),
.B1(n_88),
.B2(n_86),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_954),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_890),
.B(n_35),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_913),
.A2(n_914),
.B(n_958),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_SL g1137 ( 
.A1(n_876),
.A2(n_82),
.B(n_80),
.C(n_75),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_965),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_840),
.A2(n_895),
.B1(n_1004),
.B2(n_911),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_855),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1004),
.A2(n_74),
.B1(n_69),
.B2(n_64),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_981),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_992),
.B(n_36),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_876),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_978),
.B(n_39),
.Y(n_1145)
);

BUFx4f_ASAP7_75t_SL g1146 ( 
.A(n_981),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_888),
.A2(n_885),
.B(n_879),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_854),
.A2(n_63),
.B(n_44),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_951),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_862),
.A2(n_43),
.B(n_44),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_860),
.A2(n_47),
.B(n_52),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1010),
.B(n_971),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1052),
.B(n_965),
.Y(n_1153)
);

CKINVDCx8_ASAP7_75t_R g1154 ( 
.A(n_1051),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1029),
.A2(n_859),
.A3(n_1003),
.B(n_935),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1092),
.A2(n_830),
.B(n_845),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1046),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1026),
.B(n_1000),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1019),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1034),
.B(n_1000),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_1113),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1014),
.A2(n_863),
.B(n_880),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1038),
.A2(n_872),
.B(n_874),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1031),
.B(n_959),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1022),
.B(n_1129),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1069),
.A2(n_941),
.B(n_946),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_SL g1167 ( 
.A1(n_1023),
.A2(n_891),
.B(n_867),
.C(n_979),
.Y(n_1167)
);

AO21x2_ASAP7_75t_L g1168 ( 
.A1(n_1147),
.A2(n_984),
.B(n_940),
.Y(n_1168)
);

AO31x2_ASAP7_75t_L g1169 ( 
.A1(n_1093),
.A2(n_969),
.A3(n_988),
.B(n_975),
.Y(n_1169)
);

AOI221xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1067),
.A2(n_924),
.B1(n_901),
.B2(n_897),
.C(n_968),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1082),
.B(n_1036),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1131),
.B(n_960),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1013),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1103),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1134),
.B(n_980),
.Y(n_1175)
);

OA21x2_ASAP7_75t_L g1176 ( 
.A1(n_1039),
.A2(n_853),
.B(n_928),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_SL g1177 ( 
.A1(n_1125),
.A2(n_891),
.B(n_867),
.C(n_976),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1009),
.B(n_980),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1106),
.A2(n_953),
.B(n_963),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1132),
.A2(n_949),
.B(n_947),
.Y(n_1180)
);

AO221x1_ASAP7_75t_L g1181 ( 
.A1(n_1141),
.A2(n_1000),
.B1(n_994),
.B2(n_986),
.C(n_940),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1006),
.A2(n_1028),
.B(n_1064),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1018),
.B(n_974),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1009),
.B(n_967),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1098),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1101),
.A2(n_884),
.B(n_918),
.C(n_985),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1011),
.A2(n_972),
.B(n_962),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1101),
.A2(n_964),
.B(n_999),
.C(n_997),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1015),
.A2(n_1001),
.B(n_995),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1094),
.B(n_986),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1070),
.A2(n_994),
.B(n_54),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1094),
.A2(n_52),
.B1(n_54),
.B2(n_57),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1149),
.B(n_57),
.Y(n_1193)
);

AOI221xp5_ASAP7_75t_L g1194 ( 
.A1(n_1140),
.A2(n_58),
.B1(n_59),
.B2(n_1151),
.C(n_1090),
.Y(n_1194)
);

AOI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1041),
.A2(n_1024),
.B(n_1021),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1035),
.A2(n_1037),
.B(n_1027),
.Y(n_1196)
);

CKINVDCx6p67_ASAP7_75t_R g1197 ( 
.A(n_1068),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_1043),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1018),
.B(n_1032),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1109),
.B(n_1126),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1058),
.B(n_1032),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_L g1202 ( 
.A(n_1150),
.B(n_1140),
.C(n_1072),
.Y(n_1202)
);

AOI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1007),
.A2(n_1012),
.B(n_1111),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1033),
.B(n_1088),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_SL g1205 ( 
.A(n_1016),
.B(n_1008),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_SL g1206 ( 
.A(n_1045),
.B(n_1079),
.C(n_1067),
.Y(n_1206)
);

BUFx10_ASAP7_75t_L g1207 ( 
.A(n_1008),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1066),
.A2(n_1144),
.B(n_1074),
.C(n_1115),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1099),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1075),
.B(n_1083),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1097),
.A2(n_1109),
.B1(n_1126),
.B2(n_1135),
.Y(n_1211)
);

AOI221x1_ASAP7_75t_L g1212 ( 
.A1(n_1148),
.A2(n_1108),
.B1(n_1114),
.B2(n_1118),
.C(n_1086),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1048),
.A2(n_1017),
.A3(n_1050),
.B(n_1056),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1135),
.A2(n_1062),
.B1(n_1059),
.B2(n_1063),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1065),
.A2(n_1091),
.B(n_1077),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1081),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1089),
.A2(n_1039),
.B(n_1119),
.Y(n_1217)
);

OAI22x1_ASAP7_75t_L g1218 ( 
.A1(n_1127),
.A2(n_1143),
.B1(n_1084),
.B2(n_1125),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1124),
.A2(n_1055),
.A3(n_1057),
.B(n_1145),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_SL g1220 ( 
.A1(n_1079),
.A2(n_1088),
.B(n_1133),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_SL g1221 ( 
.A1(n_1137),
.A2(n_1049),
.B(n_1060),
.C(n_1111),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1107),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1102),
.A2(n_1030),
.B(n_1104),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1146),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1081),
.B(n_1117),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1085),
.A2(n_1102),
.B(n_1073),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1047),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1112),
.A2(n_1042),
.A3(n_1078),
.B(n_1110),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1042),
.A2(n_1076),
.A3(n_1116),
.B(n_1025),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1104),
.A2(n_1100),
.B(n_1042),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1095),
.A2(n_1096),
.B(n_1137),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1121),
.A2(n_1105),
.B(n_1053),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1053),
.A2(n_1117),
.B1(n_1128),
.B2(n_1138),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1123),
.A2(n_1122),
.A3(n_1105),
.B(n_1020),
.Y(n_1234)
);

AOI221x1_ASAP7_75t_L g1235 ( 
.A1(n_1143),
.A2(n_1122),
.B1(n_1071),
.B2(n_1087),
.C(n_1040),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1128),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1061),
.B(n_1047),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1105),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1071),
.A2(n_1087),
.B(n_1072),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1142),
.B(n_1040),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1122),
.A2(n_1120),
.B(n_1080),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1040),
.A2(n_1130),
.A3(n_1054),
.B(n_1121),
.Y(n_1242)
);

OR2x6_ASAP7_75t_L g1243 ( 
.A(n_1121),
.B(n_1142),
.Y(n_1243)
);

AO21x2_ASAP7_75t_L g1244 ( 
.A1(n_1120),
.A2(n_1040),
.B(n_1130),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1130),
.A2(n_1142),
.B(n_1146),
.C(n_1054),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1130),
.B(n_1054),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1044),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1029),
.A2(n_1139),
.A3(n_1093),
.B(n_956),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1136),
.A2(n_1092),
.B(n_1014),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1026),
.B(n_1031),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1026),
.B(n_920),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1010),
.A2(n_909),
.B(n_755),
.C(n_1023),
.Y(n_1252)
);

OAI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1010),
.A2(n_496),
.B1(n_909),
.B2(n_755),
.Y(n_1253)
);

INVx8_ASAP7_75t_L g1254 ( 
.A(n_1121),
.Y(n_1254)
);

AOI211x1_ASAP7_75t_L g1255 ( 
.A1(n_1151),
.A2(n_836),
.B(n_749),
.C(n_1150),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1013),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1038),
.A2(n_666),
.B(n_665),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1136),
.A2(n_1092),
.B(n_1014),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1052),
.A2(n_684),
.B1(n_870),
.B2(n_619),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1136),
.A2(n_1092),
.B(n_1014),
.Y(n_1260)
);

AOI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1092),
.A2(n_1106),
.B(n_1139),
.Y(n_1261)
);

OR2x6_ASAP7_75t_L g1262 ( 
.A(n_1013),
.B(n_873),
.Y(n_1262)
);

OAI22x1_ASAP7_75t_L g1263 ( 
.A1(n_1052),
.A2(n_443),
.B1(n_554),
.B2(n_626),
.Y(n_1263)
);

BUFx2_ASAP7_75t_SL g1264 ( 
.A(n_1013),
.Y(n_1264)
);

AOI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1092),
.A2(n_1106),
.B(n_1139),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1038),
.A2(n_666),
.B(n_665),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1010),
.B(n_528),
.Y(n_1267)
);

CKINVDCx14_ASAP7_75t_R g1268 ( 
.A(n_1008),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1010),
.B(n_528),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1023),
.A2(n_909),
.B(n_717),
.C(n_556),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1029),
.A2(n_1139),
.A3(n_1093),
.B(n_956),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1038),
.A2(n_666),
.B(n_665),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1038),
.A2(n_666),
.B(n_665),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1038),
.A2(n_666),
.B(n_665),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1010),
.A2(n_909),
.B(n_755),
.C(n_1023),
.Y(n_1275)
);

INVx8_ASAP7_75t_L g1276 ( 
.A(n_1121),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1023),
.A2(n_1029),
.B(n_909),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1136),
.A2(n_1092),
.B(n_1014),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1051),
.B(n_615),
.Y(n_1279)
);

INVx3_ASAP7_75t_SL g1280 ( 
.A(n_1051),
.Y(n_1280)
);

AO32x2_ASAP7_75t_L g1281 ( 
.A1(n_1139),
.A2(n_1144),
.A3(n_934),
.B1(n_1132),
.B2(n_1141),
.Y(n_1281)
);

AOI221x1_ASAP7_75t_L g1282 ( 
.A1(n_1151),
.A2(n_1150),
.B1(n_1023),
.B2(n_1029),
.C(n_939),
.Y(n_1282)
);

OA22x2_ASAP7_75t_L g1283 ( 
.A1(n_1018),
.A2(n_443),
.B1(n_626),
.B2(n_554),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1010),
.B(n_528),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1146),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1038),
.A2(n_666),
.B(n_665),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1010),
.A2(n_835),
.B1(n_663),
.B2(n_1029),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1010),
.A2(n_835),
.B1(n_663),
.B2(n_1029),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1010),
.B(n_755),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1023),
.A2(n_1029),
.B(n_909),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1026),
.B(n_1031),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1038),
.A2(n_666),
.B(n_665),
.Y(n_1292)
);

INVxp67_ASAP7_75t_SL g1293 ( 
.A(n_1018),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1013),
.Y(n_1294)
);

AOI22x1_ASAP7_75t_L g1295 ( 
.A1(n_1151),
.A2(n_1150),
.B1(n_1118),
.B2(n_1127),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1013),
.Y(n_1296)
);

OAI22x1_ASAP7_75t_L g1297 ( 
.A1(n_1052),
.A2(n_443),
.B1(n_554),
.B2(n_626),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1038),
.A2(n_666),
.B(n_665),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1026),
.B(n_920),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1038),
.A2(n_666),
.B(n_665),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1013),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1206),
.A2(n_1194),
.B1(n_1202),
.B2(n_1290),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1259),
.A2(n_1250),
.B1(n_1291),
.B2(n_1220),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1161),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1161),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1251),
.B(n_1299),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1277),
.A2(n_1204),
.B1(n_1283),
.B2(n_1200),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1253),
.A2(n_1152),
.B1(n_1211),
.B2(n_1297),
.Y(n_1308)
);

AO22x1_ASAP7_75t_L g1309 ( 
.A1(n_1289),
.A2(n_1165),
.B1(n_1280),
.B2(n_1267),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1295),
.A2(n_1171),
.B1(n_1182),
.B2(n_1237),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1287),
.A2(n_1288),
.B1(n_1205),
.B2(n_1191),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1262),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1269),
.A2(n_1284),
.B1(n_1270),
.B2(n_1164),
.Y(n_1313)
);

BUFx4_ASAP7_75t_R g1314 ( 
.A(n_1207),
.Y(n_1314)
);

BUFx10_ASAP7_75t_L g1315 ( 
.A(n_1173),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1201),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_SL g1317 ( 
.A1(n_1181),
.A2(n_1227),
.B1(n_1196),
.B2(n_1268),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1241),
.A2(n_1190),
.B1(n_1293),
.B2(n_1192),
.Y(n_1318)
);

CKINVDCx11_ASAP7_75t_R g1319 ( 
.A(n_1154),
.Y(n_1319)
);

INVx6_ASAP7_75t_L g1320 ( 
.A(n_1207),
.Y(n_1320)
);

INVx8_ASAP7_75t_L g1321 ( 
.A(n_1254),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1247),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1264),
.A2(n_1153),
.B1(n_1161),
.B2(n_1301),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1262),
.Y(n_1324)
);

AOI21xp33_ASAP7_75t_L g1325 ( 
.A1(n_1252),
.A2(n_1275),
.B(n_1208),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1263),
.A2(n_1158),
.B1(n_1218),
.B2(n_1214),
.Y(n_1326)
);

INVx6_ASAP7_75t_L g1327 ( 
.A(n_1254),
.Y(n_1327)
);

BUFx2_ASAP7_75t_SL g1328 ( 
.A(n_1224),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1216),
.A2(n_1256),
.B1(n_1296),
.B2(n_1294),
.Y(n_1329)
);

OAI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1282),
.A2(n_1197),
.B1(n_1193),
.B2(n_1279),
.Y(n_1330)
);

INVx4_ASAP7_75t_L g1331 ( 
.A(n_1276),
.Y(n_1331)
);

INVx4_ASAP7_75t_L g1332 ( 
.A(n_1276),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1225),
.Y(n_1333)
);

OAI21xp33_ASAP7_75t_L g1334 ( 
.A1(n_1199),
.A2(n_1172),
.B(n_1184),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1236),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1174),
.A2(n_1198),
.B1(n_1239),
.B2(n_1183),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1224),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1240),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1255),
.A2(n_1174),
.B1(n_1157),
.B2(n_1178),
.Y(n_1339)
);

BUFx8_ASAP7_75t_L g1340 ( 
.A(n_1210),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1185),
.B(n_1209),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1185),
.A2(n_1209),
.B1(n_1222),
.B2(n_1233),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1229),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1175),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1210),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1222),
.A2(n_1160),
.B1(n_1285),
.B2(n_1217),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1160),
.Y(n_1347)
);

BUFx4f_ASAP7_75t_SL g1348 ( 
.A(n_1240),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1229),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1246),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1244),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1168),
.A2(n_1223),
.B1(n_1180),
.B2(n_1232),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1244),
.Y(n_1353)
);

INVx8_ASAP7_75t_L g1354 ( 
.A(n_1243),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1243),
.Y(n_1355)
);

INVx8_ASAP7_75t_L g1356 ( 
.A(n_1242),
.Y(n_1356)
);

INVx6_ASAP7_75t_L g1357 ( 
.A(n_1245),
.Y(n_1357)
);

OAI21xp33_ASAP7_75t_L g1358 ( 
.A1(n_1186),
.A2(n_1188),
.B(n_1195),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1234),
.B(n_1271),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1238),
.Y(n_1360)
);

CKINVDCx11_ASAP7_75t_R g1361 ( 
.A(n_1238),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1168),
.A2(n_1187),
.B1(n_1298),
.B2(n_1292),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1234),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1234),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1230),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1155),
.Y(n_1366)
);

INVx6_ASAP7_75t_L g1367 ( 
.A(n_1167),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1257),
.A2(n_1300),
.B1(n_1266),
.B2(n_1286),
.Y(n_1368)
);

INVx6_ASAP7_75t_L g1369 ( 
.A(n_1221),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1155),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1272),
.A2(n_1274),
.B(n_1273),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1231),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_SL g1373 ( 
.A1(n_1212),
.A2(n_1235),
.B(n_1179),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1163),
.A2(n_1166),
.B1(n_1176),
.B2(n_1189),
.Y(n_1374)
);

INVx6_ASAP7_75t_L g1375 ( 
.A(n_1177),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1155),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1219),
.Y(n_1377)
);

OAI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1281),
.A2(n_1203),
.B1(n_1261),
.B2(n_1265),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1176),
.A2(n_1226),
.B1(n_1215),
.B2(n_1162),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1219),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1281),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1249),
.A2(n_1278),
.B1(n_1260),
.B2(n_1258),
.Y(n_1382)
);

INVx8_ASAP7_75t_L g1383 ( 
.A(n_1219),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1281),
.A2(n_1271),
.B1(n_1248),
.B2(n_1170),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1248),
.B(n_1271),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1248),
.B(n_1213),
.Y(n_1386)
);

BUFx2_ASAP7_75t_SL g1387 ( 
.A(n_1213),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1213),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1169),
.A2(n_1140),
.B1(n_1200),
.B2(n_1211),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1156),
.A2(n_1206),
.B1(n_1194),
.B2(n_1202),
.Y(n_1390)
);

CKINVDCx8_ASAP7_75t_R g1391 ( 
.A(n_1228),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1169),
.A2(n_684),
.B1(n_1259),
.B2(n_364),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1169),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1228),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1220),
.A2(n_759),
.B(n_1206),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1257),
.A2(n_1272),
.B(n_1266),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1200),
.A2(n_1140),
.B1(n_1211),
.B2(n_1267),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1283),
.A2(n_496),
.B1(n_1290),
.B2(n_1277),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1200),
.A2(n_1140),
.B1(n_1211),
.B2(n_1267),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1154),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1159),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1301),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_SL g1403 ( 
.A1(n_1283),
.A2(n_1297),
.B1(n_1263),
.B2(n_594),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1206),
.A2(n_1194),
.B1(n_1202),
.B2(n_1277),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1250),
.B(n_1291),
.Y(n_1405)
);

INVx4_ASAP7_75t_SL g1406 ( 
.A(n_1242),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1259),
.A2(n_496),
.B1(n_1200),
.B2(n_1211),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1200),
.A2(n_1140),
.B1(n_1211),
.B2(n_1267),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1259),
.A2(n_684),
.B1(n_364),
.B2(n_385),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1283),
.A2(n_496),
.B1(n_1290),
.B2(n_1277),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1161),
.Y(n_1411)
);

BUFx10_ASAP7_75t_L g1412 ( 
.A(n_1173),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1262),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1262),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1259),
.A2(n_684),
.B1(n_364),
.B2(n_385),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1262),
.Y(n_1416)
);

OAI21xp33_ASAP7_75t_L g1417 ( 
.A1(n_1200),
.A2(n_496),
.B(n_1211),
.Y(n_1417)
);

INVx6_ASAP7_75t_L g1418 ( 
.A(n_1207),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1283),
.A2(n_496),
.B1(n_1290),
.B2(n_1277),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1259),
.A2(n_684),
.B1(n_364),
.B2(n_385),
.Y(n_1420)
);

OAI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1200),
.A2(n_496),
.B1(n_1211),
.B2(n_1010),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1262),
.Y(n_1422)
);

INVx6_ASAP7_75t_L g1423 ( 
.A(n_1207),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1220),
.A2(n_759),
.B(n_1206),
.Y(n_1424)
);

OAI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1259),
.A2(n_496),
.B1(n_1200),
.B2(n_1211),
.Y(n_1425)
);

BUFx12f_ASAP7_75t_L g1426 ( 
.A(n_1207),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1200),
.A2(n_1140),
.B1(n_1211),
.B2(n_1267),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1360),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1366),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1379),
.A2(n_1382),
.B(n_1396),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1370),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1351),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1359),
.B(n_1381),
.Y(n_1433)
);

INVxp67_ASAP7_75t_L g1434 ( 
.A(n_1306),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1376),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_SL g1436 ( 
.A1(n_1403),
.A2(n_1421),
.B1(n_1399),
.B2(n_1397),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_SL g1437 ( 
.A1(n_1339),
.A2(n_1341),
.B(n_1325),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1405),
.Y(n_1438)
);

BUFx4f_ASAP7_75t_SL g1439 ( 
.A(n_1426),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1406),
.B(n_1393),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1356),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1381),
.B(n_1307),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1353),
.B(n_1388),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1343),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1381),
.B(n_1365),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1333),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1322),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1334),
.B(n_1333),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1377),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1385),
.B(n_1308),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1396),
.A2(n_1374),
.B(n_1371),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1409),
.B(n_1415),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1383),
.B(n_1387),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1349),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1417),
.B(n_1398),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1371),
.A2(n_1380),
.B(n_1352),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1363),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1319),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1385),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1394),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1386),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1386),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1320),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1320),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1410),
.A2(n_1419),
.B1(n_1424),
.B2(n_1395),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1378),
.A2(n_1373),
.B(n_1368),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1316),
.B(n_1350),
.Y(n_1467)
);

AO21x1_ASAP7_75t_SL g1468 ( 
.A1(n_1325),
.A2(n_1302),
.B(n_1404),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1340),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1339),
.Y(n_1470)
);

AO21x2_ASAP7_75t_L g1471 ( 
.A1(n_1373),
.A2(n_1368),
.B(n_1358),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1338),
.B(n_1372),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1384),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1372),
.A2(n_1362),
.B(n_1313),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1384),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1407),
.B(n_1425),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1320),
.Y(n_1477)
);

OAI211xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1395),
.A2(n_1424),
.B(n_1303),
.C(n_1326),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1389),
.A2(n_1392),
.B(n_1330),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1335),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1391),
.Y(n_1481)
);

A2O1A1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1311),
.A2(n_1408),
.B(n_1399),
.C(n_1397),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1316),
.B(n_1390),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1401),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1340),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1346),
.A2(n_1389),
.B(n_1341),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1375),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1313),
.A2(n_1342),
.B(n_1336),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1367),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1335),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1418),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1375),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1361),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1375),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1344),
.A2(n_1427),
.B(n_1408),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1310),
.B(n_1318),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1345),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1414),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1309),
.B(n_1427),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1369),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1364),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1318),
.Y(n_1502)
);

AO21x2_ASAP7_75t_L g1503 ( 
.A1(n_1420),
.A2(n_1317),
.B(n_1357),
.Y(n_1503)
);

OR2x6_ASAP7_75t_L g1504 ( 
.A(n_1354),
.B(n_1328),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1357),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1357),
.Y(n_1506)
);

OA21x2_ASAP7_75t_L g1507 ( 
.A1(n_1312),
.A2(n_1324),
.B(n_1422),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1354),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1354),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1355),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1413),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1348),
.A2(n_1337),
.B(n_1314),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1416),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1329),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1323),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1482),
.A2(n_1321),
.B(n_1305),
.C(n_1411),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1446),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1465),
.A2(n_1347),
.B1(n_1423),
.B2(n_1418),
.Y(n_1518)
);

AO32x2_ASAP7_75t_L g1519 ( 
.A1(n_1459),
.A2(n_1332),
.A3(n_1331),
.B1(n_1304),
.B2(n_1305),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1445),
.B(n_1402),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1507),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1480),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1433),
.B(n_1443),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1452),
.A2(n_1478),
.B1(n_1465),
.B2(n_1436),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1474),
.A2(n_1476),
.B(n_1488),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1496),
.A2(n_1423),
.B1(n_1418),
.B2(n_1411),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1499),
.B(n_1423),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1490),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1467),
.B(n_1315),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1496),
.A2(n_1321),
.B(n_1327),
.C(n_1400),
.Y(n_1530)
);

OAI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1488),
.A2(n_1331),
.B(n_1315),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1450),
.B(n_1412),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1447),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1499),
.B(n_1327),
.Y(n_1534)
);

AO32x2_ASAP7_75t_L g1535 ( 
.A1(n_1459),
.A2(n_1462),
.A3(n_1477),
.B1(n_1491),
.B2(n_1464),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1450),
.B(n_1412),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1434),
.B(n_1327),
.Y(n_1537)
);

AOI221xp5_ASAP7_75t_L g1538 ( 
.A1(n_1502),
.A2(n_1437),
.B1(n_1455),
.B2(n_1514),
.C(n_1479),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_SL g1539 ( 
.A(n_1469),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1483),
.B(n_1449),
.Y(n_1540)
);

OAI211xp5_ASAP7_75t_L g1541 ( 
.A1(n_1502),
.A2(n_1514),
.B(n_1448),
.C(n_1515),
.Y(n_1541)
);

OAI211xp5_ASAP7_75t_L g1542 ( 
.A1(n_1515),
.A2(n_1506),
.B(n_1505),
.C(n_1511),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1507),
.B(n_1428),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1507),
.B(n_1428),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1507),
.B(n_1438),
.Y(n_1545)
);

AOI221xp5_ASAP7_75t_L g1546 ( 
.A1(n_1437),
.A2(n_1479),
.B1(n_1513),
.B2(n_1511),
.C(n_1475),
.Y(n_1546)
);

OAI211xp5_ASAP7_75t_L g1547 ( 
.A1(n_1505),
.A2(n_1506),
.B(n_1513),
.C(n_1498),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1495),
.A2(n_1451),
.B(n_1486),
.Y(n_1548)
);

OR2x6_ASAP7_75t_L g1549 ( 
.A(n_1453),
.B(n_1441),
.Y(n_1549)
);

OA21x2_ASAP7_75t_L g1550 ( 
.A1(n_1430),
.A2(n_1456),
.B(n_1475),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1442),
.B(n_1471),
.Y(n_1551)
);

AND2x2_ASAP7_75t_SL g1552 ( 
.A(n_1440),
.B(n_1462),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1501),
.B(n_1442),
.Y(n_1553)
);

AOI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1479),
.A2(n_1473),
.B1(n_1470),
.B2(n_1503),
.C(n_1471),
.Y(n_1554)
);

CKINVDCx6p67_ASAP7_75t_R g1555 ( 
.A(n_1469),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1458),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1501),
.B(n_1510),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1497),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1471),
.B(n_1484),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1503),
.A2(n_1493),
.B1(n_1468),
.B2(n_1466),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1468),
.A2(n_1503),
.B1(n_1493),
.B2(n_1485),
.Y(n_1561)
);

AOI21xp33_ASAP7_75t_L g1562 ( 
.A1(n_1466),
.A2(n_1481),
.B(n_1470),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1466),
.B(n_1473),
.Y(n_1563)
);

AO32x1_ASAP7_75t_L g1564 ( 
.A1(n_1457),
.A2(n_1460),
.A3(n_1461),
.B1(n_1444),
.B2(n_1454),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1453),
.B(n_1456),
.Y(n_1565)
);

BUFx4f_ASAP7_75t_SL g1566 ( 
.A(n_1469),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1551),
.B(n_1461),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1551),
.B(n_1559),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1524),
.A2(n_1493),
.B1(n_1485),
.B2(n_1481),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1560),
.B(n_1489),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1533),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1543),
.B(n_1432),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1521),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1544),
.B(n_1432),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1563),
.B(n_1460),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1565),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1563),
.B(n_1431),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1521),
.B(n_1435),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1535),
.B(n_1431),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1545),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1550),
.B(n_1429),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1516),
.A2(n_1492),
.B1(n_1487),
.B2(n_1494),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1519),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1549),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1550),
.B(n_1429),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1535),
.B(n_1550),
.Y(n_1586)
);

INVx5_ASAP7_75t_L g1587 ( 
.A(n_1565),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1517),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1564),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1522),
.Y(n_1590)
);

NAND2x1p5_ASAP7_75t_SL g1591 ( 
.A(n_1532),
.B(n_1509),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1525),
.A2(n_1485),
.B1(n_1472),
.B2(n_1500),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1573),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1581),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1567),
.B(n_1528),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1578),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1584),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1569),
.A2(n_1516),
.B1(n_1561),
.B2(n_1541),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1568),
.B(n_1523),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1576),
.Y(n_1600)
);

OAI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1569),
.A2(n_1561),
.B1(n_1538),
.B2(n_1530),
.C(n_1518),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1567),
.B(n_1554),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1582),
.A2(n_1542),
.B1(n_1530),
.B2(n_1552),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1583),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1567),
.B(n_1546),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1573),
.Y(n_1606)
);

INVx5_ASAP7_75t_L g1607 ( 
.A(n_1576),
.Y(n_1607)
);

OAI222xp33_ASAP7_75t_L g1608 ( 
.A1(n_1570),
.A2(n_1536),
.B1(n_1532),
.B2(n_1558),
.C1(n_1553),
.C2(n_1540),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1583),
.B(n_1548),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1568),
.B(n_1523),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1578),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1568),
.B(n_1552),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1583),
.B(n_1586),
.Y(n_1613)
);

OR2x6_ASAP7_75t_L g1614 ( 
.A(n_1576),
.B(n_1549),
.Y(n_1614)
);

INVx4_ASAP7_75t_L g1615 ( 
.A(n_1587),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1581),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1578),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1586),
.B(n_1519),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1570),
.A2(n_1536),
.B1(n_1527),
.B2(n_1539),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1575),
.B(n_1562),
.Y(n_1620)
);

NAND3xp33_ASAP7_75t_L g1621 ( 
.A(n_1592),
.B(n_1531),
.C(n_1547),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1585),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1588),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1588),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1571),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1572),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1571),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1592),
.A2(n_1527),
.B1(n_1539),
.B2(n_1557),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1579),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1576),
.Y(n_1630)
);

OAI211xp5_ASAP7_75t_L g1631 ( 
.A1(n_1582),
.A2(n_1534),
.B(n_1500),
.C(n_1494),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1590),
.A2(n_1539),
.B1(n_1534),
.B2(n_1529),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1586),
.B(n_1519),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1618),
.B(n_1580),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1602),
.B(n_1575),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1596),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1602),
.B(n_1575),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1605),
.B(n_1577),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1596),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1611),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1605),
.B(n_1577),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1618),
.B(n_1580),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1611),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1612),
.B(n_1576),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1617),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1623),
.B(n_1577),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1607),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1617),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1620),
.B(n_1572),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1606),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1623),
.B(n_1590),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1612),
.B(n_1618),
.Y(n_1652)
);

BUFx2_ASAP7_75t_L g1653 ( 
.A(n_1614),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1620),
.B(n_1572),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1594),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1626),
.B(n_1574),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1606),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1607),
.B(n_1587),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1624),
.Y(n_1659)
);

INVxp67_ASAP7_75t_SL g1660 ( 
.A(n_1593),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1594),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1625),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1612),
.B(n_1576),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1594),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1594),
.Y(n_1665)
);

NOR2xp67_ASAP7_75t_L g1666 ( 
.A(n_1607),
.B(n_1615),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1627),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1633),
.B(n_1576),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1649),
.B(n_1609),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1638),
.B(n_1599),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1638),
.B(n_1599),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1649),
.B(n_1609),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1651),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1651),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1657),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1657),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1650),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1655),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1654),
.B(n_1609),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1641),
.B(n_1599),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1650),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1655),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1636),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1659),
.B(n_1556),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1653),
.A2(n_1598),
.B1(n_1603),
.B2(n_1621),
.Y(n_1685)
);

INVxp67_ASAP7_75t_SL g1686 ( 
.A(n_1666),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1659),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1636),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1639),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1652),
.B(n_1644),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1647),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1641),
.B(n_1610),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1654),
.B(n_1604),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1653),
.B(n_1621),
.C(n_1598),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1635),
.B(n_1556),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1639),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1652),
.B(n_1633),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1635),
.B(n_1604),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1640),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1640),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1637),
.B(n_1439),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1643),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1644),
.A2(n_1603),
.B1(n_1601),
.B2(n_1619),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1637),
.B(n_1610),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1643),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1663),
.B(n_1633),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1663),
.B(n_1668),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1668),
.B(n_1630),
.Y(n_1708)
);

AOI33xp33_ASAP7_75t_L g1709 ( 
.A1(n_1668),
.A2(n_1619),
.A3(n_1613),
.B1(n_1628),
.B2(n_1632),
.B3(n_1589),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1645),
.Y(n_1710)
);

NOR2xp67_ASAP7_75t_SL g1711 ( 
.A(n_1647),
.B(n_1631),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1690),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1705),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1687),
.B(n_1566),
.Y(n_1714)
);

OR2x6_ASAP7_75t_L g1715 ( 
.A(n_1694),
.B(n_1666),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1693),
.B(n_1660),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1693),
.B(n_1660),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1685),
.B(n_1610),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1681),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1703),
.A2(n_1601),
.B(n_1631),
.Y(n_1720)
);

NAND2xp33_ASAP7_75t_SL g1721 ( 
.A(n_1711),
.B(n_1647),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1690),
.B(n_1707),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1707),
.B(n_1647),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_L g1724 ( 
.A(n_1709),
.B(n_1628),
.C(n_1632),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1709),
.B(n_1646),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1706),
.B(n_1658),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1684),
.B(n_1566),
.Y(n_1727)
);

NAND4xp25_ASAP7_75t_L g1728 ( 
.A(n_1701),
.B(n_1658),
.C(n_1615),
.D(n_1526),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1696),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1695),
.B(n_1646),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1670),
.B(n_1645),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1671),
.B(n_1648),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1706),
.B(n_1658),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1686),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1691),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1673),
.B(n_1626),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1674),
.B(n_1595),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1708),
.B(n_1595),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1708),
.B(n_1656),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1675),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1680),
.B(n_1555),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1697),
.B(n_1658),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1696),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1692),
.B(n_1648),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1676),
.B(n_1711),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1677),
.B(n_1656),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1697),
.B(n_1634),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1704),
.B(n_1555),
.Y(n_1748)
);

OR4x1_ASAP7_75t_L g1749 ( 
.A(n_1713),
.B(n_1691),
.C(n_1702),
.D(n_1700),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1720),
.A2(n_1614),
.B1(n_1615),
.B2(n_1576),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1719),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1725),
.A2(n_1608),
.B1(n_1604),
.B2(n_1710),
.C(n_1689),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1724),
.A2(n_1607),
.B1(n_1614),
.B2(n_1669),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1734),
.B(n_1669),
.Y(n_1754)
);

AOI211x1_ASAP7_75t_L g1755 ( 
.A1(n_1745),
.A2(n_1608),
.B(n_1613),
.C(n_1634),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1722),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1734),
.B(n_1672),
.Y(n_1757)
);

OAI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1715),
.A2(n_1679),
.B(n_1672),
.Y(n_1758)
);

AOI32xp33_ASAP7_75t_L g1759 ( 
.A1(n_1721),
.A2(n_1718),
.A3(n_1722),
.B1(n_1733),
.B2(n_1726),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1721),
.A2(n_1614),
.B1(n_1615),
.B2(n_1607),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_L g1761 ( 
.A(n_1715),
.B(n_1679),
.C(n_1683),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1740),
.B(n_1698),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1730),
.B(n_1698),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1712),
.B(n_1630),
.Y(n_1764)
);

OAI322xp33_ASAP7_75t_L g1765 ( 
.A1(n_1713),
.A2(n_1717),
.A3(n_1716),
.B1(n_1712),
.B2(n_1746),
.C1(n_1739),
.C2(n_1736),
.Y(n_1765)
);

NAND3xp33_ASAP7_75t_L g1766 ( 
.A(n_1715),
.B(n_1699),
.C(n_1688),
.Y(n_1766)
);

AOI21xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1714),
.A2(n_1591),
.B(n_1600),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1735),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1715),
.A2(n_1607),
.B1(n_1615),
.B2(n_1587),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1726),
.B(n_1634),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1733),
.B(n_1642),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1729),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1742),
.B(n_1642),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1743),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1768),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1756),
.B(n_1742),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1768),
.B(n_1723),
.Y(n_1777)
);

AOI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1755),
.A2(n_1723),
.B1(n_1735),
.B2(n_1716),
.C(n_1717),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1751),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1772),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1774),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1758),
.B(n_1747),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1754),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1757),
.Y(n_1784)
);

AOI21xp33_ASAP7_75t_L g1785 ( 
.A1(n_1761),
.A2(n_1727),
.B(n_1741),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1758),
.B(n_1747),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1762),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_L g1788 ( 
.A(n_1752),
.B(n_1737),
.C(n_1728),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1766),
.B(n_1738),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1749),
.Y(n_1790)
);

AOI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1753),
.A2(n_1748),
.B1(n_1607),
.B2(n_1630),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1750),
.A2(n_1607),
.B1(n_1614),
.B2(n_1613),
.Y(n_1792)
);

OAI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1760),
.A2(n_1614),
.B1(n_1600),
.B2(n_1587),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1759),
.A2(n_1614),
.B1(n_1600),
.B2(n_1597),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1775),
.Y(n_1795)
);

O2A1O1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1790),
.A2(n_1775),
.B(n_1783),
.C(n_1784),
.Y(n_1796)
);

NAND3xp33_ASAP7_75t_L g1797 ( 
.A(n_1790),
.B(n_1769),
.C(n_1763),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1777),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1777),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1789),
.B(n_1770),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1782),
.B(n_1764),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1782),
.B(n_1771),
.Y(n_1802)
);

OAI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1788),
.A2(n_1767),
.B(n_1773),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1776),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1779),
.Y(n_1805)
);

OAI31xp33_ASAP7_75t_L g1806 ( 
.A1(n_1789),
.A2(n_1765),
.A3(n_1744),
.B(n_1732),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1798),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1798),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1799),
.B(n_1787),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1799),
.Y(n_1810)
);

NAND4xp25_ASAP7_75t_L g1811 ( 
.A(n_1796),
.B(n_1785),
.C(n_1791),
.D(n_1778),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1804),
.B(n_1789),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1804),
.B(n_1800),
.Y(n_1813)
);

NAND3xp33_ASAP7_75t_L g1814 ( 
.A(n_1806),
.B(n_1786),
.C(n_1781),
.Y(n_1814)
);

NOR3xp33_ASAP7_75t_L g1815 ( 
.A(n_1797),
.B(n_1795),
.C(n_1805),
.Y(n_1815)
);

NAND3xp33_ASAP7_75t_L g1816 ( 
.A(n_1814),
.B(n_1795),
.C(n_1803),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1811),
.A2(n_1802),
.B1(n_1786),
.B2(n_1794),
.C(n_1801),
.Y(n_1817)
);

OAI211xp5_ASAP7_75t_SL g1818 ( 
.A1(n_1815),
.A2(n_1780),
.B(n_1793),
.C(n_1792),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1812),
.B(n_1801),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1813),
.B(n_1802),
.Y(n_1820)
);

NOR3xp33_ASAP7_75t_L g1821 ( 
.A(n_1816),
.B(n_1809),
.C(n_1807),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1820),
.A2(n_1808),
.B1(n_1776),
.B2(n_1810),
.Y(n_1822)
);

AOI211xp5_ASAP7_75t_L g1823 ( 
.A1(n_1819),
.A2(n_1744),
.B(n_1732),
.C(n_1731),
.Y(n_1823)
);

OA22x2_ASAP7_75t_L g1824 ( 
.A1(n_1818),
.A2(n_1817),
.B1(n_1682),
.B2(n_1678),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1816),
.A2(n_1731),
.B1(n_1600),
.B2(n_1629),
.Y(n_1825)
);

NOR3xp33_ASAP7_75t_L g1826 ( 
.A(n_1816),
.B(n_1464),
.C(n_1463),
.Y(n_1826)
);

NOR4xp75_ASAP7_75t_L g1827 ( 
.A(n_1822),
.B(n_1600),
.C(n_1477),
.D(n_1463),
.Y(n_1827)
);

NOR2x1_ASAP7_75t_L g1828 ( 
.A(n_1825),
.B(n_1678),
.Y(n_1828)
);

XNOR2x1_ASAP7_75t_L g1829 ( 
.A(n_1824),
.B(n_1512),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1821),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1826),
.Y(n_1831)
);

NAND3x1_ASAP7_75t_L g1832 ( 
.A(n_1830),
.B(n_1823),
.C(n_1642),
.Y(n_1832)
);

OAI221xp5_ASAP7_75t_SL g1833 ( 
.A1(n_1831),
.A2(n_1829),
.B1(n_1827),
.B2(n_1828),
.C(n_1682),
.Y(n_1833)
);

OAI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1830),
.A2(n_1491),
.B1(n_1597),
.B2(n_1504),
.C(n_1664),
.Y(n_1834)
);

OAI221xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1834),
.A2(n_1504),
.B1(n_1597),
.B2(n_1665),
.C(n_1664),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1835),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1836),
.Y(n_1837)
);

AO21x2_ASAP7_75t_L g1838 ( 
.A1(n_1836),
.A2(n_1832),
.B(n_1833),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1837),
.A2(n_1665),
.B1(n_1664),
.B2(n_1661),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1838),
.A2(n_1661),
.B1(n_1655),
.B2(n_1665),
.Y(n_1840)
);

AO22x2_ASAP7_75t_L g1841 ( 
.A1(n_1840),
.A2(n_1838),
.B1(n_1661),
.B2(n_1667),
.Y(n_1841)
);

XOR2xp5_ASAP7_75t_L g1842 ( 
.A(n_1839),
.B(n_1838),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1841),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1843),
.A2(n_1842),
.B1(n_1622),
.B2(n_1616),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1844),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1597),
.B1(n_1520),
.B2(n_1662),
.Y(n_1846)
);

AOI211xp5_ASAP7_75t_L g1847 ( 
.A1(n_1846),
.A2(n_1512),
.B(n_1508),
.C(n_1537),
.Y(n_1847)
);


endmodule