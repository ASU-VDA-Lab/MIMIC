module fake_jpeg_23625_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx13_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx16_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_8),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_18),
.A2(n_11),
.B(n_12),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_25),
.B1(n_26),
.B2(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

AND2x6_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_1),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_34),
.B(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_22),
.B1(n_21),
.B2(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_22),
.B1(n_21),
.B2(n_18),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_32),
.B1(n_13),
.B2(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_23),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_50),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_12),
.B(n_14),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_21),
.C(n_13),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_38),
.C(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_38),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_60),
.B(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_61),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_43),
.C(n_37),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_53),
.C(n_51),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_16),
.B1(n_21),
.B2(n_10),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_9),
.B1(n_12),
.B2(n_10),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_63),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_50),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_9),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_56),
.C(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_70),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_59),
.B1(n_9),
.B2(n_4),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_2),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_65),
.B1(n_63),
.B2(n_16),
.Y(n_71)
);

OAI31xp33_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_69),
.A3(n_9),
.B(n_16),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_2),
.C(n_3),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.A3(n_73),
.B1(n_4),
.B2(n_5),
.C1(n_3),
.C2(n_16),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_3),
.C(n_5),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_5),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_69),
.Y(n_79)
);


endmodule