module real_aes_4839_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_1297, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_1296, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_1300, n_325, n_1298, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_1299, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_1297;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_1296;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_1300;
input n_325;
input n_1298;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_1299;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_592;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_417;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_859;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1161;
wire n_686;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1162;
wire n_762;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_414;
wire n_776;
wire n_1138;
wire n_890;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_816;
wire n_625;
wire n_953;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1060;
wire n_1154;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_974;
wire n_857;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_698;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_0), .A2(n_234), .B1(n_585), .B2(n_630), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_1), .A2(n_328), .B1(n_663), .B2(n_732), .Y(n_849) );
INVx1_ASAP7_75t_L g761 ( .A(n_2), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_3), .A2(n_254), .B1(n_672), .B2(n_680), .Y(n_1258) );
INVx1_ASAP7_75t_L g558 ( .A(n_4), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_5), .A2(n_270), .B1(n_580), .B2(n_642), .Y(n_774) );
INVx1_ASAP7_75t_L g431 ( .A(n_6), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_7), .A2(n_253), .B1(n_663), .B2(n_664), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_8), .A2(n_288), .B1(n_487), .B2(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_9), .A2(n_189), .B1(n_673), .B2(n_678), .Y(n_1257) );
INVx1_ASAP7_75t_L g969 ( .A(n_10), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_11), .A2(n_190), .B1(n_601), .B2(n_656), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_12), .A2(n_308), .B1(n_588), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_13), .A2(n_296), .B1(n_568), .B2(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g997 ( .A(n_14), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_15), .A2(n_145), .B1(n_482), .B2(n_484), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_16), .A2(n_217), .B1(n_580), .B2(n_941), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_17), .A2(n_283), .B1(n_400), .B2(n_423), .C(n_430), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g885 ( .A1(n_18), .A2(n_80), .B1(n_626), .B2(n_821), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_19), .A2(n_236), .B1(n_673), .B2(n_681), .Y(n_930) );
INVx1_ASAP7_75t_L g764 ( .A(n_20), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_21), .A2(n_300), .B1(n_583), .B2(n_626), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_22), .A2(n_24), .B1(n_583), .B2(n_585), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g1276 ( .A1(n_23), .A2(n_77), .B1(n_487), .B2(n_567), .Y(n_1276) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_25), .B(n_405), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_26), .A2(n_136), .B1(n_673), .B2(n_678), .Y(n_869) );
AOI21xp33_ASAP7_75t_L g600 ( .A1(n_27), .A2(n_601), .B(n_602), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g1026 ( .A(n_28), .Y(n_1026) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_29), .A2(n_240), .B1(n_580), .B2(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g652 ( .A(n_30), .Y(n_652) );
INVx1_ASAP7_75t_L g759 ( .A(n_31), .Y(n_759) );
AOI221x1_ASAP7_75t_L g717 ( .A1(n_32), .A2(n_94), .B1(n_718), .B2(n_719), .C(n_720), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_33), .A2(n_357), .B1(n_464), .B2(n_563), .Y(n_1278) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_34), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_35), .A2(n_41), .B1(n_585), .B2(n_630), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g1011 ( .A1(n_36), .A2(n_100), .B1(n_1012), .B2(n_1014), .Y(n_1011) );
INVx1_ASAP7_75t_L g917 ( .A(n_37), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_38), .A2(n_373), .B1(n_591), .B2(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_39), .A2(n_273), .B1(n_487), .B2(n_489), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_40), .A2(n_55), .B1(n_510), .B2(n_512), .Y(n_509) );
INVx1_ASAP7_75t_L g922 ( .A(n_42), .Y(n_922) );
AOI21xp33_ASAP7_75t_L g950 ( .A1(n_43), .A2(n_650), .B(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g855 ( .A(n_44), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_45), .A2(n_153), .B1(n_644), .B2(n_646), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_46), .A2(n_124), .B1(n_472), .B2(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_47), .A2(n_245), .B1(n_598), .B2(n_599), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_48), .A2(n_115), .B1(n_675), .B2(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g556 ( .A(n_49), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_50), .A2(n_242), .B1(n_1002), .B2(n_1004), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_51), .B(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_52), .A2(n_309), .B1(n_587), .B2(n_588), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g1254 ( .A1(n_53), .A2(n_365), .B1(n_552), .B2(n_667), .Y(n_1254) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_54), .A2(n_233), .B1(n_563), .B2(n_580), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_56), .A2(n_301), .B1(n_470), .B2(n_614), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_57), .A2(n_62), .B1(n_630), .B2(n_943), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_58), .A2(n_134), .B1(n_675), .B2(n_676), .Y(n_845) );
INVx1_ASAP7_75t_L g1024 ( .A(n_59), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_60), .A2(n_243), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_61), .A2(n_360), .B1(n_666), .B2(n_766), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_63), .A2(n_343), .B1(n_666), .B2(n_667), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_64), .A2(n_111), .B1(n_464), .B2(n_563), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_65), .B(n_799), .Y(n_1288) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_66), .A2(n_143), .B1(n_525), .B2(n_526), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_67), .A2(n_371), .B1(n_577), .B2(n_578), .Y(n_823) );
OA22x2_ASAP7_75t_L g403 ( .A1(n_68), .A2(n_162), .B1(n_404), .B2(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g442 ( .A(n_68), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_69), .A2(n_141), .B1(n_675), .B2(n_676), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_70), .A2(n_321), .B1(n_680), .B2(n_681), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_71), .A2(n_114), .B1(n_592), .B2(n_598), .Y(n_948) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_72), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_73), .A2(n_152), .B1(n_591), .B2(n_880), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_74), .A2(n_367), .B1(n_580), .B2(n_678), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_75), .A2(n_226), .B1(n_588), .B2(n_628), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_76), .B(n_552), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_78), .A2(n_313), .B1(n_588), .B2(n_703), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_79), .B(n_181), .Y(n_385) );
INVx1_ASAP7_75t_L g411 ( .A(n_79), .Y(n_411) );
OAI21xp33_ASAP7_75t_L g457 ( .A1(n_79), .A2(n_162), .B(n_458), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_81), .A2(n_339), .B1(n_577), .B2(n_578), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_82), .A2(n_354), .B1(n_675), .B2(n_676), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_83), .A2(n_251), .B1(n_535), .B2(n_537), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_84), .A2(n_260), .B1(n_577), .B2(n_578), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_85), .A2(n_225), .B1(n_577), .B2(n_646), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_86), .A2(n_237), .B1(n_614), .B2(n_799), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_87), .A2(n_182), .B1(n_400), .B2(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g971 ( .A(n_88), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_89), .A2(n_230), .B1(n_492), .B2(n_565), .Y(n_1277) );
AOI21xp33_ASAP7_75t_L g831 ( .A1(n_90), .A2(n_400), .B(n_832), .Y(n_831) );
XOR2x2_ASAP7_75t_L g958 ( .A(n_91), .B(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g996 ( .A(n_92), .Y(n_996) );
AND2x4_ASAP7_75t_L g1003 ( .A(n_92), .B(n_269), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g1293 ( .A(n_92), .Y(n_1293) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_93), .A2(n_317), .B1(n_664), .B2(n_681), .Y(n_1256) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_95), .A2(n_293), .B1(n_577), .B2(n_578), .Y(n_631) );
INVx1_ASAP7_75t_L g787 ( .A(n_96), .Y(n_787) );
INVx1_ASAP7_75t_L g973 ( .A(n_97), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_98), .A2(n_359), .B1(n_487), .B2(n_578), .Y(n_802) );
AO22x1_ASAP7_75t_L g820 ( .A1(n_99), .A2(n_316), .B1(n_626), .B2(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_101), .A2(n_180), .B1(n_799), .B2(n_882), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_102), .A2(n_122), .B1(n_568), .B2(n_724), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_103), .A2(n_150), .B1(n_591), .B2(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_104), .A2(n_322), .B1(n_547), .B2(n_829), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_105), .A2(n_118), .B1(n_470), .B2(n_472), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_106), .A2(n_227), .B1(n_591), .B2(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_107), .B(n_594), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_108), .A2(n_142), .B1(n_494), .B2(n_630), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_109), .A2(n_298), .B1(n_460), .B2(n_537), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_110), .A2(n_205), .B1(n_464), .B2(n_563), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g866 ( .A1(n_112), .A2(n_333), .B1(n_821), .B2(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g994 ( .A(n_113), .Y(n_994) );
AND2x4_ASAP7_75t_L g999 ( .A(n_113), .B(n_381), .Y(n_999) );
INVx1_ASAP7_75t_SL g1013 ( .A(n_113), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_116), .A2(n_355), .B1(n_446), .B2(n_453), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g834 ( .A(n_117), .B(n_594), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g806 ( .A1(n_119), .A2(n_121), .B1(n_492), .B2(n_565), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_120), .B(n_851), .Y(n_850) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_123), .A2(n_694), .B(n_695), .Y(n_693) );
CKINVDCx16_ASAP7_75t_R g1065 ( .A(n_125), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_126), .A2(n_149), .B1(n_992), .B2(n_1045), .Y(n_1044) );
AOI33xp33_ASAP7_75t_R g888 ( .A1(n_127), .A2(n_250), .A3(n_427), .B1(n_456), .B2(n_889), .B3(n_1300), .Y(n_888) );
INVx1_ASAP7_75t_L g506 ( .A(n_128), .Y(n_506) );
INVx1_ASAP7_75t_L g573 ( .A(n_129), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_130), .A2(n_329), .B1(n_664), .B2(n_681), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_131), .A2(n_264), .B1(n_664), .B2(n_672), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_132), .A2(n_263), .B1(n_487), .B2(n_489), .Y(n_533) );
AO22x1_ASAP7_75t_L g459 ( .A1(n_133), .A2(n_319), .B1(n_460), .B2(n_464), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_135), .A2(n_232), .B1(n_460), .B2(n_897), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g1270 ( .A1(n_137), .A2(n_1271), .B1(n_1272), .B2(n_1273), .Y(n_1270) );
CKINVDCx5p33_ASAP7_75t_R g1271 ( .A(n_137), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_138), .A2(n_165), .B1(n_628), .B2(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_139), .A2(n_259), .B1(n_672), .B2(n_673), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_140), .A2(n_197), .B1(n_616), .B2(n_656), .Y(n_1289) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_144), .A2(n_304), .B1(n_649), .B2(n_650), .C(n_651), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_146), .A2(n_345), .B1(n_530), .B2(n_531), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_147), .A2(n_151), .B1(n_464), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_148), .A2(n_287), .B1(n_512), .B2(n_619), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_154), .B(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_155), .A2(n_274), .B1(n_446), .B2(n_492), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_156), .A2(n_307), .B1(n_577), .B2(n_578), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_157), .A2(n_363), .B1(n_446), .B2(n_492), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_158), .A2(n_171), .B1(n_563), .B2(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_159), .A2(n_338), .B1(n_425), .B2(n_621), .Y(n_620) );
CKINVDCx6p67_ASAP7_75t_R g783 ( .A(n_160), .Y(n_783) );
INVx1_ASAP7_75t_L g422 ( .A(n_161), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_161), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_161), .B(n_220), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_162), .B(n_282), .Y(n_384) );
XNOR2x1_ASAP7_75t_L g841 ( .A(n_163), .B(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g937 ( .A(n_164), .Y(n_937) );
INVx1_ASAP7_75t_L g905 ( .A(n_166), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_167), .A2(n_177), .B1(n_628), .B2(n_640), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_168), .B(n_650), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_169), .A2(n_188), .B1(n_678), .B2(n_680), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_170), .A2(n_256), .B1(n_460), .B2(n_464), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_172), .A2(n_277), .B1(n_583), .B2(n_585), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_173), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g1032 ( .A1(n_174), .A2(n_334), .B1(n_1016), .B2(n_1017), .Y(n_1032) );
AOI21xp5_ASAP7_75t_L g1248 ( .A1(n_175), .A2(n_425), .B(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g967 ( .A(n_176), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_178), .A2(n_194), .B1(n_472), .B2(n_669), .Y(n_965) );
INVx1_ASAP7_75t_L g549 ( .A(n_179), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_181), .B(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_183), .A2(n_208), .B1(n_563), .B2(n_565), .Y(n_980) );
INVx1_ASAP7_75t_L g553 ( .A(n_184), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g1279 ( .A1(n_185), .A2(n_348), .B1(n_460), .B2(n_804), .Y(n_1279) );
AOI22xp5_ASAP7_75t_L g1015 ( .A1(n_186), .A2(n_289), .B1(n_1016), .B2(n_1017), .Y(n_1015) );
AO22x2_ASAP7_75t_L g1242 ( .A1(n_186), .A2(n_1243), .B1(n_1260), .B2(n_1261), .Y(n_1242) );
INVxp67_ASAP7_75t_SL g1260 ( .A(n_186), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g1267 ( .A1(n_186), .A2(n_1268), .B1(n_1270), .B2(n_1290), .Y(n_1267) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_187), .A2(n_326), .B1(n_515), .B2(n_517), .Y(n_514) );
INVx1_ASAP7_75t_L g910 ( .A(n_191), .Y(n_910) );
INVx1_ASAP7_75t_L g1067 ( .A(n_192), .Y(n_1067) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_193), .A2(n_306), .B1(n_460), .B2(n_804), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g736 ( .A(n_195), .Y(n_736) );
INVx1_ASAP7_75t_L g952 ( .A(n_196), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_198), .B(n_482), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_199), .A2(n_366), .B1(n_673), .B2(n_678), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_200), .A2(n_340), .B1(n_591), .B2(n_614), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_201), .A2(n_374), .B1(n_591), .B2(n_829), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_202), .A2(n_302), .B1(n_992), .B2(n_1039), .Y(n_1038) );
INVx1_ASAP7_75t_L g754 ( .A(n_203), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_204), .A2(n_238), .B1(n_640), .B2(n_672), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_206), .A2(n_368), .B1(n_650), .B2(n_669), .Y(n_668) );
BUFx2_ASAP7_75t_L g1251 ( .A(n_207), .Y(n_1251) );
INVx1_ASAP7_75t_L g916 ( .A(n_209), .Y(n_916) );
INVx1_ASAP7_75t_L g861 ( .A(n_210), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g1031 ( .A1(n_211), .A2(n_350), .B1(n_1012), .B2(n_1014), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_212), .A2(n_318), .B1(n_492), .B2(n_494), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_213), .A2(n_281), .B1(n_1004), .B2(n_1036), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_214), .A2(n_278), .B1(n_672), .B2(n_680), .Y(n_727) );
XOR2x2_ASAP7_75t_L g875 ( .A(n_215), .B(n_876), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g978 ( .A1(n_216), .A2(n_299), .B1(n_489), .B2(n_979), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_218), .A2(n_276), .B1(n_649), .B2(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_219), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g409 ( .A(n_220), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_221), .A2(n_358), .B1(n_675), .B2(n_676), .Y(n_933) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_222), .A2(n_336), .B1(n_591), .B2(n_654), .Y(n_699) );
INVx1_ASAP7_75t_L g397 ( .A(n_223), .Y(n_397) );
OAI222xp33_ASAP7_75t_L g467 ( .A1(n_223), .A2(n_468), .B1(n_486), .B2(n_491), .C1(n_1296), .C2(n_1297), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_223), .B(n_491), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g738 ( .A(n_224), .Y(n_738) );
INVx1_ASAP7_75t_L g635 ( .A(n_228), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_229), .A2(n_356), .B1(n_664), .B2(n_672), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_231), .A2(n_241), .B1(n_1036), .B2(n_1037), .Y(n_1035) );
INVx1_ASAP7_75t_L g1287 ( .A(n_235), .Y(n_1287) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_239), .A2(n_291), .B1(n_587), .B2(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_244), .A2(n_362), .B1(n_650), .B2(n_667), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_246), .A2(n_266), .B1(n_992), .B2(n_1039), .Y(n_1050) );
OAI21x1_ASAP7_75t_L g815 ( .A1(n_247), .A2(n_816), .B(n_835), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_247), .B(n_819), .Y(n_838) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_248), .A2(n_341), .B1(n_649), .B2(n_851), .C(n_860), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_249), .A2(n_258), .B1(n_512), .B2(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_252), .A2(n_320), .B1(n_492), .B2(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g794 ( .A(n_255), .Y(n_794) );
INVx1_ASAP7_75t_L g603 ( .A(n_257), .Y(n_603) );
INVx1_ASAP7_75t_L g544 ( .A(n_261), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_262), .A2(n_297), .B1(n_588), .B2(n_628), .Y(n_770) );
INVx1_ASAP7_75t_L g962 ( .A(n_265), .Y(n_962) );
INVx1_ASAP7_75t_L g689 ( .A(n_266), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_266), .B(n_706), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_267), .A2(n_290), .B1(n_1002), .B2(n_1037), .Y(n_1049) );
AOI21xp5_ASAP7_75t_L g1283 ( .A1(n_268), .A2(n_1284), .B(n_1286), .Y(n_1283) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_269), .Y(n_386) );
AND2x4_ASAP7_75t_L g995 ( .A(n_269), .B(n_996), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_271), .A2(n_280), .B1(n_680), .B2(n_681), .Y(n_679) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_272), .Y(n_733) );
XNOR2x1_ASAP7_75t_L g856 ( .A(n_275), .B(n_857), .Y(n_856) );
AOI211x1_ASAP7_75t_L g901 ( .A1(n_279), .A2(n_902), .B(n_904), .C(n_912), .Y(n_901) );
INVx1_ASAP7_75t_L g420 ( .A(n_282), .Y(n_420) );
INVxp67_ASAP7_75t_L g480 ( .A(n_282), .Y(n_480) );
INVx1_ASAP7_75t_L g833 ( .A(n_284), .Y(n_833) );
INVx1_ASAP7_75t_L g788 ( .A(n_285), .Y(n_788) );
AOI21xp33_ASAP7_75t_SL g1245 ( .A1(n_286), .A2(n_598), .B(n_1246), .Y(n_1245) );
INVxp67_ASAP7_75t_R g1069 ( .A(n_292), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_294), .A2(n_332), .B1(n_487), .B2(n_489), .Y(n_486) );
INVx2_ASAP7_75t_L g381 ( .A(n_295), .Y(n_381) );
INVx1_ASAP7_75t_SL g716 ( .A(n_302), .Y(n_716) );
NOR3xp33_ASAP7_75t_L g744 ( .A(n_302), .B(n_745), .C(n_746), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_303), .A2(n_347), .B1(n_601), .B2(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g756 ( .A(n_305), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_310), .A2(n_311), .B1(n_663), .B2(n_667), .Y(n_926) );
AOI21xp33_ASAP7_75t_L g853 ( .A1(n_312), .A2(n_649), .B(n_854), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_314), .A2(n_335), .B1(n_592), .B2(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_315), .A2(n_330), .B1(n_649), .B2(n_666), .Y(n_925) );
INVx1_ASAP7_75t_L g1247 ( .A(n_323), .Y(n_1247) );
INVx1_ASAP7_75t_L g696 ( .A(n_324), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_325), .B(n_482), .Y(n_883) );
INVx1_ASAP7_75t_L g792 ( .A(n_327), .Y(n_792) );
XOR2xp5_ASAP7_75t_L g658 ( .A(n_331), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g1022 ( .A(n_337), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_342), .A2(n_346), .B1(n_552), .B2(n_592), .Y(n_827) );
INVx1_ASAP7_75t_L g632 ( .A(n_344), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_349), .A2(n_372), .B1(n_799), .B2(n_851), .Y(n_927) );
AO22x2_ASAP7_75t_L g748 ( .A1(n_350), .A2(n_749), .B1(n_750), .B2(n_751), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_350), .Y(n_749) );
AND2x2_ASAP7_75t_L g720 ( .A(n_351), .B(n_526), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_352), .A2(n_369), .B1(n_804), .B2(n_976), .Y(n_975) );
BUFx2_ASAP7_75t_L g1253 ( .A(n_353), .Y(n_1253) );
INVx1_ASAP7_75t_L g914 ( .A(n_361), .Y(n_914) );
INVx1_ASAP7_75t_L g1000 ( .A(n_364), .Y(n_1000) );
INVx1_ASAP7_75t_L g796 ( .A(n_370), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_387), .B(n_985), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx4_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
NAND3xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_382), .C(n_386), .Y(n_378) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_379), .B(n_1265), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_379), .B(n_1266), .Y(n_1269) );
AOI21xp5_ASAP7_75t_L g1294 ( .A1(n_379), .A2(n_386), .B(n_1013), .Y(n_1294) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AO21x1_ASAP7_75t_L g1291 ( .A1(n_380), .A2(n_1292), .B(n_1294), .Y(n_1291) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g993 ( .A(n_381), .B(n_994), .Y(n_993) );
AND3x4_ASAP7_75t_L g1012 ( .A(n_381), .B(n_995), .C(n_1013), .Y(n_1012) );
NOR2xp33_ASAP7_75t_L g1265 ( .A(n_382), .B(n_1266), .Y(n_1265) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AO21x2_ASAP7_75t_L g434 ( .A1(n_383), .A2(n_435), .B(n_437), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g1266 ( .A(n_386), .Y(n_1266) );
XNOR2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_810), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_683), .B2(n_684), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_605), .B1(n_606), .B2(n_682), .Y(n_390) );
INVx1_ASAP7_75t_L g682 ( .A(n_391), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_538), .B2(n_604), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_504), .B2(n_505), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_396), .B(n_497), .Y(n_395) );
AOI21x1_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_467), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_443), .Y(n_398) );
BUFx2_ASAP7_75t_L g498 ( .A(n_399), .Y(n_498) );
INVx4_ASAP7_75t_L g557 ( .A(n_400), .Y(n_557) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g516 ( .A(n_401), .Y(n_516) );
BUFx3_ASAP7_75t_L g598 ( .A(n_401), .Y(n_598) );
BUFx3_ASAP7_75t_L g619 ( .A(n_401), .Y(n_619) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_412), .Y(n_401) );
AND2x4_ASAP7_75t_L g483 ( .A(n_402), .B(n_428), .Y(n_483) );
AND2x4_ASAP7_75t_L g649 ( .A(n_402), .B(n_412), .Y(n_649) );
AND2x2_ASAP7_75t_L g851 ( .A(n_402), .B(n_428), .Y(n_851) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_406), .Y(n_402) );
AND2x2_ASAP7_75t_L g427 ( .A(n_403), .B(n_407), .Y(n_427) );
INVx1_ASAP7_75t_L g449 ( .A(n_403), .Y(n_449) );
AND2x2_ASAP7_75t_L g478 ( .A(n_403), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_404), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2xp33_ASAP7_75t_L g408 ( .A(n_405), .B(n_409), .Y(n_408) );
INVx3_ASAP7_75t_L g415 ( .A(n_405), .Y(n_415) );
NAND2xp33_ASAP7_75t_L g421 ( .A(n_405), .B(n_422), .Y(n_421) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_405), .Y(n_436) );
INVx1_ASAP7_75t_L g458 ( .A(n_405), .Y(n_458) );
AND2x4_ASAP7_75t_L g448 ( .A(n_406), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_409), .B(n_442), .Y(n_441) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_411), .A2(n_458), .B(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g471 ( .A(n_412), .B(n_427), .Y(n_471) );
AND2x4_ASAP7_75t_L g488 ( .A(n_412), .B(n_448), .Y(n_488) );
AND2x4_ASAP7_75t_L g663 ( .A(n_412), .B(n_427), .Y(n_663) );
AND2x4_ASAP7_75t_L g675 ( .A(n_412), .B(n_448), .Y(n_675) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_417), .Y(n_412) );
INVx2_ASAP7_75t_L g429 ( .A(n_413), .Y(n_429) );
OR2x2_ASAP7_75t_L g451 ( .A(n_413), .B(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g462 ( .A(n_413), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g475 ( .A(n_413), .B(n_476), .Y(n_475) );
AND2x4_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_415), .B(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g439 ( .A(n_415), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_416), .B(n_438), .C(n_440), .Y(n_437) );
AND2x4_ASAP7_75t_L g428 ( .A(n_417), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g452 ( .A(n_418), .Y(n_452) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g545 ( .A(n_423), .Y(n_545) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI21xp33_ASAP7_75t_L g763 ( .A1(n_424), .A2(n_764), .B(n_765), .Y(n_763) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g523 ( .A(n_426), .Y(n_523) );
INVx3_ASAP7_75t_L g595 ( .A(n_426), .Y(n_595) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
AND2x2_ASAP7_75t_L g461 ( .A(n_427), .B(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g465 ( .A(n_427), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g584 ( .A(n_427), .B(n_462), .Y(n_584) );
AND2x2_ASAP7_75t_L g650 ( .A(n_427), .B(n_428), .Y(n_650) );
AND2x4_ASAP7_75t_L g673 ( .A(n_427), .B(n_450), .Y(n_673) );
AND2x4_ASAP7_75t_L g678 ( .A(n_427), .B(n_462), .Y(n_678) );
AND2x4_ASAP7_75t_L g485 ( .A(n_428), .B(n_456), .Y(n_485) );
AND2x2_ASAP7_75t_L g490 ( .A(n_428), .B(n_448), .Y(n_490) );
AND2x4_ASAP7_75t_L g667 ( .A(n_428), .B(n_456), .Y(n_667) );
AND2x4_ASAP7_75t_L g676 ( .A(n_428), .B(n_448), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx4_ASAP7_75t_L g547 ( .A(n_432), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_432), .B(n_603), .Y(n_602) );
INVx4_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx3_ASAP7_75t_L g527 ( .A(n_433), .Y(n_527) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_434), .Y(n_623) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_436), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_439), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g456 ( .A(n_440), .B(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_459), .Y(n_443) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g502 ( .A(n_445), .B(n_486), .Y(n_502) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_447), .Y(n_565) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_447), .Y(n_588) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_447), .Y(n_640) );
AND2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_450), .Y(n_447) );
AND2x4_ASAP7_75t_L g493 ( .A(n_448), .B(n_462), .Y(n_493) );
AND2x4_ASAP7_75t_L g664 ( .A(n_448), .B(n_466), .Y(n_664) );
AND2x4_ASAP7_75t_L g672 ( .A(n_448), .B(n_462), .Y(n_672) );
AND2x4_ASAP7_75t_L g455 ( .A(n_450), .B(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g681 ( .A(n_450), .B(n_456), .Y(n_681) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g466 ( .A(n_451), .Y(n_466) );
INVx1_ASAP7_75t_L g463 ( .A(n_452), .Y(n_463) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g531 ( .A(n_454), .Y(n_531) );
INVx3_ASAP7_75t_L g642 ( .A(n_454), .Y(n_642) );
INVx2_ASAP7_75t_L g703 ( .A(n_454), .Y(n_703) );
INVx5_ASAP7_75t_L g821 ( .A(n_454), .Y(n_821) );
INVx2_ASAP7_75t_L g941 ( .A(n_454), .Y(n_941) );
INVx6_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx12f_ASAP7_75t_L g563 ( .A(n_455), .Y(n_563) );
AND2x4_ASAP7_75t_L g496 ( .A(n_456), .B(n_462), .Y(n_496) );
AND2x4_ASAP7_75t_L g680 ( .A(n_456), .B(n_462), .Y(n_680) );
INVx1_ASAP7_75t_L g503 ( .A(n_459), .Y(n_503) );
BUFx8_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_461), .Y(n_536) );
HB1xp67_ASAP7_75t_L g889 ( .A(n_462), .Y(n_889) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx3_ASAP7_75t_L g530 ( .A(n_465), .Y(n_530) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_465), .Y(n_580) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_465), .Y(n_626) );
INVx1_ASAP7_75t_L g501 ( .A(n_468), .Y(n_501) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_481), .Y(n_468) );
INVx2_ASAP7_75t_L g915 ( .A(n_470), .Y(n_915) );
BUFx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g519 ( .A(n_471), .Y(n_519) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_471), .Y(n_591) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g525 ( .A(n_473), .Y(n_525) );
INVx4_ASAP7_75t_L g599 ( .A(n_473), .Y(n_599) );
INVx2_ASAP7_75t_L g654 ( .A(n_473), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g1286 ( .A1(n_473), .A2(n_1287), .B(n_1288), .Y(n_1286) );
INVx5_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g614 ( .A(n_474), .Y(n_614) );
BUFx4f_ASAP7_75t_L g829 ( .A(n_474), .Y(n_829) );
BUFx2_ASAP7_75t_L g880 ( .A(n_474), .Y(n_880) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_478), .Y(n_474) );
AND2x2_ASAP7_75t_L g666 ( .A(n_475), .B(n_478), .Y(n_666) );
AND2x4_ASAP7_75t_L g732 ( .A(n_475), .B(n_478), .Y(n_732) );
INVx2_ASAP7_75t_L g968 ( .A(n_482), .Y(n_968) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g511 ( .A(n_483), .Y(n_511) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_483), .Y(n_552) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_483), .Y(n_601) );
INVx2_ASAP7_75t_L g617 ( .A(n_483), .Y(n_617) );
BUFx8_ASAP7_75t_SL g718 ( .A(n_483), .Y(n_718) );
INVx4_ASAP7_75t_L g554 ( .A(n_484), .Y(n_554) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx3_ASAP7_75t_L g513 ( .A(n_485), .Y(n_513) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_485), .Y(n_592) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx12f_ASAP7_75t_L g577 ( .A(n_488), .Y(n_577) );
INVx3_ASAP7_75t_L g645 ( .A(n_488), .Y(n_645) );
BUFx5_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g569 ( .A(n_490), .Y(n_569) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_490), .Y(n_578) );
BUFx3_ASAP7_75t_L g646 ( .A(n_490), .Y(n_646) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_493), .Y(n_587) );
BUFx12f_ASAP7_75t_L g628 ( .A(n_493), .Y(n_628) );
INVx4_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g537 ( .A(n_495), .Y(n_537) );
INVx4_ASAP7_75t_L g585 ( .A(n_495), .Y(n_585) );
INVx1_ASAP7_75t_L g705 ( .A(n_495), .Y(n_705) );
INVx4_ASAP7_75t_L g804 ( .A(n_495), .Y(n_804) );
INVx1_ASAP7_75t_L g897 ( .A(n_495), .Y(n_897) );
INVx2_ASAP7_75t_SL g943 ( .A(n_495), .Y(n_943) );
INVx8_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND4xp75_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .C(n_502), .D(n_503), .Y(n_497) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
XNOR2x1_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_506), .A2(n_998), .B1(n_1021), .B2(n_1022), .Y(n_1020) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_528), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g508 ( .A(n_509), .B(n_514), .C(n_520), .D(n_524), .Y(n_508) );
INVx2_ASAP7_75t_L g793 ( .A(n_510), .Y(n_793) );
INVx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
OAI21xp5_ASAP7_75t_SL g909 ( .A1(n_511), .A2(n_910), .B(n_911), .Y(n_909) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g656 ( .A(n_513), .Y(n_656) );
INVx2_ASAP7_75t_L g698 ( .A(n_513), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_513), .A2(n_792), .B1(n_793), .B2(n_794), .Y(n_791) );
INVx2_ASAP7_75t_L g972 ( .A(n_515), .Y(n_972) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g694 ( .A(n_516), .Y(n_694) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g560 ( .A(n_518), .Y(n_560) );
INVx2_ASAP7_75t_L g1282 ( .A(n_518), .Y(n_1282) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g790 ( .A(n_519), .Y(n_790) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g964 ( .A(n_522), .Y(n_964) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g882 ( .A(n_523), .Y(n_882) );
INVx4_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g1246 ( .A(n_527), .B(n_1247), .Y(n_1246) );
NAND4xp25_ASAP7_75t_L g528 ( .A(n_529), .B(n_532), .C(n_533), .D(n_534), .Y(n_528) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g604 ( .A(n_538), .Y(n_604) );
XOR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_571), .Y(n_538) );
XNOR2xp5_ASAP7_75t_SL g539 ( .A(n_540), .B(n_541), .Y(n_539) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_561), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_548), .C(n_555), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .B(n_546), .Y(n_543) );
OAI22xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B1(n_553), .B2(n_554), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g760 ( .A(n_552), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_554), .A2(n_967), .B1(n_968), .B2(n_969), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_557), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_786) );
INVxp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND4x1_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .C(n_566), .D(n_570), .Y(n_561) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
XNOR2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NOR4xp75_ASAP7_75t_L g574 ( .A(n_575), .B(n_581), .C(n_589), .D(n_596), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_586), .Y(n_581) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx4f_ASAP7_75t_L g630 ( .A(n_584), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_593), .Y(n_589) );
INVx3_ASAP7_75t_L g757 ( .A(n_591), .Y(n_757) );
INVx3_ASAP7_75t_L g762 ( .A(n_592), .Y(n_762) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g719 ( .A(n_595), .Y(n_719) );
INVx2_ASAP7_75t_L g863 ( .A(n_595), .Y(n_863) );
INVx2_ASAP7_75t_L g907 ( .A(n_595), .Y(n_907) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_597), .B(n_600), .Y(n_596) );
INVx2_ASAP7_75t_L g903 ( .A(n_598), .Y(n_903) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
XNOR2x1_ASAP7_75t_L g607 ( .A(n_608), .B(n_633), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
XOR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_632), .Y(n_610) );
NOR2x1_ASAP7_75t_L g611 ( .A(n_612), .B(n_624), .Y(n_611) );
NAND4xp25_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .C(n_618), .D(n_620), .Y(n_612) );
INVx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g755 ( .A(n_619), .Y(n_755) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_622), .B(n_652), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_622), .B(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_622), .B(n_833), .Y(n_832) );
NOR2xp67_ASAP7_75t_SL g860 ( .A(n_622), .B(n_861), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_622), .B(n_952), .Y(n_951) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g669 ( .A(n_623), .Y(n_669) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_623), .Y(n_767) );
INVx2_ASAP7_75t_L g799 ( .A(n_623), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_623), .B(n_855), .Y(n_854) );
NAND4xp25_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .C(n_629), .D(n_631), .Y(n_624) );
BUFx12f_ASAP7_75t_L g976 ( .A(n_628), .Y(n_976) );
XNOR2x1_ASAP7_75t_L g633 ( .A(n_634), .B(n_657), .Y(n_633) );
XNOR2x1_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_637), .B(n_647), .Y(n_636) );
NAND4xp25_ASAP7_75t_SL g637 ( .A(n_638), .B(n_639), .C(n_641), .D(n_643), .Y(n_637) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g724 ( .A(n_645), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_653), .C(n_655), .Y(n_647) );
INVx2_ASAP7_75t_L g737 ( .A(n_649), .Y(n_737) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_670), .Y(n_659) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .C(n_665), .D(n_668), .Y(n_660) );
INVx2_ASAP7_75t_L g739 ( .A(n_663), .Y(n_739) );
INVx2_ASAP7_75t_L g734 ( .A(n_667), .Y(n_734) );
NAND4xp25_ASAP7_75t_L g670 ( .A(n_671), .B(n_674), .C(n_677), .D(n_679), .Y(n_670) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_680), .Y(n_867) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AO22x2_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B1(n_778), .B2(n_809), .Y(n_684) );
INVx2_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
AO22x2_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_747), .B1(n_775), .B2(n_776), .Y(n_686) );
INVx1_ASAP7_75t_L g775 ( .A(n_687), .Y(n_775) );
XNOR2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_712), .Y(n_687) );
OAI21x1_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B(n_709), .Y(n_688) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_700), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_691), .B(n_710), .C(n_711), .Y(n_709) );
AND4x1_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .C(n_697), .D(n_699), .Y(n_691) );
INVx1_ASAP7_75t_L g913 ( .A(n_698), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_706), .Y(n_700) );
INVxp67_ASAP7_75t_SL g711 ( .A(n_701), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g781 ( .A(n_712), .Y(n_781) );
NAND2x1_ASAP7_75t_L g712 ( .A(n_713), .B(n_740), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_721), .C(n_726), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_717), .B2(n_1298), .Y(n_714) );
INVx1_ASAP7_75t_L g745 ( .A(n_715), .Y(n_745) );
NOR2xp67_ASAP7_75t_L g721 ( .A(n_716), .B(n_722), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_716), .A2(n_727), .B1(n_728), .B2(n_1299), .Y(n_726) );
INVx1_ASAP7_75t_L g742 ( .A(n_717), .Y(n_742) );
INVx1_ASAP7_75t_L g797 ( .A(n_719), .Y(n_797) );
INVx1_ASAP7_75t_L g1285 ( .A(n_719), .Y(n_1285) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_722), .B(n_741), .C(n_744), .Y(n_740) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
BUFx4f_ASAP7_75t_L g979 ( .A(n_724), .Y(n_979) );
INVx1_ASAP7_75t_L g746 ( .A(n_727), .Y(n_746) );
INVx1_ASAP7_75t_L g743 ( .A(n_728), .Y(n_743) );
NOR2x1_ASAP7_75t_L g728 ( .A(n_729), .B(n_735), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B1(n_733), .B2(n_734), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g1249 ( .A1(n_731), .A2(n_739), .B1(n_1250), .B2(n_1252), .Y(n_1249) );
INVx4_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g777 ( .A(n_748), .Y(n_777) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_768), .Y(n_751) );
NOR3xp33_ASAP7_75t_SL g752 ( .A(n_753), .B(n_758), .C(n_763), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_761), .B2(n_762), .Y(n_758) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_772), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_779), .Y(n_809) );
OAI22xp5_ASAP7_75t_SL g779 ( .A1(n_780), .A2(n_781), .B1(n_782), .B2(n_808), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVxp67_ASAP7_75t_SL g808 ( .A(n_782), .Y(n_808) );
XNOR2x1_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_783), .A2(n_991), .B1(n_998), .B2(n_1065), .Y(n_1064) );
NAND2x1_ASAP7_75t_L g784 ( .A(n_785), .B(n_800), .Y(n_784) );
NOR3xp33_ASAP7_75t_SL g785 ( .A(n_786), .B(n_791), .C(n_795), .Y(n_785) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OAI21xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_797), .B(n_798), .Y(n_795) );
NOR2x1_ASAP7_75t_L g800 ( .A(n_801), .B(n_805), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_890), .B1(n_983), .B2(n_984), .Y(n_810) );
INVx1_ASAP7_75t_L g983 ( .A(n_811), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_813), .B1(n_872), .B2(n_873), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
OA22x2_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_839), .B1(n_840), .B2(n_871), .Y(n_813) );
INVx2_ASAP7_75t_L g871 ( .A(n_814), .Y(n_871) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g816 ( .A(n_817), .B(n_825), .Y(n_816) );
NOR3xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_820), .C(n_822), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NOR3xp33_ASAP7_75t_L g837 ( .A(n_820), .B(n_830), .C(n_838), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_822), .B(n_826), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_830), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_834), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
XNOR2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_856), .Y(n_840) );
OR2x2_ASAP7_75t_L g842 ( .A(n_843), .B(n_848), .Y(n_842) );
NAND4xp25_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .C(n_846), .D(n_847), .Y(n_843) );
NAND4xp25_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .C(n_852), .D(n_853), .Y(n_848) );
NOR2x1_ASAP7_75t_L g857 ( .A(n_858), .B(n_865), .Y(n_857) );
NAND3xp33_ASAP7_75t_L g858 ( .A(n_859), .B(n_862), .C(n_864), .Y(n_858) );
NAND4xp25_ASAP7_75t_L g865 ( .A(n_866), .B(n_868), .C(n_869), .D(n_870), .Y(n_865) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NOR2x1_ASAP7_75t_L g876 ( .A(n_877), .B(n_884), .Y(n_876) );
NAND4xp25_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .C(n_881), .D(n_883), .Y(n_877) );
NAND4xp25_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .C(n_887), .D(n_888), .Y(n_884) );
INVx1_ASAP7_75t_L g984 ( .A(n_890), .Y(n_984) );
AOI22xp5_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_956), .B1(n_981), .B2(n_982), .Y(n_890) );
INVx2_ASAP7_75t_SL g982 ( .A(n_891), .Y(n_982) );
OA22x2_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_918), .B1(n_919), .B2(n_955), .Y(n_891) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g955 ( .A(n_893), .Y(n_955) );
XNOR2x1_ASAP7_75t_L g893 ( .A(n_894), .B(n_917), .Y(n_893) );
NAND2x1_ASAP7_75t_L g894 ( .A(n_895), .B(n_901), .Y(n_894) );
AND4x1_ASAP7_75t_L g895 ( .A(n_896), .B(n_898), .C(n_899), .D(n_900), .Y(n_895) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
OAI21xp5_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .B(n_908), .Y(n_904) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_914), .B1(n_915), .B2(n_916), .Y(n_912) );
OAI22xp33_ASAP7_75t_L g970 ( .A1(n_915), .A2(n_971), .B1(n_972), .B2(n_973), .Y(n_970) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
AOI22x1_ASAP7_75t_L g919 ( .A1(n_920), .A2(n_934), .B1(n_953), .B2(n_954), .Y(n_919) );
INVx2_ASAP7_75t_L g954 ( .A(n_920), .Y(n_954) );
XNOR2x1_ASAP7_75t_L g957 ( .A(n_920), .B(n_958), .Y(n_957) );
INVx3_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
XNOR2x1_ASAP7_75t_L g921 ( .A(n_922), .B(n_923), .Y(n_921) );
OR2x2_ASAP7_75t_L g923 ( .A(n_924), .B(n_929), .Y(n_923) );
NAND4xp25_ASAP7_75t_L g924 ( .A(n_925), .B(n_926), .C(n_927), .D(n_928), .Y(n_924) );
NAND4xp25_ASAP7_75t_L g929 ( .A(n_930), .B(n_931), .C(n_932), .D(n_933), .Y(n_929) );
INVxp67_ASAP7_75t_SL g934 ( .A(n_935), .Y(n_934) );
BUFx2_ASAP7_75t_L g953 ( .A(n_935), .Y(n_953) );
XNOR2x1_ASAP7_75t_L g935 ( .A(n_936), .B(n_938), .Y(n_935) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_937), .Y(n_936) );
NOR2x1_ASAP7_75t_L g938 ( .A(n_939), .B(n_946), .Y(n_938) );
NAND4xp25_ASAP7_75t_L g939 ( .A(n_940), .B(n_942), .C(n_944), .D(n_945), .Y(n_939) );
NAND4xp25_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .C(n_949), .D(n_950), .Y(n_946) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g981 ( .A(n_957), .Y(n_981) );
NAND2x1_ASAP7_75t_L g959 ( .A(n_960), .B(n_974), .Y(n_959) );
NOR3xp33_ASAP7_75t_L g960 ( .A(n_961), .B(n_966), .C(n_970), .Y(n_960) );
OAI21xp5_ASAP7_75t_L g961 ( .A1(n_962), .A2(n_963), .B(n_965), .Y(n_961) );
INVx2_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
AND4x1_ASAP7_75t_L g974 ( .A(n_975), .B(n_977), .C(n_978), .D(n_980), .Y(n_974) );
OAI221xp5_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_1235), .B1(n_1237), .B2(n_1262), .C(n_1267), .Y(n_985) );
AOI211xp5_ASAP7_75t_L g986 ( .A1(n_987), .A2(n_1005), .B(n_1139), .C(n_1202), .Y(n_986) );
HB1xp67_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
CKINVDCx16_ASAP7_75t_R g1153 ( .A(n_988), .Y(n_1153) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_989), .B(n_1179), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_989), .B(n_1042), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_989), .B(n_1073), .Y(n_1220) );
BUFx3_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx2_ASAP7_75t_L g1171 ( .A(n_990), .Y(n_1171) );
OAI221xp5_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_997), .B1(n_998), .B2(n_1000), .C(n_1001), .Y(n_990) );
INVx3_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
AND2x4_ASAP7_75t_L g992 ( .A(n_993), .B(n_995), .Y(n_992) );
AND2x4_ASAP7_75t_L g1002 ( .A(n_993), .B(n_1003), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_993), .B(n_1003), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_993), .B(n_1003), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_995), .B(n_999), .Y(n_998) );
AND2x4_ASAP7_75t_L g1014 ( .A(n_995), .B(n_999), .Y(n_1014) );
AND2x4_ASAP7_75t_L g1039 ( .A(n_995), .B(n_999), .Y(n_1039) );
AND2x4_ASAP7_75t_L g1004 ( .A(n_999), .B(n_1003), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_999), .B(n_1003), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_999), .B(n_1003), .Y(n_1037) );
INVx3_ASAP7_75t_L g1068 ( .A(n_1002), .Y(n_1068) );
BUFx2_ASAP7_75t_L g1236 ( .A(n_1002), .Y(n_1236) );
INVx2_ASAP7_75t_L g1070 ( .A(n_1004), .Y(n_1070) );
NAND4xp25_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1094), .C(n_1117), .D(n_1135), .Y(n_1005) );
AOI211xp5_ASAP7_75t_SL g1006 ( .A1(n_1007), .A2(n_1040), .B(n_1051), .C(n_1076), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1018), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_1008), .B(n_1061), .Y(n_1084) );
NOR2xp33_ASAP7_75t_L g1197 ( .A(n_1008), .B(n_1033), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1008), .B(n_1033), .Y(n_1212) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1010), .B(n_1057), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1010), .B(n_1075), .Y(n_1074) );
CKINVDCx6p67_ASAP7_75t_R g1081 ( .A(n_1010), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1010), .B(n_1161), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1170 ( .A(n_1010), .B(n_1030), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1010), .B(n_1030), .Y(n_1190) );
NOR2xp33_ASAP7_75t_L g1206 ( .A(n_1010), .B(n_1029), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1015), .Y(n_1010) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1012), .Y(n_1021) );
INVx2_ASAP7_75t_SL g1046 ( .A(n_1014), .Y(n_1046) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1016), .Y(n_1027) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1017), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1028), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_1019), .B(n_1056), .Y(n_1055) );
CKINVDCx6p67_ASAP7_75t_R g1061 ( .A(n_1019), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1019), .B(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1019), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1019), .B(n_1134), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1019), .B(n_1092), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_1019), .A2(n_1110), .B1(n_1174), .B2(n_1176), .Y(n_1173) );
NOR2xp33_ASAP7_75t_L g1198 ( .A(n_1019), .B(n_1063), .Y(n_1198) );
NAND4xp25_ASAP7_75t_L g1201 ( .A(n_1019), .B(n_1029), .C(n_1153), .D(n_1157), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1019), .B(n_1072), .Y(n_1230) );
OR2x6_ASAP7_75t_SL g1019 ( .A(n_1020), .B(n_1023), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_1024), .A2(n_1025), .B1(n_1026), .B2(n_1027), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1028), .B(n_1084), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1028), .B(n_1061), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1028), .B(n_1093), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1033), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1029), .B(n_1034), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1029), .B(n_1084), .Y(n_1109) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_1030), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1030), .B(n_1033), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1030), .B(n_1034), .Y(n_1092) );
OAI32xp33_ASAP7_75t_L g1125 ( .A1(n_1030), .A2(n_1103), .A3(n_1126), .B1(n_1130), .B2(n_1133), .Y(n_1125) );
AND2x4_ASAP7_75t_SL g1030 ( .A(n_1031), .B(n_1032), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1033), .B(n_1081), .Y(n_1134) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1033), .Y(n_1144) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1038), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1040), .B(n_1124), .Y(n_1123) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
O2A1O1Ixp33_ASAP7_75t_L g1166 ( .A1(n_1041), .A2(n_1167), .B(n_1168), .C(n_1171), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1047), .Y(n_1041) );
INVx3_ASAP7_75t_L g1073 ( .A(n_1042), .Y(n_1073) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1042), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1042), .B(n_1048), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1042), .B(n_1062), .Y(n_1116) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1042), .B(n_1128), .Y(n_1127) );
OR2x2_ASAP7_75t_L g1132 ( .A(n_1042), .B(n_1047), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1042), .B(n_1158), .Y(n_1157) );
AND2x4_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1044), .Y(n_1042) );
INVx2_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVx3_ASAP7_75t_L g1053 ( .A(n_1047), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1047), .B(n_1063), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1047), .B(n_1073), .Y(n_1137) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1048), .B(n_1063), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1048), .B(n_1072), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1112 ( .A(n_1048), .B(n_1063), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1050), .Y(n_1048) );
OAI21xp33_ASAP7_75t_L g1051 ( .A1(n_1052), .A2(n_1054), .B(n_1058), .Y(n_1051) );
AOI21xp5_ASAP7_75t_L g1204 ( .A1(n_1052), .A2(n_1159), .B(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx3_ASAP7_75t_L g1179 ( .A(n_1053), .Y(n_1179) );
INVxp67_ASAP7_75t_SL g1054 ( .A(n_1055), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1056), .B(n_1183), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1057), .B(n_1084), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1119 ( .A(n_1057), .B(n_1075), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1057), .B(n_1128), .Y(n_1165) );
AND2x2_ASAP7_75t_SL g1175 ( .A(n_1057), .B(n_1081), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1057), .B(n_1093), .Y(n_1184) );
OAI21xp5_ASAP7_75t_L g1058 ( .A1(n_1059), .A2(n_1071), .B(n_1074), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1062), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1061), .B(n_1081), .Y(n_1093) );
NOR2xp33_ASAP7_75t_L g1120 ( .A(n_1061), .B(n_1112), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1061), .B(n_1108), .Y(n_1145) );
NOR2x1p5_ASAP7_75t_L g1169 ( .A(n_1061), .B(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1061), .Y(n_1194) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1062), .Y(n_1155) );
INVx3_ASAP7_75t_L g1072 ( .A(n_1063), .Y(n_1072) );
INVx2_ASAP7_75t_L g1087 ( .A(n_1063), .Y(n_1087) );
OR2x2_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1066), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_1067), .A2(n_1068), .B1(n_1069), .B2(n_1070), .Y(n_1066) );
AOI322xp5_ASAP7_75t_L g1231 ( .A1(n_1071), .A2(n_1078), .A3(n_1086), .B1(n_1120), .B2(n_1206), .C1(n_1232), .C2(n_1233), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1073), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1072), .B(n_1097), .Y(n_1096) );
NOR2xp33_ASAP7_75t_L g1131 ( .A(n_1072), .B(n_1132), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1072), .B(n_1083), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1072), .B(n_1107), .Y(n_1223) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1073), .Y(n_1107) );
HB1xp67_ASAP7_75t_L g1148 ( .A(n_1073), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1074), .B(n_1128), .Y(n_1138) );
NOR2xp33_ASAP7_75t_L g1174 ( .A(n_1074), .B(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1075), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1075), .B(n_1081), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1075), .B(n_1115), .Y(n_1114) );
A2O1A1Ixp33_ASAP7_75t_L g1076 ( .A1(n_1077), .A2(n_1082), .B(n_1085), .C(n_1089), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
NOR2xp33_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1080), .Y(n_1078) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1080), .Y(n_1102) );
NOR2xp33_ASAP7_75t_L g1118 ( .A(n_1081), .B(n_1119), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1081), .B(n_1092), .Y(n_1122) );
NOR2xp33_ASAP7_75t_L g1151 ( .A(n_1081), .B(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1084), .B(n_1092), .Y(n_1097) );
NOR2xp33_ASAP7_75t_L g1149 ( .A(n_1085), .B(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
NOR2xp33_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1088), .Y(n_1086) );
NOR2xp33_ASAP7_75t_L g1090 ( .A(n_1087), .B(n_1091), .Y(n_1090) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1087), .Y(n_1124) );
BUFx2_ASAP7_75t_L g1183 ( .A(n_1087), .Y(n_1183) );
INVxp67_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1091), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1093), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1092), .B(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1092), .Y(n_1152) );
AOI211xp5_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1098), .B(n_1099), .C(n_1113), .Y(n_1094) );
INVxp67_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1097), .B(n_1124), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1098), .B(n_1169), .Y(n_1168) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1098), .Y(n_1228) );
OAI222xp33_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1103), .B1(n_1105), .B2(n_1109), .C1(n_1110), .C2(n_1112), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
NOR2xp33_ASAP7_75t_L g1226 ( .A(n_1103), .B(n_1171), .Y(n_1226) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
AOI322xp5_ASAP7_75t_L g1188 ( .A1(n_1104), .A2(n_1147), .A3(n_1189), .B1(n_1191), .B2(n_1193), .C1(n_1195), .C2(n_1199), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1108), .Y(n_1105) );
INVx3_ASAP7_75t_L g1176 ( .A(n_1106), .Y(n_1176) );
INVx3_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1108), .B(n_1128), .Y(n_1214) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1111), .B(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1112), .Y(n_1158) );
INVxp67_ASAP7_75t_SL g1113 ( .A(n_1114), .Y(n_1113) );
O2A1O1Ixp33_ASAP7_75t_L g1162 ( .A1(n_1115), .A2(n_1163), .B(n_1164), .C(n_1166), .Y(n_1162) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
AOI221xp5_ASAP7_75t_L g1117 ( .A1(n_1118), .A2(n_1120), .B1(n_1121), .B2(n_1123), .C(n_1125), .Y(n_1117) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
INVxp33_ASAP7_75t_SL g1126 ( .A(n_1127), .Y(n_1126) );
INVx3_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1132), .Y(n_1187) );
INVxp67_ASAP7_75t_SL g1135 ( .A(n_1136), .Y(n_1135) );
NOR2xp33_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1138), .Y(n_1136) );
NAND5xp2_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1172), .C(n_1180), .D(n_1188), .E(n_1201), .Y(n_1139) );
O2A1O1Ixp33_ASAP7_75t_L g1140 ( .A1(n_1141), .A2(n_1149), .B(n_1153), .C(n_1154), .Y(n_1140) );
O2A1O1Ixp33_ASAP7_75t_SL g1141 ( .A1(n_1142), .A2(n_1145), .B(n_1146), .C(n_1148), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
A2O1A1Ixp33_ASAP7_75t_L g1154 ( .A1(n_1155), .A2(n_1156), .B(n_1159), .C(n_1162), .Y(n_1154) );
AOI21xp33_ASAP7_75t_L g1207 ( .A1(n_1155), .A2(n_1193), .B(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
AOI222xp33_ASAP7_75t_L g1172 ( .A1(n_1157), .A2(n_1158), .B1(n_1173), .B2(n_1175), .C1(n_1177), .C2(n_1179), .Y(n_1172) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
OAI31xp33_ASAP7_75t_L g1180 ( .A1(n_1160), .A2(n_1181), .A3(n_1185), .B(n_1187), .Y(n_1180) );
INVxp67_ASAP7_75t_L g1216 ( .A(n_1161), .Y(n_1216) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
CKINVDCx16_ASAP7_75t_R g1209 ( .A(n_1171), .Y(n_1209) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1175), .Y(n_1208) );
INVx3_ASAP7_75t_L g1232 ( .A(n_1176), .Y(n_1232) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1184), .Y(n_1181) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1182), .Y(n_1217) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
AOI211xp5_ASAP7_75t_L g1221 ( .A1(n_1184), .A2(n_1222), .B(n_1224), .C(n_1227), .Y(n_1221) );
INVxp33_ASAP7_75t_SL g1185 ( .A(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
CKINVDCx14_ASAP7_75t_R g1193 ( .A(n_1194), .Y(n_1193) );
INVxp67_ASAP7_75t_SL g1195 ( .A(n_1196), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1198), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1198), .B(n_1206), .Y(n_1205) );
CKINVDCx14_ASAP7_75t_R g1199 ( .A(n_1200), .Y(n_1199) );
AOI21xp33_ASAP7_75t_SL g1227 ( .A1(n_1200), .A2(n_1228), .B(n_1229), .Y(n_1227) );
NAND4xp25_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1210), .C(n_1221), .D(n_1231), .Y(n_1202) );
OAI21xp5_ASAP7_75t_SL g1203 ( .A1(n_1204), .A2(n_1207), .B(n_1209), .Y(n_1203) );
A2O1A1Ixp33_ASAP7_75t_L g1215 ( .A1(n_1208), .A2(n_1216), .B(n_1217), .C(n_1218), .Y(n_1215) );
A2O1A1Ixp33_ASAP7_75t_L g1210 ( .A1(n_1211), .A2(n_1213), .B(n_1215), .C(n_1219), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1212), .B(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
INVxp67_ASAP7_75t_SL g1224 ( .A(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
CKINVDCx5p33_ASAP7_75t_R g1235 ( .A(n_1236), .Y(n_1235) );
INVxp67_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1243), .Y(n_1261) );
NOR2x1_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1255), .Y(n_1243) );
NAND3xp33_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1248), .C(n_1254), .Y(n_1244) );
CKINVDCx16_ASAP7_75t_R g1250 ( .A(n_1251), .Y(n_1250) );
CKINVDCx9p33_ASAP7_75t_R g1252 ( .A(n_1253), .Y(n_1252) );
NAND4xp25_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1257), .C(n_1258), .D(n_1259), .Y(n_1255) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
HB1xp67_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
BUFx2_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
HB1xp67_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
NOR2x1_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1280), .Y(n_1274) );
NAND4xp25_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1277), .C(n_1278), .D(n_1279), .Y(n_1275) );
NAND3xp33_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1283), .C(n_1289), .Y(n_1280) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
BUFx3_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
CKINVDCx5p33_ASAP7_75t_R g1292 ( .A(n_1293), .Y(n_1292) );
endmodule