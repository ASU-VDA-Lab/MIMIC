module fake_jpeg_19963_n_164 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_36),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_20),
.B(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_1),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_23),
.C(n_25),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_47),
.B(n_52),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_30),
.B1(n_20),
.B2(n_18),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_30),
.B1(n_16),
.B2(n_26),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_59),
.B1(n_22),
.B2(n_32),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_24),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_15),
.B1(n_18),
.B2(n_27),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_45),
.B1(n_54),
.B2(n_62),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_33),
.B(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_29),
.Y(n_69)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_77),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_54),
.B1(n_53),
.B2(n_48),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_29),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_87),
.B(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_27),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_82),
.B1(n_50),
.B2(n_19),
.Y(n_103)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_81),
.Y(n_105)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_31),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_41),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_19),
.Y(n_100)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_31),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_15),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_64),
.B1(n_67),
.B2(n_85),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_53),
.B1(n_41),
.B2(n_31),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_96),
.B1(n_80),
.B2(n_74),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_53),
.B1(n_25),
.B2(n_23),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_64),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_84),
.C(n_87),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_103),
.B(n_75),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_78),
.B(n_75),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_102),
.B(n_88),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_115),
.B(n_103),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_71),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_110),
.C(n_120),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_70),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_114),
.C(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_113),
.B(n_92),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_101),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_80),
.B(n_74),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_74),
.B1(n_65),
.B2(n_76),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_97),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_76),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_66),
.C(n_81),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_105),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_123),
.B(n_129),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_94),
.B(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_127),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_95),
.C(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_96),
.B1(n_93),
.B2(n_19),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_109),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_114),
.B1(n_119),
.B2(n_111),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_138),
.B1(n_128),
.B2(n_141),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_140),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_126),
.B(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_105),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_108),
.B1(n_117),
.B2(n_82),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_109),
.B(n_128),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_122),
.B(n_142),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_148),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_138),
.C(n_58),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_5),
.A3(n_9),
.B1(n_7),
.B2(n_14),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_6),
.B(n_13),
.C(n_12),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_R g156 ( 
.A(n_150),
.B(n_9),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_143),
.B(n_146),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_153),
.B(n_149),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_155),
.B(n_156),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_154),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

OAI321xp33_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_151),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_1),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_162),
.A2(n_163),
.B(n_159),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_2),
.B(n_4),
.Y(n_163)
);


endmodule