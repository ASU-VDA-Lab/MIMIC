module fake_netlist_5_93_n_197 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_197);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_197;

wire n_137;
wire n_168;
wire n_164;
wire n_191;
wire n_91;
wire n_82;
wire n_122;
wire n_194;
wire n_142;
wire n_176;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_182;
wire n_143;
wire n_132;
wire n_83;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_189;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_195;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_139;
wire n_38;
wire n_123;
wire n_113;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_30;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_193;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_192;
wire n_53;
wire n_160;
wire n_188;
wire n_190;
wire n_158;
wire n_44;
wire n_154;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_40;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_183;
wire n_185;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_196;
wire n_99;
wire n_181;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_64;
wire n_77;
wire n_106;
wire n_102;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_134;
wire n_187;
wire n_32;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx4_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_27),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_0),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp67_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_R g73 ( 
.A(n_44),
.B(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_71),
.B(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_32),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

OR2x2_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_36),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_46),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_56),
.B(n_72),
.C(n_70),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_67),
.B(n_45),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_67),
.B1(n_41),
.B2(n_39),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_58),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_76),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_74),
.B(n_72),
.C(n_70),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_59),
.B(n_37),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

OAI21x1_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_85),
.B(n_86),
.Y(n_104)
);

OAI21x1_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_86),
.B(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_51),
.B1(n_45),
.B2(n_47),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_92),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_SL g111 ( 
.A(n_109),
.B(n_65),
.C(n_66),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

BUFx4f_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_81),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_81),
.Y(n_115)
);

AO31x2_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_46),
.A3(n_37),
.B(n_47),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_101),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_110),
.B1(n_101),
.B2(n_96),
.Y(n_118)
);

INVxp33_ASAP7_75t_SL g119 ( 
.A(n_112),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_110),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_111),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_116),
.Y(n_124)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_110),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_79),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_116),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_116),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_103),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_111),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

AO21x2_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_105),
.B(n_104),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_128),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_128),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_132),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_136),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_SL g147 ( 
.A(n_136),
.B(n_133),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_132),
.B(n_125),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_134),
.Y(n_149)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_55),
.B1(n_51),
.B2(n_61),
.C(n_93),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_147),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_126),
.B(n_76),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_53),
.B(n_50),
.C(n_150),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_53),
.B(n_50),
.Y(n_161)
);

AOI211xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_74),
.B(n_73),
.C(n_64),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_151),
.A2(n_1),
.B(n_2),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_154),
.B(n_113),
.Y(n_164)
);

OAI211xp5_ASAP7_75t_L g165 ( 
.A1(n_158),
.A2(n_95),
.B(n_100),
.C(n_102),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_113),
.B(n_125),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_149),
.A3(n_103),
.B1(n_87),
.B2(n_78),
.C1(n_8),
.C2(n_9),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_157),
.Y(n_168)
);

AND4x2_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_157),
.C(n_152),
.D(n_5),
.Y(n_169)
);

AOI222xp33_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_83),
.B1(n_89),
.B2(n_87),
.C1(n_78),
.C2(n_90),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_152),
.B1(n_90),
.B2(n_83),
.C(n_91),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_162),
.B(n_165),
.C(n_167),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_125),
.B1(n_137),
.B2(n_83),
.Y(n_174)
);

AND3x4_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_91),
.C(n_92),
.Y(n_175)
);

AOI221xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_40),
.B1(n_2),
.B2(n_6),
.C(n_9),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_172),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_174),
.Y(n_178)
);

AOI221xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_1),
.B1(n_6),
.B2(n_10),
.C(n_11),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_175),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_170),
.A2(n_176),
.B1(n_171),
.B2(n_137),
.Y(n_182)
);

NAND4xp75_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_12),
.C(n_13),
.D(n_108),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_12),
.B1(n_13),
.B2(n_92),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_137),
.B(n_105),
.Y(n_189)
);

OAI22x1_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_182),
.B1(n_183),
.B2(n_108),
.Y(n_190)
);

AO22x2_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_108),
.B1(n_106),
.B2(n_18),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_185),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_189),
.B1(n_184),
.B2(n_106),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_193),
.A2(n_105),
.B1(n_104),
.B2(n_98),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_196),
.A2(n_195),
.B1(n_194),
.B2(n_104),
.Y(n_197)
);


endmodule