module fake_aes_7675_n_21 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_21;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
AOI22xp33_ASAP7_75t_L g11 ( .A1(n_1), .A2(n_4), .B1(n_2), .B2(n_7), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
INVx4_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
NAND2xp5_ASAP7_75t_SL g14 ( .A(n_5), .B(n_8), .Y(n_14) );
AOI21xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_6), .B(n_10), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_15), .B(n_13), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
AOI222xp33_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_11), .B1(n_16), .B2(n_12), .C1(n_13), .C2(n_0), .Y(n_18) );
NAND4xp75_ASAP7_75t_L g19 ( .A(n_18), .B(n_1), .C(n_2), .D(n_3), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_19), .B(n_12), .Y(n_20) );
AOI22x1_ASAP7_75t_SL g21 ( .A1(n_20), .A2(n_3), .B1(n_4), .B2(n_12), .Y(n_21) );
endmodule