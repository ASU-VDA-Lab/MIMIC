module fake_jpeg_29089_n_63 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_31),
.B1(n_34),
.B2(n_4),
.Y(n_36)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_27),
.B1(n_25),
.B2(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_5),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_7),
.B1(n_10),
.B2(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_14),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_6),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_7),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_29),
.C(n_34),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_20),
.C(n_21),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_33),
.B1(n_8),
.B2(n_9),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_48),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_40),
.B(n_43),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_55),
.C(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_44),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_22),
.C(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_52),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_60),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_61),
.Y(n_63)
);


endmodule