module real_jpeg_8822_n_16 (n_5, n_4, n_8, n_0, n_12, n_324, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_324;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_1),
.A2(n_33),
.B1(n_49),
.B2(n_50),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_1),
.A2(n_33),
.B1(n_65),
.B2(n_66),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_2),
.A2(n_50),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_2),
.B(n_50),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_2),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_2),
.A2(n_89),
.B1(n_92),
.B2(n_182),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_2),
.B(n_104),
.Y(n_228)
);

AOI21xp33_ASAP7_75t_L g246 ( 
.A1(n_2),
.A2(n_25),
.B(n_27),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_180),
.Y(n_261)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_4),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g46 ( 
.A(n_7),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_8),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_8),
.A2(n_36),
.B1(n_65),
.B2(n_66),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_10),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_162),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_162),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_162),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_11),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_11),
.A2(n_65),
.B1(n_66),
.B2(n_171),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_171),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_171),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_54),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_12),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_13),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_144),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_144),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_144),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_15),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_71),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_71),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_122),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_20),
.B(n_105),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.C(n_85),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_21),
.A2(n_73),
.B1(n_74),
.B2(n_150),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_21),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_40),
.B2(n_41),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_22),
.A2(n_23),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_23),
.B(n_59),
.C(n_72),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_29),
.B(n_32),
.C(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_24),
.A2(n_30),
.B1(n_38),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_24),
.A2(n_38),
.B1(n_263),
.B2(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_24),
.A2(n_38),
.B1(n_143),
.B2(n_272),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_24)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_27),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_45),
.Y(n_47)
);

HAxp5_ASAP7_75t_SL g205 ( 
.A(n_27),
.B(n_180),
.CON(n_205),
.SN(n_205)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_29),
.A2(n_32),
.B(n_180),
.C(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_35),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_37),
.A2(n_104),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_38),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_38),
.A2(n_143),
.B(n_145),
.Y(n_142)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_59),
.B1(n_60),
.B2(n_72),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_52),
.B(n_55),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_43),
.A2(n_58),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_43),
.A2(n_58),
.B1(n_223),
.B2(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_43),
.A2(n_114),
.B(n_259),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_48),
.B1(n_53),
.B2(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_44),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_44),
.A2(n_48),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_44),
.A2(n_56),
.B(n_115),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_45),
.B(n_50),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_47),
.A2(n_49),
.B1(n_205),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_115),
.Y(n_114)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_62),
.Y(n_63)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_58),
.A2(n_77),
.B(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_58),
.B(n_180),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_59),
.A2(n_60),
.B1(n_113),
.B2(n_118),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_64),
.B(n_69),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_61),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_61),
.A2(n_64),
.B1(n_96),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_61),
.A2(n_64),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_61),
.A2(n_64),
.B1(n_170),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_61),
.A2(n_64),
.B1(n_195),
.B2(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_61),
.A2(n_79),
.B(n_203),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_63),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_64),
.B(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_64),
.A2(n_81),
.B(n_140),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_65),
.B(n_68),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_65),
.B(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_66),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_172)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_70),
.A2(n_84),
.B(n_98),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_74),
.A2(n_75),
.B(n_78),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_85),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_99),
.B(n_100),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_86),
.A2(n_87),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_95),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_99),
.B1(n_100),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_88),
.A2(n_95),
.B1(n_99),
.B2(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B(n_93),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_89),
.A2(n_92),
.B1(n_161),
.B2(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_89),
.A2(n_138),
.B(n_164),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_89),
.A2(n_93),
.B(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_89),
.A2(n_92),
.B1(n_227),
.B2(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_89),
.A2(n_213),
.B(n_249),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_90),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_90),
.A2(n_91),
.B1(n_160),
.B2(n_163),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_91),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_94),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_91),
.B(n_137),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_92),
.B(n_180),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_92),
.A2(n_136),
.B(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_95),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_102),
.B(n_104),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_120),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_119),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_151),
.B(n_322),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_148),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_124),
.B(n_148),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.C(n_132),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_131),
.Y(n_314)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_132),
.A2(n_133),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_141),
.C(n_146),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_134),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_135),
.B(n_139),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_141),
.A2(n_142),
.B1(n_146),
.B2(n_147),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

AOI321xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_298),
.A3(n_310),
.B1(n_315),
.B2(n_321),
.C(n_324),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_265),
.C(n_294),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_239),
.B(n_264),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_216),
.B(n_238),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_198),
.B(n_215),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_189),
.B(n_197),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_177),
.B(n_188),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_159),
.B(n_165),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_172),
.B2(n_176),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_166),
.B(n_176),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_169),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_172),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_183),
.B(n_187),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_190),
.B(n_191),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_192),
.B(n_199),
.Y(n_215)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.CI(n_196),
.CON(n_192),
.SN(n_192)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_209),
.B2(n_214),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_204),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_208),
.C(n_214),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_206),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_209),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_212),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_218),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_232),
.B2(n_233),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_235),
.C(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_224),
.B1(n_225),
.B2(n_231),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_221),
.Y(n_231)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_226),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_228),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_229),
.C(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_234),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_235),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_241),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_253),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_243),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_243),
.B(n_252),
.C(n_253),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_248),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_248),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_250),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_260),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_257),
.C(n_260),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_281),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_266),
.B(n_281),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_275),
.C(n_279),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_297),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_270),
.C(n_274),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_273),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_278),
.Y(n_284)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_290),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_290),
.C(n_291),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_284),
.B(n_286),
.C(n_289),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_296),
.Y(n_318)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_299),
.A2(n_316),
.B(n_320),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_300),
.B(n_301),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_309),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_307),
.C(n_309),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_312),
.Y(n_321)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B(n_319),
.Y(n_316)
);


endmodule