module real_jpeg_13297_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_4),
.A2(n_26),
.B1(n_28),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_83),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_83),
.Y(n_148)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_56),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_8),
.A2(n_27),
.B1(n_68),
.B2(n_69),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_8),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_8),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_26),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_10),
.A2(n_38),
.B1(n_49),
.B2(n_50),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_92),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_14),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_15),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_15),
.B(n_50),
.C(n_89),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_71),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_15),
.A2(n_46),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_15),
.B(n_123),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_116),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_114),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_96),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_19),
.B(n_96),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_58),
.B2(n_59),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_45),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_23),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_34),
.B2(n_37),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_25),
.A2(n_30),
.B1(n_112),
.B2(n_123),
.Y(n_122)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_28),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_26),
.A2(n_43),
.B(n_67),
.C(n_72),
.Y(n_66)
);

HAxp5_ASAP7_75t_SL g112 ( 
.A(n_26),
.B(n_71),
.CON(n_112),
.SN(n_112)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_26),
.B(n_33),
.C(n_36),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_44),
.C(n_68),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_29),
.A2(n_34),
.B1(n_37),
.B2(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

OA22x2_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_32),
.A2(n_35),
.B(n_112),
.C(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_35),
.A2(n_36),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_35),
.B(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_39),
.A2(n_40),
.B1(n_45),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_67),
.B1(n_75),
.B2(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_77),
.Y(n_76)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_44),
.B1(n_68),
.B2(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B(n_53),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_55),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_46),
.B(n_71),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_46),
.A2(n_146),
.B1(n_154),
.B2(n_155),
.Y(n_158)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_49),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_47),
.A2(n_57),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_47),
.B(n_109),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_50),
.B1(n_87),
.B2(n_89),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_49),
.B(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_57),
.Y(n_155)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.CON(n_67),
.SN(n_67)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_71),
.B(n_143),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_95),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_91),
.B(n_93),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_85),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_85),
.A2(n_126),
.B1(n_142),
.B2(n_143),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_SL g89 ( 
.A(n_87),
.Y(n_89)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_102),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.C(n_105),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_105),
.B1(n_106),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_131),
.B(n_178),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_128),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_128),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_124),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_119),
.A2(n_120),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_124),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_172),
.B(n_177),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_161),
.B(n_171),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_149),
.B(n_160),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_144),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_155),
.B(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_156),
.B(n_159),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_158),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_163),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_176),
.Y(n_177)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);


endmodule