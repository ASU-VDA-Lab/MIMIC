module real_jpeg_18807_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_596;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_586;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_612),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_0),
.B(n_613),
.Y(n_612)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_1),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_1),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_1),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_1),
.Y(n_449)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_2),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_3),
.A2(n_62),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_3),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_3),
.A2(n_245),
.B1(n_272),
.B2(n_274),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g462 ( 
.A1(n_3),
.A2(n_245),
.B1(n_463),
.B2(n_465),
.Y(n_462)
);

OAI22xp33_ASAP7_75t_L g521 ( 
.A1(n_3),
.A2(n_245),
.B1(n_522),
.B2(n_525),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_4),
.A2(n_312),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_4),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_4),
.A2(n_314),
.B1(n_387),
.B2(n_392),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_4),
.A2(n_314),
.B1(n_514),
.B2(n_517),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_4),
.A2(n_314),
.B1(n_555),
.B2(n_558),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_5),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_5),
.A2(n_33),
.B1(n_230),
.B2(n_233),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_5),
.A2(n_33),
.B1(n_297),
.B2(n_300),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_5),
.A2(n_33),
.B1(n_335),
.B2(n_338),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_6),
.A2(n_61),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_6),
.A2(n_61),
.B1(n_203),
.B2(n_206),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_6),
.A2(n_61),
.B1(n_233),
.B2(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_7),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_7),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_7),
.A2(n_96),
.B1(n_143),
.B2(n_147),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_7),
.A2(n_96),
.B1(n_255),
.B2(n_257),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_7),
.A2(n_59),
.B1(n_96),
.B2(n_343),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_8),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_8),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_8),
.A2(n_108),
.B1(n_153),
.B2(n_157),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_8),
.A2(n_108),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_8),
.A2(n_108),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_9),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_9),
.Y(n_95)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_9),
.Y(n_223)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_9),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_9),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_9),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_10),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_10),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_10),
.Y(n_253)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_10),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_11),
.A2(n_238),
.B1(n_239),
.B2(n_241),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_11),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_11),
.A2(n_241),
.B1(n_366),
.B2(n_371),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_11),
.A2(n_241),
.B1(n_455),
.B2(n_461),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_11),
.A2(n_241),
.B1(n_537),
.B2(n_540),
.Y(n_536)
);

OAI32xp33_ASAP7_75t_L g278 ( 
.A1(n_12),
.A2(n_279),
.A3(n_283),
.B1(n_285),
.B2(n_291),
.Y(n_278)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_12),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_12),
.A2(n_59),
.B1(n_290),
.B2(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_12),
.B(n_43),
.Y(n_397)
);

OAI32xp33_ASAP7_75t_L g434 ( 
.A1(n_12),
.A2(n_335),
.A3(n_435),
.B1(n_440),
.B2(n_443),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_12),
.A2(n_290),
.B1(n_470),
.B2(n_472),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g531 ( 
.A(n_12),
.B(n_116),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_12),
.B(n_212),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_12),
.B(n_67),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_13),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_15),
.Y(n_135)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_16),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_16),
.Y(n_259)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_181),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_179),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_172),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_22),
.B(n_172),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_150),
.C(n_159),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_23),
.A2(n_150),
.B1(n_590),
.B2(n_591),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_23),
.Y(n_590)
);

XNOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_65),
.Y(n_23)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_24),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_34),
.B1(n_55),
.B2(n_64),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_25),
.A2(n_64),
.B(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_29),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_30),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_31),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_32),
.Y(n_238)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_32),
.Y(n_345)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_34),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_34),
.A2(n_55),
.B(n_174),
.Y(n_173)
);

OAI22x1_ASAP7_75t_SL g236 ( 
.A1(n_34),
.A2(n_64),
.B1(n_237),
.B2(n_242),
.Y(n_236)
);

OAI21x1_ASAP7_75t_L g340 ( 
.A1(n_34),
.A2(n_242),
.B(n_341),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_34),
.A2(n_64),
.B1(n_311),
.B2(n_359),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_34),
.A2(n_174),
.B(n_417),
.Y(n_416)
);

OR2x6_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_43),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_39),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_39),
.Y(n_363)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_40),
.Y(n_284)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_43),
.B(n_152),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_43),
.A2(n_158),
.B1(n_310),
.B2(n_317),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_43),
.B(n_342),
.Y(n_341)
);

AO22x2_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_51),
.B2(n_53),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_45),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_49),
.Y(n_164)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_50),
.Y(n_337)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_52),
.Y(n_139)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_60),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_62),
.B(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_102),
.B1(n_103),
.B2(n_149),
.Y(n_65)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_66),
.B(n_150),
.C(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_66),
.B(n_160),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_78),
.B(n_90),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_67),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_67),
.B(n_221),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_67),
.A2(n_78),
.B1(n_510),
.B2(n_513),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_67),
.A2(n_78),
.B1(n_454),
.B2(n_513),
.Y(n_530)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_68),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_68),
.B(n_91),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_68),
.A2(n_263),
.B1(n_453),
.B2(n_462),
.Y(n_452)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_71),
.Y(n_205)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_71),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_71),
.Y(n_218)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_71),
.Y(n_527)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_75),
.Y(n_208)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_75),
.Y(n_256)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_75),
.Y(n_496)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_75),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_78),
.B(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_78),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_78),
.A2(n_413),
.B(n_477),
.Y(n_476)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_84),
.B2(n_87),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_80),
.Y(n_504)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_82),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_82),
.Y(n_512)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AO22x2_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_117),
.B1(n_120),
.B2(n_123),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_89),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_89),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_89),
.Y(n_518)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g357 ( 
.A1(n_91),
.A2(n_263),
.B(n_327),
.Y(n_357)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_94),
.Y(n_227)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_102),
.B(n_149),
.C(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AO21x1_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_114),
.B(n_140),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_104),
.B(n_116),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_104),
.Y(n_333)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_114),
.A2(n_161),
.B(n_170),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_114),
.A2(n_116),
.B(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_114),
.A2(n_140),
.B(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_114),
.A2(n_116),
.B1(n_161),
.B2(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_115),
.A2(n_142),
.B(n_171),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_115),
.A2(n_141),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_115),
.A2(n_141),
.B1(n_271),
.B2(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_115),
.A2(n_141),
.B1(n_365),
.B2(n_386),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_115),
.A2(n_141),
.B1(n_386),
.B2(n_469),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_128),
.Y(n_115)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_121),
.Y(n_232)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_122),
.Y(n_267)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_132),
.B1(n_136),
.B2(n_138),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_135),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_135),
.Y(n_289)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_138),
.Y(n_276)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_146),
.Y(n_370)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_150),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_150),
.A2(n_591),
.B1(n_595),
.B2(n_596),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_158),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_155),
.Y(n_313)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_159),
.B(n_589),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_163),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_169),
.Y(n_273)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_169),
.Y(n_374)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g615 ( 
.A(n_172),
.Y(n_615)
);

FAx1_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_175),
.CI(n_177),
.CON(n_172),
.SN(n_172)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_586),
.B(n_609),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_423),
.Y(n_183)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_349),
.B(n_400),
.C(n_401),
.D(n_422),
.Y(n_184)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_185),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_318),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_186),
.B(n_318),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_247),
.C(n_268),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_188),
.A2(n_247),
.B1(n_248),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_188),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_235),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_189),
.B(n_236),
.C(n_246),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_219),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_190),
.B(n_219),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_202),
.B(n_209),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_191),
.A2(n_202),
.B1(n_296),
.B2(n_304),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_191),
.A2(n_209),
.B(n_451),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_191),
.A2(n_535),
.B1(n_545),
.B2(n_546),
.Y(n_534)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_192),
.B(n_214),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_192),
.A2(n_254),
.B(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_192),
.A2(n_521),
.B(n_528),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_192),
.A2(n_212),
.B1(n_290),
.B2(n_554),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_192),
.A2(n_536),
.B1(n_554),
.B2(n_568),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_195),
.Y(n_539)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_196),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_197),
.Y(n_544)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_198),
.Y(n_569)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_208),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_218),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_228),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g412 ( 
.A(n_220),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_223),
.Y(n_442)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_234),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_246),
.Y(n_235)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_261),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_249),
.B(n_261),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_260),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_250),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_251),
.Y(n_399)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_254),
.Y(n_451)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_259),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_260),
.A2(n_296),
.B(n_399),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g326 ( 
.A1(n_263),
.A2(n_264),
.B(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_268),
.B(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_277),
.C(n_309),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_269),
.B(n_309),
.Y(n_355)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_277),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_295),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_278),
.B(n_295),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_282),
.Y(n_391)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_290),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_289),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_290),
.B(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_290),
.B(n_503),
.Y(n_502)
);

OAI21xp33_ASAP7_75t_SL g510 ( 
.A1(n_290),
.A2(n_502),
.B(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_303),
.Y(n_524)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_308),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_319),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_329),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_320),
.B(n_329),
.C(n_346),
.Y(n_403)
);

OAI22xp33_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_325),
.B1(n_326),
.B2(n_328),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_321),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_321),
.A2(n_328),
.B1(n_416),
.B2(n_418),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_321),
.B(n_326),
.Y(n_419)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI21xp33_ASAP7_75t_L g600 ( 
.A1(n_328),
.A2(n_418),
.B(n_601),
.Y(n_600)
);

XNOR2x1_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_330),
.B(n_340),
.C(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_340),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_334),
.Y(n_410)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_337),
.Y(n_339)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_342),
.Y(n_417)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.C(n_376),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_350),
.B(n_353),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.C(n_375),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_375),
.Y(n_378)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.C(n_364),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_364),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_377),
.B(n_379),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_382),
.C(n_384),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_380),
.B(n_583),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_382),
.A2(n_383),
.B1(n_384),
.B2(n_584),
.Y(n_583)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_384),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_396),
.C(n_398),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_385),
.B(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_387),
.Y(n_472)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_393),
.Y(n_471)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_396),
.A2(n_397),
.B1(n_398),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_398),
.Y(n_481)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

NOR3xp33_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_425),
.C(n_428),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_404),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_407),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_405),
.B(n_420),
.C(n_604),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_414),
.B1(n_420),
.B2(n_421),
.Y(n_407)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_408),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_409),
.B(n_411),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_414),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_414),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_419),
.Y(n_414)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_416),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g601 ( 
.A(n_419),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_429),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_580),
.B(n_585),
.Y(n_429)
);

AOI21x1_ASAP7_75t_SL g430 ( 
.A1(n_431),
.A2(n_483),
.B(n_579),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_473),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_432),
.B(n_473),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_452),
.C(n_468),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_433),
.B(n_576),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_450),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_434),
.B(n_450),
.Y(n_475)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_439),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_446),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_452),
.B(n_468),
.Y(n_576)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_462),
.Y(n_477)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_478),
.B1(n_479),
.B2(n_482),
.Y(n_473)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_474),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_475),
.B(n_476),
.C(n_478),
.Y(n_581)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_484),
.A2(n_574),
.B(n_578),
.Y(n_483)
);

AOI21x1_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_532),
.B(n_573),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_519),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_486),
.B(n_519),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_508),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_487),
.A2(n_508),
.B1(n_509),
.B2(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_487),
.Y(n_550)
);

OAI32xp33_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_493),
.A3(n_497),
.B1(n_502),
.B2(n_505),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx8_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_529),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_520),
.B(n_530),
.C(n_531),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_521),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_531),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_533),
.A2(n_551),
.B(n_572),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_549),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_534),
.B(n_549),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_552),
.A2(n_566),
.B(n_571),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_553),
.B(n_561),
.Y(n_552)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_562),
.B(n_563),
.Y(n_561)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_567),
.B(n_570),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_567),
.B(n_570),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

NOR2xp67_ASAP7_75t_SL g574 ( 
.A(n_575),
.B(n_577),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_575),
.B(n_577),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_581),
.B(n_582),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_581),
.B(n_582),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_587),
.B(n_602),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_587),
.A2(n_610),
.B(n_611),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_SL g587 ( 
.A(n_588),
.B(n_592),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_588),
.B(n_592),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_593),
.B(n_597),
.C(n_599),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_594),
.A2(n_597),
.B1(n_598),
.B2(n_608),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_594),
.Y(n_608)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_595),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_599),
.A2(n_600),
.B1(n_606),
.B2(n_607),
.Y(n_605)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_603),
.B(n_605),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_603),
.B(n_605),
.Y(n_610)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);


endmodule