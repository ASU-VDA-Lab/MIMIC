module fake_aes_3609_n_520 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_520);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_520;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g75 ( .A(n_50), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_22), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_16), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_67), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_9), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_65), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_13), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_9), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_27), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_71), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_30), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_32), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_68), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_47), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_25), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_42), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_41), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_55), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_45), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_34), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_43), .Y(n_95) );
OR2x2_ASAP7_75t_L g96 ( .A(n_63), .B(n_18), .Y(n_96) );
INVx1_ASAP7_75t_SL g97 ( .A(n_70), .Y(n_97) );
BUFx10_ASAP7_75t_L g98 ( .A(n_62), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_72), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_15), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_60), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_39), .Y(n_102) );
BUFx10_ASAP7_75t_L g103 ( .A(n_1), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_19), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_44), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_52), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_21), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_69), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_87), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_86), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_86), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g112 ( .A(n_98), .B(n_0), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_87), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_100), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_103), .B(n_0), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_76), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_86), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_77), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_83), .Y(n_119) );
INVxp33_ASAP7_75t_SL g120 ( .A(n_92), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_88), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_86), .Y(n_122) );
INVx2_ASAP7_75t_SL g123 ( .A(n_98), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_79), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_89), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_98), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_75), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_100), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_103), .B(n_1), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_126), .B(n_81), .Y(n_131) );
INVx4_ASAP7_75t_L g132 ( .A(n_126), .Y(n_132) );
INVx2_ASAP7_75t_SL g133 ( .A(n_126), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_127), .Y(n_134) );
AND2x6_ASAP7_75t_L g135 ( .A(n_115), .B(n_102), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_126), .B(n_92), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_127), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_127), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_124), .B(n_103), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_123), .B(n_116), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_127), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_123), .B(n_95), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_120), .B(n_91), .Y(n_144) );
OR2x2_ASAP7_75t_L g145 ( .A(n_124), .B(n_82), .Y(n_145) );
AND2x6_ASAP7_75t_L g146 ( .A(n_115), .B(n_101), .Y(n_146) );
NAND2xp33_ASAP7_75t_SL g147 ( .A(n_130), .B(n_105), .Y(n_147) );
AO21x2_ASAP7_75t_L g148 ( .A1(n_112), .A2(n_99), .B(n_104), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_116), .B(n_108), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_127), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_110), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_117), .Y(n_152) );
INVx4_ASAP7_75t_SL g153 ( .A(n_110), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_110), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_141), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_141), .B(n_130), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_141), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_137), .Y(n_159) );
INVxp67_ASAP7_75t_L g160 ( .A(n_139), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_141), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_139), .A2(n_105), .B1(n_118), .B2(n_125), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_135), .A2(n_129), .B1(n_118), .B2(n_125), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_132), .B(n_119), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_150), .Y(n_165) );
INVx4_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_135), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_143), .B(n_119), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_135), .Y(n_170) );
BUFx4f_ASAP7_75t_L g171 ( .A(n_135), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_131), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_132), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_131), .B(n_129), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_135), .A2(n_121), .B1(n_75), .B2(n_107), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_147), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_132), .B(n_121), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_131), .B(n_106), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_131), .B(n_78), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
BUFx2_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
NAND2x1p5_ASAP7_75t_L g182 ( .A(n_133), .B(n_96), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_136), .A2(n_108), .B(n_85), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_145), .B(n_80), .Y(n_184) );
NAND3xp33_ASAP7_75t_SL g185 ( .A(n_144), .B(n_114), .C(n_128), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_145), .B(n_84), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_160), .B(n_109), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_165), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_168), .A2(n_149), .B(n_85), .C(n_94), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_156), .A2(n_135), .B1(n_146), .B2(n_148), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_165), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_165), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_173), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_173), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_167), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_166), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_164), .A2(n_148), .B(n_138), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_174), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_167), .Y(n_201) );
BUFx4f_ASAP7_75t_L g202 ( .A(n_170), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_161), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_174), .B(n_146), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_171), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_162), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_176), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_177), .A2(n_148), .B(n_138), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_174), .B(n_113), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_157), .B(n_146), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_165), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_184), .B(n_146), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_176), .B(n_146), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_156), .B(n_146), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_165), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_172), .A2(n_78), .B(n_94), .C(n_107), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_187), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_166), .Y(n_218) );
AO31x2_ASAP7_75t_L g219 ( .A1(n_190), .A2(n_183), .A3(n_122), .B(n_117), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_194), .Y(n_220) );
BUFx2_ASAP7_75t_SL g221 ( .A(n_215), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_206), .A2(n_146), .B1(n_170), .B2(n_181), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_198), .A2(n_187), .B(n_163), .Y(n_223) );
NAND2x1p5_ASAP7_75t_L g224 ( .A(n_202), .B(n_171), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_194), .Y(n_225) );
OAI22xp33_ASAP7_75t_L g226 ( .A1(n_202), .A2(n_171), .B1(n_181), .B2(n_185), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_200), .B(n_179), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_202), .B(n_166), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_207), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_216), .A2(n_180), .B(n_175), .C(n_179), .Y(n_230) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_208), .A2(n_182), .B(n_180), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_188), .B(n_186), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_199), .B(n_179), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_215), .Y(n_234) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_189), .A2(n_182), .B(n_142), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_199), .B(n_182), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_209), .B(n_178), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_204), .A2(n_97), .B1(n_93), .B2(n_150), .Y(n_238) );
INVxp67_ASAP7_75t_SL g239 ( .A(n_196), .Y(n_239) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_189), .A2(n_140), .B(n_142), .Y(n_240) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_189), .A2(n_134), .B(n_140), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_197), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_203), .B(n_150), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_237), .B(n_209), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_237), .A2(n_203), .B1(n_210), .B2(n_212), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_223), .A2(n_191), .B(n_193), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_220), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_236), .A2(n_195), .B1(n_217), .B2(n_213), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_230), .A2(n_193), .B(n_211), .Y(n_249) );
CKINVDCx11_ASAP7_75t_R g250 ( .A(n_229), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_232), .A2(n_214), .B(n_218), .C(n_197), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_220), .Y(n_252) );
OAI21xp33_ASAP7_75t_L g253 ( .A1(n_236), .A2(n_217), .B(n_193), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_233), .A2(n_195), .B1(n_217), .B2(n_218), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_225), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_233), .B(n_211), .Y(n_256) );
OAI211xp5_ASAP7_75t_SL g257 ( .A1(n_222), .A2(n_122), .B(n_134), .C(n_154), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_229), .B(n_192), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_225), .B(n_197), .Y(n_259) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_228), .A2(n_197), .B1(n_215), .B2(n_201), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_231), .A2(n_192), .B(n_215), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_228), .A2(n_201), .B1(n_196), .B2(n_215), .Y(n_262) );
INVx6_ASAP7_75t_L g263 ( .A(n_234), .Y(n_263) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_227), .A2(n_201), .B1(n_196), .B2(n_122), .C(n_154), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_258), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_247), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_252), .B(n_234), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_255), .B(n_231), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_256), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_259), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_254), .B(n_235), .Y(n_271) );
AO21x2_ASAP7_75t_L g272 ( .A1(n_246), .A2(n_235), .B(n_241), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_254), .B(n_221), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_259), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_244), .B(n_221), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_263), .Y(n_276) );
NOR4xp25_ASAP7_75t_SL g277 ( .A(n_253), .B(n_239), .C(n_219), .D(n_226), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_263), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_263), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_262), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_248), .B(n_219), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_260), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_245), .B(n_219), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_245), .B(n_242), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_248), .B(n_219), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_266), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_269), .B(n_251), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_269), .B(n_219), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_266), .Y(n_289) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_272), .A2(n_261), .B(n_249), .Y(n_290) );
NOR2x1_ASAP7_75t_SL g291 ( .A(n_273), .B(n_260), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_266), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_268), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_268), .Y(n_294) );
NOR2xp67_ASAP7_75t_L g295 ( .A(n_282), .B(n_242), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_285), .B(n_2), .Y(n_296) );
INVx4_ASAP7_75t_L g297 ( .A(n_268), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_285), .B(n_2), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_283), .B(n_3), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_268), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_267), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_272), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_283), .B(n_3), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_265), .B(n_250), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_267), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_271), .B(n_4), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_275), .B(n_228), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_271), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_279), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_281), .B(n_4), .Y(n_310) );
OAI33xp33_ASAP7_75t_L g311 ( .A1(n_281), .A2(n_238), .A3(n_257), .B1(n_7), .B2(n_8), .B3(n_10), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_273), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_272), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_274), .B(n_5), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_282), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_312), .B(n_282), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_297), .B(n_282), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_299), .B(n_284), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_286), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_308), .B(n_280), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_286), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_311), .A2(n_275), .B1(n_274), .B2(n_270), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_297), .B(n_274), .Y(n_323) );
OAI33xp33_ASAP7_75t_L g324 ( .A1(n_310), .A2(n_270), .A3(n_278), .B1(n_276), .B2(n_8), .B3(n_10), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_312), .B(n_277), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_289), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_308), .B(n_277), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_299), .B(n_278), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_310), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_303), .B(n_278), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_289), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_288), .B(n_276), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_300), .B(n_267), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_304), .B(n_5), .Y(n_334) );
NAND4xp25_ASAP7_75t_L g335 ( .A(n_296), .B(n_276), .C(n_267), .D(n_264), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_292), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_297), .B(n_6), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_303), .B(n_6), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_309), .B(n_7), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_292), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_302), .Y(n_341) );
NAND2x1_ASAP7_75t_L g342 ( .A(n_297), .B(n_111), .Y(n_342) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_307), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_309), .B(n_11), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_306), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_300), .B(n_111), .Y(n_346) );
INVx1_ASAP7_75t_SL g347 ( .A(n_314), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_293), .B(n_111), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_296), .B(n_11), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_302), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_298), .B(n_287), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_298), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_293), .B(n_111), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_293), .B(n_111), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_294), .B(n_111), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_294), .B(n_12), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_294), .B(n_110), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_302), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_320), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_320), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_316), .B(n_315), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_329), .B(n_314), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_352), .B(n_301), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_353), .B(n_301), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_321), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_316), .B(n_315), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_345), .B(n_305), .Y(n_368) );
OAI21xp33_ASAP7_75t_L g369 ( .A1(n_334), .A2(n_313), .B(n_315), .Y(n_369) );
OR2x6_ASAP7_75t_L g370 ( .A(n_317), .B(n_295), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_333), .B(n_313), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_351), .B(n_305), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_332), .B(n_313), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_326), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_332), .B(n_305), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_333), .B(n_291), .Y(n_376) );
NAND2x1_ASAP7_75t_L g377 ( .A(n_337), .B(n_305), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_336), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_343), .B(n_290), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_341), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_327), .B(n_291), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_337), .B(n_295), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_327), .B(n_290), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_340), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_325), .B(n_290), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_341), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_319), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_347), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_325), .B(n_110), .Y(n_389) );
INVx4_ASAP7_75t_L g390 ( .A(n_357), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_323), .B(n_110), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_323), .B(n_12), .Y(n_392) );
BUFx2_ASAP7_75t_L g393 ( .A(n_323), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_328), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_338), .B(n_13), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_318), .B(n_152), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_324), .A2(n_344), .B1(n_339), .B2(n_349), .C(n_322), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_317), .B(n_14), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_330), .B(n_152), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_350), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_317), .B(n_17), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_319), .B(n_20), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_350), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_331), .B(n_23), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_331), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_359), .B(n_24), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_357), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_346), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_346), .B(n_26), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_359), .B(n_28), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_388), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_397), .A2(n_335), .B1(n_356), .B2(n_355), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_360), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_361), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_366), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_377), .A2(n_342), .B1(n_358), .B2(n_355), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_374), .Y(n_417) );
OAI21xp5_ASAP7_75t_SL g418 ( .A1(n_369), .A2(n_224), .B(n_356), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_378), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_384), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_364), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_375), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_387), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_381), .B(n_354), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_395), .A2(n_358), .B1(n_354), .B2(n_348), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_373), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_382), .A2(n_342), .B(n_348), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_376), .B(n_29), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_394), .B(n_31), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_382), .A2(n_224), .B1(n_243), .B2(n_240), .Y(n_430) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_392), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g432 ( .A(n_389), .B(n_155), .C(n_151), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_373), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_365), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_405), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_405), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_375), .A2(n_224), .B1(n_205), .B2(n_155), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_371), .Y(n_438) );
OAI221xp5_ASAP7_75t_L g439 ( .A1(n_379), .A2(n_205), .B1(n_155), .B2(n_151), .C(n_37), .Y(n_439) );
AOI322xp5_ASAP7_75t_L g440 ( .A1(n_381), .A2(n_205), .A3(n_155), .B1(n_151), .B2(n_38), .C1(n_40), .C2(n_46), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_407), .B(n_33), .Y(n_441) );
AOI21xp33_ASAP7_75t_L g442 ( .A1(n_389), .A2(n_35), .B(n_36), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_392), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_371), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_383), .B(n_48), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_390), .B(n_241), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_368), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_372), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_390), .A2(n_151), .B1(n_51), .B2(n_53), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_379), .Y(n_450) );
INVxp67_ASAP7_75t_L g451 ( .A(n_391), .Y(n_451) );
AOI21xp33_ASAP7_75t_SL g452 ( .A1(n_370), .A2(n_49), .B(n_54), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_408), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_422), .B(n_376), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_412), .A2(n_385), .B1(n_383), .B2(n_393), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_411), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_415), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_431), .B(n_363), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_421), .B(n_393), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_434), .B(n_390), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_450), .B(n_385), .Y(n_461) );
AOI31xp33_ASAP7_75t_L g462 ( .A1(n_452), .A2(n_443), .A3(n_416), .B(n_427), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_423), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_447), .B(n_362), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_424), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_413), .A2(n_396), .B1(n_367), .B2(n_362), .C(n_391), .Y(n_466) );
AOI211xp5_ASAP7_75t_L g467 ( .A1(n_418), .A2(n_401), .B(n_398), .C(n_367), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_448), .B(n_400), .Y(n_468) );
AOI21xp33_ASAP7_75t_SL g469 ( .A1(n_418), .A2(n_370), .B(n_401), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
OAI211xp5_ASAP7_75t_SL g471 ( .A1(n_440), .A2(n_399), .B(n_409), .C(n_402), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_419), .Y(n_472) );
INVxp67_ASAP7_75t_L g473 ( .A(n_414), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_420), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_451), .B(n_398), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_446), .A2(n_370), .B(n_406), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_438), .B(n_399), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_425), .A2(n_370), .B1(n_400), .B2(n_403), .Y(n_479) );
AOI221x1_ASAP7_75t_L g480 ( .A1(n_449), .A2(n_404), .B1(n_410), .B2(n_406), .C(n_403), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_444), .B(n_386), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_455), .A2(n_424), .B1(n_453), .B2(n_426), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_462), .A2(n_432), .B1(n_428), .B2(n_433), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_463), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_463), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g486 ( .A1(n_469), .A2(n_445), .B1(n_439), .B2(n_430), .C(n_429), .Y(n_486) );
NAND4xp25_ASAP7_75t_L g487 ( .A(n_480), .B(n_432), .C(n_442), .D(n_437), .Y(n_487) );
OAI21xp33_ASAP7_75t_SL g488 ( .A1(n_465), .A2(n_458), .B(n_454), .Y(n_488) );
O2A1O1Ixp5_ASAP7_75t_SL g489 ( .A1(n_456), .A2(n_441), .B(n_436), .C(n_410), .Y(n_489) );
AOI211xp5_ASAP7_75t_L g490 ( .A1(n_479), .A2(n_386), .B(n_380), .C(n_240), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_457), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_470), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g493 ( .A1(n_473), .A2(n_380), .B1(n_169), .B2(n_159), .C(n_59), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_472), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_460), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_477), .A2(n_56), .B(n_57), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_459), .B(n_461), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g498 ( .A1(n_483), .A2(n_467), .B1(n_466), .B2(n_471), .C(n_476), .Y(n_498) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_488), .A2(n_475), .B1(n_478), .B2(n_468), .C(n_471), .Y(n_499) );
AOI21xp33_ASAP7_75t_SL g500 ( .A1(n_484), .A2(n_481), .B(n_464), .Y(n_500) );
XNOR2x1_ASAP7_75t_L g501 ( .A(n_482), .B(n_474), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_485), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_491), .Y(n_503) );
XOR2xp5_ASAP7_75t_L g504 ( .A(n_487), .B(n_58), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_492), .Y(n_505) );
XNOR2xp5_ASAP7_75t_L g506 ( .A(n_495), .B(n_61), .Y(n_506) );
AOI221x1_ASAP7_75t_L g507 ( .A1(n_505), .A2(n_496), .B1(n_487), .B2(n_494), .C(n_497), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_502), .B(n_486), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_499), .A2(n_490), .B1(n_493), .B2(n_489), .C(n_159), .Y(n_509) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_501), .B(n_64), .Y(n_510) );
NOR4xp25_ASAP7_75t_L g511 ( .A(n_508), .B(n_498), .C(n_503), .D(n_504), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_509), .B(n_498), .C(n_500), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_507), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_513), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_511), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_514), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_516), .B(n_515), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_517), .A2(n_510), .B1(n_512), .B2(n_506), .Y(n_518) );
AOI22x1_ASAP7_75t_L g519 ( .A1(n_518), .A2(n_66), .B1(n_73), .B2(n_74), .Y(n_519) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_519), .A2(n_153), .B1(n_169), .B2(n_513), .C1(n_514), .C2(n_515), .Y(n_520) );
endmodule