module fake_jpeg_2055_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_46),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_38),
.B1(n_45),
.B2(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_44),
.Y(n_66)
);

OR2x4_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_2),
.Y(n_94)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_65),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_36),
.B(n_51),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_82),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_50),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_54),
.B1(n_53),
.B2(n_49),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_26),
.B1(n_34),
.B2(n_33),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_41),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_90),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_53),
.B1(n_57),
.B2(n_18),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_1),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_96),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_8),
.B(n_9),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_100),
.B1(n_104),
.B2(n_96),
.Y(n_115)
);

CKINVDCx12_ASAP7_75t_R g102 ( 
.A(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_102),
.B(n_88),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_17),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_106),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_7),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_113),
.Y(n_118)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_111),
.A2(n_112),
.B(n_88),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_8),
.B(n_9),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_113),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_15),
.B(n_22),
.C(n_28),
.D(n_29),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_123),
.C(n_124),
.Y(n_129)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_30),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_126),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_122),
.C(n_107),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_133),
.A2(n_127),
.B1(n_131),
.B2(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_136),
.B(n_118),
.C(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_121),
.B(n_125),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_112),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_125),
.C(n_32),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_31),
.Y(n_143)
);


endmodule