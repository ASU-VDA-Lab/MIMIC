module fake_jpeg_3243_n_680 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_680);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_680;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_19),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_8),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_60),
.Y(n_174)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_63),
.Y(n_193)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_66),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_68),
.Y(n_183)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g202 ( 
.A(n_69),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_70),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_10),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_71),
.A2(n_75),
.B(n_52),
.C(n_6),
.Y(n_182)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_72),
.Y(n_170)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_74),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_35),
.B(n_10),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_79),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_81),
.Y(n_225)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_85),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_34),
.Y(n_86)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_87),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_88),
.B(n_18),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_89),
.Y(n_220)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_29),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g163 ( 
.A1(n_91),
.A2(n_127),
.B1(n_34),
.B2(n_35),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_92),
.Y(n_213)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_20),
.B(n_7),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_57),
.Y(n_148)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_98),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_99),
.Y(n_217)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_109),
.Y(n_206)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_112),
.Y(n_208)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_29),
.Y(n_113)
);

CKINVDCx6p67_ASAP7_75t_R g205 ( 
.A(n_113),
.Y(n_205)
);

BUFx12_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_118),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_22),
.Y(n_119)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_119),
.Y(n_215)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_22),
.Y(n_121)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_121),
.Y(n_227)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_123),
.Y(n_187)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_22),
.Y(n_124)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_125),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_126),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_37),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_22),
.Y(n_128)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_128),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_22),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_129),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_131),
.B(n_14),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_75),
.A2(n_23),
.B1(n_20),
.B2(n_25),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_134),
.A2(n_178),
.B1(n_218),
.B2(n_223),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_24),
.B1(n_49),
.B2(n_39),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_139),
.A2(n_146),
.B1(n_149),
.B2(n_155),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_71),
.A2(n_64),
.B1(n_84),
.B2(n_81),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_148),
.B(n_177),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_62),
.A2(n_23),
.B1(n_25),
.B2(n_44),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_70),
.B(n_57),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_151),
.A2(n_165),
.B(n_172),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_87),
.A2(n_39),
.B1(n_28),
.B2(n_49),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_152),
.A2(n_169),
.B1(n_195),
.B2(n_183),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_66),
.A2(n_36),
.B1(n_44),
.B2(n_55),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_86),
.A2(n_40),
.B1(n_28),
.B2(n_24),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_162),
.A2(n_173),
.B(n_221),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_163),
.A2(n_223),
.B1(n_4),
.B2(n_5),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_98),
.B(n_36),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_104),
.A2(n_34),
.B1(n_40),
.B2(n_42),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_171),
.B(n_182),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_98),
.B(n_11),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_60),
.A2(n_40),
.B1(n_34),
.B2(n_52),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_72),
.B(n_7),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_67),
.A2(n_52),
.B1(n_42),
.B2(n_11),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_90),
.B(n_6),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_181),
.B(n_222),
.Y(n_263)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_191),
.Y(n_315)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_199),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_201),
.B(n_229),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_89),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g219 ( 
.A(n_92),
.B(n_14),
.C(n_13),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_219),
.B(n_5),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_124),
.A2(n_18),
.B1(n_14),
.B2(n_13),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_114),
.B(n_12),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_99),
.A2(n_12),
.B1(n_6),
.B2(n_2),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_132),
.B(n_12),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_228),
.B(n_230),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_68),
.B(n_12),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_74),
.B(n_6),
.Y(n_230)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_233),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_235),
.Y(n_338)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_236),
.Y(n_346)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_237),
.Y(n_325)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_238),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_175),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_239),
.B(n_253),
.Y(n_342)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_141),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_243),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_152),
.A2(n_115),
.B1(n_112),
.B2(n_103),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_244),
.A2(n_268),
.B1(n_285),
.B2(n_291),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_145),
.Y(n_245)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_245),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_SL g247 ( 
.A1(n_163),
.A2(n_91),
.B(n_127),
.C(n_102),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_247),
.A2(n_293),
.B1(n_300),
.B2(n_307),
.Y(n_353)
);

OR2x2_ASAP7_75t_SL g248 ( 
.A(n_148),
.B(n_79),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_248),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_193),
.Y(n_249)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

INVx4_ASAP7_75t_SL g250 ( 
.A(n_140),
.Y(n_250)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_250),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_251),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_191),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_252),
.A2(n_303),
.B(n_273),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_165),
.Y(n_253)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_255),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_135),
.B(n_0),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_257),
.B(n_276),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_196),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_259),
.B(n_260),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_151),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_205),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_261),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_141),
.Y(n_264)
);

INVx8_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_174),
.Y(n_265)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_265),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_164),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_266),
.Y(n_360)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_154),
.Y(n_267)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_230),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_159),
.Y(n_269)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_269),
.Y(n_348)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_176),
.Y(n_270)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_270),
.Y(n_352)
);

INVx11_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_271),
.Y(n_361)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_161),
.Y(n_272)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_193),
.Y(n_273)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_273),
.Y(n_379)
);

INVx4_ASAP7_75t_SL g274 ( 
.A(n_153),
.Y(n_274)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_274),
.Y(n_351)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_166),
.Y(n_275)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_275),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_2),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_184),
.Y(n_277)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_277),
.Y(n_355)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_206),
.Y(n_278)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_278),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_3),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_279),
.B(n_281),
.Y(n_331)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_167),
.Y(n_280)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_280),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_158),
.B(n_4),
.Y(n_281)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_150),
.Y(n_282)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_282),
.Y(n_367)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_144),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_283),
.Y(n_378)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_189),
.Y(n_284)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_284),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_180),
.A2(n_4),
.B1(n_5),
.B2(n_209),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_215),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_287),
.Y(n_322)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_190),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_289),
.Y(n_327)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_212),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g290 ( 
.A(n_185),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_290),
.B(n_295),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_292),
.B(n_297),
.Y(n_358)
);

INVx11_ASAP7_75t_L g293 ( 
.A(n_205),
.Y(n_293)
);

OA22x2_ASAP7_75t_SL g294 ( 
.A1(n_163),
.A2(n_219),
.B1(n_218),
.B2(n_173),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_294),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_156),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_196),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_296),
.B(n_304),
.Y(n_362)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_194),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_211),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_299),
.Y(n_336)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_147),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_167),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_301),
.A2(n_183),
.B1(n_195),
.B2(n_224),
.Y(n_350)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_208),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_302),
.B(n_303),
.Y(n_373)
);

INVx3_ASAP7_75t_SL g303 ( 
.A(n_202),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_133),
.B(n_138),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_202),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_305),
.B(n_309),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_306),
.A2(n_312),
.B1(n_213),
.B2(n_217),
.Y(n_319)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_150),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_177),
.A2(n_181),
.B1(n_143),
.B2(n_160),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_308),
.A2(n_137),
.B1(n_225),
.B2(n_244),
.Y(n_357)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_179),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_174),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_310),
.A2(n_313),
.B1(n_314),
.B2(n_316),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_197),
.A2(n_220),
.B1(n_142),
.B2(n_160),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_136),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_187),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_157),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_172),
.B(n_231),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_200),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_319),
.A2(n_345),
.B1(n_357),
.B2(n_372),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_248),
.B(n_315),
.C(n_241),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_320),
.B(n_356),
.C(n_290),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_330),
.B(n_366),
.Y(n_398)
);

AND2x2_ASAP7_75t_SL g335 ( 
.A(n_315),
.B(n_203),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_335),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_226),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_341),
.B(n_363),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_234),
.A2(n_162),
.B1(n_221),
.B2(n_169),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_350),
.A2(n_364),
.B1(n_293),
.B2(n_271),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_232),
.A2(n_225),
.B1(n_224),
.B2(n_207),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_354),
.A2(n_370),
.B1(n_261),
.B2(n_299),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_256),
.B(n_198),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_263),
.B(n_256),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_301),
.A2(n_308),
.B1(n_232),
.B2(n_254),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_262),
.B(n_292),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_365),
.B(n_358),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_294),
.A2(n_247),
.B1(n_291),
.B2(n_240),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_294),
.A2(n_285),
.B1(n_252),
.B2(n_280),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_380),
.A2(n_386),
.B1(n_388),
.B2(n_389),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_324),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_381),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_342),
.B(n_314),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_382),
.Y(n_459)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_379),
.Y(n_383)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_258),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_384),
.B(n_399),
.C(n_411),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_370),
.A2(n_243),
.B1(n_300),
.B2(n_264),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_379),
.Y(n_387)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_387),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_368),
.A2(n_238),
.B1(n_288),
.B2(n_236),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_368),
.A2(n_242),
.B1(n_246),
.B2(n_297),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_366),
.A2(n_249),
.B(n_289),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_390),
.A2(n_401),
.B(n_403),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_391),
.A2(n_400),
.B1(n_424),
.B2(n_347),
.Y(n_465)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_318),
.Y(n_392)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_392),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_341),
.B(n_363),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_393),
.B(n_413),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_319),
.A2(n_309),
.B1(n_298),
.B2(n_270),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_394),
.A2(n_410),
.B1(n_347),
.B2(n_352),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_324),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_395),
.B(n_404),
.Y(n_450)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_397),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_320),
.B(n_245),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_372),
.A2(n_250),
.B1(n_274),
.B2(n_310),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_358),
.A2(n_235),
.B(n_265),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_402),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_339),
.A2(n_295),
.B(n_251),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_335),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_322),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_405),
.B(n_408),
.Y(n_460)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_375),
.Y(n_406)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_406),
.Y(n_454)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_374),
.Y(n_407)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_407),
.Y(n_457)
);

NAND3xp33_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_290),
.C(n_282),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_322),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_339),
.A2(n_307),
.B1(n_353),
.B2(n_330),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_349),
.B(n_335),
.C(n_326),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_354),
.B(n_362),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_412),
.B(n_327),
.Y(n_432)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_375),
.Y(n_414)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_414),
.Y(n_462)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_326),
.Y(n_415)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_415),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_331),
.B(n_323),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_416),
.B(n_336),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_345),
.A2(n_357),
.B1(n_343),
.B2(n_327),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g455 ( 
.A1(n_417),
.A2(n_346),
.B1(n_367),
.B2(n_344),
.Y(n_455)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_359),
.Y(n_418)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_418),
.Y(n_471)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_419),
.B(n_420),
.Y(n_463)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_374),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_358),
.B(n_376),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_421),
.B(n_373),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_340),
.B(n_333),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_422),
.B(n_423),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_360),
.B(n_355),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_343),
.A2(n_355),
.B1(n_344),
.B2(n_327),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_322),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_425),
.B(n_427),
.Y(n_467)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_328),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_360),
.B(n_361),
.Y(n_428)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_428),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_361),
.B(n_337),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_429),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_432),
.B(n_437),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_446),
.C(n_447),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_389),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_440),
.B(n_441),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_388),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_398),
.A2(n_337),
.B(n_351),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_444),
.A2(n_452),
.B(n_455),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_396),
.B(n_393),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_445),
.B(n_421),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_378),
.C(n_321),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_384),
.B(n_351),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_385),
.A2(n_344),
.B1(n_371),
.B2(n_332),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_449),
.A2(n_461),
.B1(n_464),
.B2(n_465),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_451),
.B(n_416),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_403),
.A2(n_367),
.B(n_346),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_396),
.B(n_321),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_453),
.B(n_458),
.C(n_442),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_409),
.B(n_325),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_385),
.A2(n_332),
.B1(n_334),
.B2(n_325),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_412),
.Y(n_466)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_466),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_456),
.A2(n_424),
.B1(n_386),
.B2(n_380),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_472),
.A2(n_509),
.B1(n_470),
.B2(n_462),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_468),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_473),
.B(n_480),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_466),
.A2(n_400),
.B1(n_390),
.B2(n_412),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_474),
.A2(n_492),
.B1(n_506),
.B2(n_377),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g476 ( 
.A(n_444),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_476),
.B(n_432),
.Y(n_513)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_479),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_463),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_481),
.B(n_484),
.Y(n_542)
);

NOR2x1_ASAP7_75t_SL g482 ( 
.A(n_451),
.B(n_411),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_482),
.Y(n_541)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_430),
.Y(n_483)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_483),
.Y(n_514)
);

AO22x1_ASAP7_75t_L g484 ( 
.A1(n_465),
.A2(n_410),
.B1(n_394),
.B2(n_425),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_434),
.Y(n_485)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_485),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_431),
.A2(n_426),
.B(n_404),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_487),
.A2(n_489),
.B(n_491),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_463),
.Y(n_488)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_488),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_431),
.A2(n_413),
.B(n_392),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_443),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_490),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_460),
.A2(n_401),
.B(n_405),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_456),
.A2(n_445),
.B1(n_440),
.B2(n_441),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_493),
.B(n_438),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_437),
.Y(n_494)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_494),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_498),
.Y(n_516)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_496),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_443),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_497),
.B(n_438),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_442),
.B(n_451),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_460),
.Y(n_499)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_499),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_467),
.B(n_406),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_500),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_452),
.A2(n_395),
.B(n_381),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_501),
.Y(n_543)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_503),
.Y(n_518)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_435),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_458),
.B(n_387),
.C(n_397),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_505),
.C(n_447),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_439),
.B(n_383),
.C(n_415),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_461),
.A2(n_419),
.B1(n_414),
.B2(n_418),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_464),
.A2(n_402),
.B1(n_427),
.B2(n_407),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_453),
.B(n_420),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_510),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_511),
.B(n_519),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_513),
.B(n_537),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_517),
.B(n_481),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_446),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_475),
.B(n_450),
.C(n_459),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_520),
.B(n_524),
.C(n_532),
.Y(n_554)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_522),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_475),
.B(n_450),
.C(n_433),
.Y(n_524)
);

AOI21x1_ASAP7_75t_L g525 ( 
.A1(n_501),
.A2(n_436),
.B(n_470),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_525),
.A2(n_536),
.B(n_538),
.Y(n_552)
);

OAI22x1_ASAP7_75t_L g528 ( 
.A1(n_507),
.A2(n_449),
.B1(n_468),
.B2(n_436),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_528),
.A2(n_484),
.B1(n_474),
.B2(n_477),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_531),
.A2(n_472),
.B1(n_484),
.B2(n_480),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_498),
.B(n_433),
.C(n_454),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_490),
.A2(n_469),
.B1(n_462),
.B2(n_454),
.Y(n_533)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_533),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_497),
.A2(n_448),
.B1(n_471),
.B2(n_468),
.Y(n_535)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_535),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_508),
.A2(n_457),
.B(n_471),
.Y(n_536)
);

INVxp33_ASAP7_75t_SL g537 ( 
.A(n_494),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_508),
.A2(n_457),
.B(n_448),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_478),
.A2(n_328),
.B1(n_352),
.B2(n_378),
.Y(n_540)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_540),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_505),
.B(n_334),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_544),
.B(n_483),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_546),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_504),
.B(n_377),
.C(n_348),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_547),
.B(n_548),
.C(n_510),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_493),
.B(n_348),
.C(n_369),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_550),
.B(n_546),
.Y(n_602)
);

XNOR2x1_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_487),
.Y(n_553)
);

XNOR2x1_ASAP7_75t_L g585 ( 
.A(n_553),
.B(n_569),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_515),
.A2(n_489),
.B(n_491),
.Y(n_555)
);

OAI21x1_ASAP7_75t_SL g599 ( 
.A1(n_555),
.A2(n_560),
.B(n_562),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_519),
.B(n_489),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_557),
.B(n_566),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_558),
.B(n_559),
.Y(n_587)
);

FAx1_ASAP7_75t_L g560 ( 
.A(n_515),
.B(n_482),
.CI(n_492),
.CON(n_560),
.SN(n_560)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_561),
.A2(n_576),
.B1(n_577),
.B2(n_525),
.Y(n_592)
);

FAx1_ASAP7_75t_L g562 ( 
.A(n_542),
.B(n_486),
.CI(n_507),
.CON(n_562),
.SN(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_518),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_563),
.B(n_568),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_516),
.B(n_486),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_518),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_SL g569 ( 
.A(n_517),
.B(n_500),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_570),
.B(n_539),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_516),
.B(n_477),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_571),
.B(n_573),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_511),
.B(n_488),
.C(n_496),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_572),
.B(n_575),
.C(n_578),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_520),
.B(n_478),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_518),
.Y(n_574)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_574),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_524),
.B(n_485),
.C(n_503),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_528),
.A2(n_542),
.B1(n_523),
.B2(n_538),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_523),
.A2(n_506),
.B1(n_509),
.B2(n_479),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_541),
.B(n_502),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_556),
.B(n_554),
.C(n_572),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_581),
.B(n_583),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_556),
.B(n_547),
.C(n_548),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_554),
.B(n_541),
.C(n_543),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_586),
.B(n_588),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_575),
.B(n_543),
.C(n_536),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_551),
.Y(n_589)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_589),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_571),
.B(n_521),
.C(n_534),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_590),
.B(n_593),
.Y(n_611)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_577),
.Y(n_591)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_591),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_592),
.A2(n_603),
.B1(n_604),
.B2(n_562),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_549),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_557),
.B(n_534),
.C(n_529),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_594),
.B(n_597),
.Y(n_613)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_565),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_595),
.B(n_598),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_573),
.B(n_558),
.C(n_566),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_564),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_553),
.B(n_578),
.C(n_555),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_601),
.B(n_579),
.C(n_576),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_602),
.B(n_527),
.Y(n_620)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_561),
.Y(n_603)
);

BUFx24_ASAP7_75t_SL g605 ( 
.A(n_596),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_605),
.B(n_609),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_607),
.B(n_624),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_584),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_599),
.A2(n_562),
.B1(n_560),
.B2(n_530),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_610),
.A2(n_618),
.B1(n_621),
.B2(n_545),
.Y(n_634)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_612),
.Y(n_636)
);

BUFx24_ASAP7_75t_SL g614 ( 
.A(n_587),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_614),
.B(n_583),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_581),
.B(n_552),
.C(n_560),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_616),
.B(n_619),
.C(n_625),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_SL g617 ( 
.A(n_585),
.B(n_559),
.Y(n_617)
);

XNOR2x1_ASAP7_75t_L g633 ( 
.A(n_617),
.B(n_620),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_592),
.A2(n_530),
.B1(n_552),
.B2(n_539),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_580),
.B(n_550),
.C(n_569),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_602),
.A2(n_567),
.B1(n_529),
.B2(n_514),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_586),
.B(n_473),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_600),
.B(n_512),
.Y(n_625)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_622),
.Y(n_627)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_627),
.Y(n_649)
);

INVx11_ASAP7_75t_L g628 ( 
.A(n_611),
.Y(n_628)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_628),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_618),
.B(n_601),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_629),
.B(n_630),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_610),
.B(n_590),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_620),
.A2(n_594),
.B(n_588),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_631),
.A2(n_638),
.B(n_613),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_632),
.B(n_635),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_634),
.A2(n_643),
.B1(n_625),
.B2(n_615),
.Y(n_644)
);

INVx11_ASAP7_75t_L g635 ( 
.A(n_606),
.Y(n_635)
);

INVx11_ASAP7_75t_L g637 ( 
.A(n_621),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_637),
.B(n_338),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_623),
.A2(n_585),
.B(n_580),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_624),
.B(n_526),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_641),
.A2(n_617),
.B(n_369),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_616),
.A2(n_526),
.B1(n_512),
.B2(n_514),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_642),
.B(n_630),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_607),
.A2(n_587),
.B1(n_600),
.B2(n_582),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_644),
.A2(n_647),
.B(n_650),
.Y(n_658)
);

INVxp67_ASAP7_75t_SL g660 ( 
.A(n_646),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g647 ( 
.A(n_632),
.B(n_608),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_639),
.B(n_619),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_636),
.A2(n_545),
.B1(n_582),
.B2(n_597),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_651),
.A2(n_654),
.B1(n_637),
.B2(n_631),
.Y(n_659)
);

NOR2xp67_ASAP7_75t_L g662 ( 
.A(n_652),
.B(n_649),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_653),
.B(n_630),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_636),
.A2(n_329),
.B1(n_338),
.B2(n_634),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_655),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_657),
.B(n_659),
.Y(n_669)
);

O2A1O1Ixp33_ASAP7_75t_SL g661 ( 
.A1(n_656),
.A2(n_628),
.B(n_629),
.C(n_633),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_661),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_662),
.B(n_663),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_SL g663 ( 
.A(n_648),
.B(n_626),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_646),
.B(n_626),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_664),
.B(n_644),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_667),
.A2(n_670),
.B(n_671),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g670 ( 
.A(n_658),
.B(n_650),
.C(n_645),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_L g671 ( 
.A(n_660),
.B(n_640),
.C(n_665),
.Y(n_671)
);

OAI21xp33_ASAP7_75t_L g672 ( 
.A1(n_666),
.A2(n_651),
.B(n_638),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_SL g675 ( 
.A1(n_672),
.A2(n_673),
.B(n_668),
.C(n_629),
.Y(n_675)
);

AOI321xp33_ASAP7_75t_SL g673 ( 
.A1(n_668),
.A2(n_661),
.A3(n_629),
.B1(n_640),
.B2(n_635),
.C(n_643),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_SL g677 ( 
.A1(n_675),
.A2(n_676),
.B(n_641),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g676 ( 
.A(n_674),
.B(n_669),
.C(n_639),
.Y(n_676)
);

BUFx24_ASAP7_75t_SL g678 ( 
.A(n_677),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_678),
.B(n_654),
.C(n_627),
.Y(n_679)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_633),
.C(n_329),
.Y(n_680)
);


endmodule