module fake_netlist_6_4007_n_1332 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1332);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1332;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_532;
wire n_1308;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_814;
wire n_389;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_924;
wire n_475;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_129),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_287),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_222),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_215),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_166),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_212),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_172),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_151),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_291),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_231),
.Y(n_337)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_186),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_240),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_111),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_161),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_97),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_125),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_25),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_81),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_74),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_133),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_5),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_107),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_144),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_206),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_154),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_80),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_16),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_124),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_214),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_273),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_236),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_126),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_216),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_37),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_256),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_292),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_325),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_87),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_40),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_173),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_305),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_103),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_181),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_160),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_178),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_261),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_260),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_297),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_245),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_197),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_146),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_175),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_179),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_69),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_247),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_168),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_293),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_28),
.B(n_99),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_229),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_94),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_290),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_165),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_134),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_283),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_268),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_221),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_180),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_152),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_118),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_243),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_116),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_185),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_278),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_220),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_55),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_284),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_277),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_254),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_140),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_115),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_114),
.Y(n_409)
);

BUFx8_ASAP7_75t_SL g410 ( 
.A(n_158),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_42),
.B(n_207),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_241),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_46),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_187),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_190),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_269),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_170),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_286),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_113),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_322),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_301),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_162),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_272),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_58),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_49),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_282),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_16),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_142),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_137),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_66),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_57),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_237),
.B(n_156),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_44),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_234),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_169),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_182),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_249),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_90),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_8),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_274),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_25),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_17),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_250),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_2),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_53),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_92),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_171),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_72),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_91),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_40),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_65),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_34),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_208),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_128),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_285),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_75),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_223),
.Y(n_458)
);

BUFx10_ASAP7_75t_L g459 ( 
.A(n_82),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_259),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_211),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_10),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_300),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_123),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_188),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_314),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_139),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_218),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_267),
.Y(n_469)
);

NOR2xp67_ASAP7_75t_L g470 ( 
.A(n_46),
.B(n_112),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_202),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_153),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_68),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_77),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_271),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_63),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_58),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_226),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_264),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_302),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_213),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_174),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_219),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_288),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_280),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_317),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_132),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_233),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_2),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_100),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_176),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_217),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_45),
.Y(n_493)
);

BUFx10_ASAP7_75t_L g494 ( 
.A(n_296),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_326),
.B(n_246),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_21),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_84),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_163),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_8),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_96),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_276),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_157),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_1),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_86),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_195),
.Y(n_505)
);

INVxp33_ASAP7_75t_SL g506 ( 
.A(n_85),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_255),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_324),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_88),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_209),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_266),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_238),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_307),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_253),
.Y(n_514)
);

BUFx2_ASAP7_75t_SL g515 ( 
.A(n_194),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_258),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_109),
.Y(n_517)
);

BUFx2_ASAP7_75t_SL g518 ( 
.A(n_159),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_98),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_257),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_51),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_281),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_150),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_59),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_1),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_224),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_225),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_108),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_34),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_306),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_117),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_318),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_198),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_248),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_24),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_0),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_228),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_20),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_104),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_200),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_71),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_167),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_304),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_235),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_361),
.B(n_0),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_538),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_348),
.Y(n_547)
);

OA21x2_ASAP7_75t_L g548 ( 
.A1(n_339),
.A2(n_3),
.B(n_4),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_334),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g550 ( 
.A1(n_341),
.A2(n_3),
.B(n_4),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_538),
.B(n_5),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_379),
.B(n_6),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_334),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_538),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_538),
.B(n_6),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_338),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_453),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_366),
.B(n_7),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_477),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_434),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_348),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_443),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_369),
.B(n_11),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_338),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_334),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_488),
.B(n_418),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_338),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_354),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_344),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_334),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_350),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_377),
.B(n_12),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_436),
.B(n_13),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_336),
.A2(n_61),
.B(n_60),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_338),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_351),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_377),
.B(n_14),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_338),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_440),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_425),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_481),
.B(n_14),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_426),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_428),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_451),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_350),
.Y(n_585)
);

OA21x2_ASAP7_75t_L g586 ( 
.A1(n_347),
.A2(n_15),
.B(n_17),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_489),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_499),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_535),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_357),
.A2(n_64),
.B(n_62),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_414),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_529),
.B(n_18),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_459),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_351),
.B(n_67),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_351),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_438),
.B(n_18),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_351),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_478),
.B(n_19),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_328),
.B(n_19),
.Y(n_599)
);

CKINVDCx6p67_ASAP7_75t_R g600 ( 
.A(n_345),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_391),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_485),
.B(n_20),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_494),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_391),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_497),
.B(n_21),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_391),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_391),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_410),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_443),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_411),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_411),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_363),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_365),
.A2(n_544),
.B(n_372),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_405),
.B(n_22),
.Y(n_614)
);

BUFx8_ASAP7_75t_SL g615 ( 
.A(n_329),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_368),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_527),
.B(n_22),
.Y(n_617)
);

OAI22x1_ASAP7_75t_SL g618 ( 
.A1(n_362),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_411),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_375),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_458),
.B(n_26),
.Y(n_621)
);

AOI22x1_ASAP7_75t_SL g622 ( 
.A1(n_403),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_330),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_411),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_427),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_R g626 ( 
.A1(n_432),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_367),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_331),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_442),
.Y(n_629)
);

OA21x2_ASAP7_75t_L g630 ( 
.A1(n_376),
.A2(n_31),
.B(n_32),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_383),
.Y(n_631)
);

AOI22x1_ASAP7_75t_SL g632 ( 
.A1(n_446),
.A2(n_462),
.B1(n_496),
.B2(n_493),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_445),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_385),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_427),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_507),
.B(n_33),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_393),
.B(n_35),
.Y(n_637)
);

BUFx12f_ASAP7_75t_L g638 ( 
.A(n_503),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_394),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_536),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_395),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_521),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_427),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_427),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_437),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_437),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_400),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_525),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_401),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_467),
.B(n_39),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_332),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_474),
.B(n_41),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_SL g653 ( 
.A1(n_340),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_507),
.B(n_43),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_437),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_404),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_437),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_333),
.B(n_45),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_355),
.B(n_47),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_396),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_396),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_396),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_386),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_335),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_408),
.B(n_47),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_439),
.Y(n_666)
);

INVx5_ASAP7_75t_L g667 ( 
.A(n_439),
.Y(n_667)
);

AOI22x1_ASAP7_75t_SL g668 ( 
.A1(n_342),
.A2(n_364),
.B1(n_384),
.B2(n_356),
.Y(n_668)
);

OA21x2_ASAP7_75t_L g669 ( 
.A1(n_409),
.A2(n_48),
.B(n_49),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_500),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_469),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_469),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_413),
.A2(n_193),
.B(n_323),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_470),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_417),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_337),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_412),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_460),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_469),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_343),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_419),
.B(n_48),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_420),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_463),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_421),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_424),
.Y(n_685)
);

BUFx8_ASAP7_75t_SL g686 ( 
.A(n_498),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_429),
.B(n_50),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_430),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_346),
.Y(n_689)
);

NAND2x1p5_ASAP7_75t_L g690 ( 
.A(n_495),
.B(n_70),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_444),
.Y(n_691)
);

BUFx8_ASAP7_75t_SL g692 ( 
.A(n_508),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_546),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_607),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_554),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_640),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_599),
.B(n_523),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_660),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_615),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_660),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_629),
.B(n_373),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_599),
.B(n_652),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_652),
.B(n_506),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_611),
.Y(n_704)
);

INVx8_ASAP7_75t_L g705 ( 
.A(n_670),
.Y(n_705)
);

BUFx6f_ASAP7_75t_SL g706 ( 
.A(n_608),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_660),
.Y(n_707)
);

CKINVDCx14_ASAP7_75t_R g708 ( 
.A(n_600),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_661),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_661),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_661),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_672),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_624),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_625),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_614),
.B(n_422),
.Y(n_715)
);

BUFx6f_ASAP7_75t_SL g716 ( 
.A(n_585),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_635),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_678),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_651),
.B(n_448),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_621),
.B(n_473),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_645),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_549),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_549),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_629),
.B(n_491),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_549),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_553),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_623),
.Y(n_727)
);

AO21x2_ASAP7_75t_L g728 ( 
.A1(n_552),
.A2(n_433),
.B(n_452),
.Y(n_728)
);

BUFx6f_ASAP7_75t_SL g729 ( 
.A(n_593),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_628),
.B(n_664),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_672),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_676),
.B(n_455),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_670),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_553),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_552),
.B(n_534),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_553),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_565),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_565),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_565),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_672),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_568),
.B(n_540),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_570),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_680),
.B(n_461),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_570),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_557),
.Y(n_745)
);

INVx5_ASAP7_75t_L g746 ( 
.A(n_594),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_662),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_603),
.B(n_349),
.Y(n_748)
);

INVx6_ASAP7_75t_L g749 ( 
.A(n_684),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_666),
.Y(n_750)
);

AOI21x1_ASAP7_75t_L g751 ( 
.A1(n_556),
.A2(n_465),
.B(n_464),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_650),
.B(n_510),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_570),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_677),
.B(n_472),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_573),
.B(n_520),
.Y(n_755)
);

BUFx6f_ASAP7_75t_SL g756 ( 
.A(n_571),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_573),
.B(n_532),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_576),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_576),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_576),
.Y(n_760)
);

AOI21x1_ASAP7_75t_L g761 ( 
.A1(n_564),
.A2(n_480),
.B(n_476),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_597),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_L g763 ( 
.A(n_558),
.B(n_352),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_L g764 ( 
.A(n_563),
.B(n_353),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_581),
.B(n_358),
.Y(n_765)
);

BUFx10_ASAP7_75t_L g766 ( 
.A(n_566),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_638),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_679),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_677),
.B(n_490),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_682),
.Y(n_770)
);

INVx5_ASAP7_75t_L g771 ( 
.A(n_594),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_685),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_653),
.B(n_515),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_678),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_689),
.B(n_566),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_663),
.B(n_359),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_691),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_597),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_663),
.B(n_360),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_601),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_559),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_601),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_601),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_604),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_674),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_604),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_604),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_606),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_545),
.B(n_605),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_735),
.B(n_567),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_728),
.B(n_575),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_728),
.B(n_578),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_722),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_741),
.B(n_605),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_789),
.B(n_613),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_789),
.B(n_655),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_722),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_694),
.B(n_655),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_696),
.B(n_617),
.Y(n_799)
);

AO221x1_ASAP7_75t_L g800 ( 
.A1(n_785),
.A2(n_561),
.B1(n_642),
.B2(n_627),
.C(n_653),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_L g801 ( 
.A(n_697),
.B(n_659),
.C(n_658),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_701),
.B(n_667),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_724),
.B(n_667),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_748),
.B(n_667),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_754),
.A2(n_577),
.B(n_654),
.C(n_572),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_744),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_776),
.B(n_674),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_715),
.B(n_636),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_702),
.A2(n_683),
.B1(n_636),
.B2(n_648),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_732),
.B(n_743),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_718),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_766),
.Y(n_812)
);

INVxp33_ASAP7_75t_L g813 ( 
.A(n_754),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_715),
.B(n_545),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_720),
.B(n_690),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_720),
.B(n_690),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_766),
.B(n_596),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_719),
.B(n_572),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_703),
.B(n_594),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_775),
.B(n_671),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_723),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_765),
.B(n_671),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_705),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_725),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_726),
.B(n_671),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_774),
.B(n_596),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_726),
.B(n_671),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_734),
.Y(n_828)
);

NOR3xp33_ASAP7_75t_L g829 ( 
.A(n_702),
.B(n_654),
.C(n_577),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_730),
.B(n_637),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_779),
.B(n_591),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_734),
.B(n_595),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_727),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_727),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_736),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_736),
.Y(n_836)
);

AND2x6_ASAP7_75t_L g837 ( 
.A(n_730),
.B(n_637),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_737),
.Y(n_838)
);

OR2x6_ASAP7_75t_L g839 ( 
.A(n_705),
.B(n_560),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_738),
.B(n_595),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_745),
.B(n_592),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_769),
.A2(n_602),
.B1(n_598),
.B2(n_550),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_738),
.B(n_595),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_703),
.B(n_598),
.Y(n_844)
);

INVxp67_ASAP7_75t_SL g845 ( 
.A(n_744),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_739),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_781),
.B(n_591),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_739),
.B(n_595),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_769),
.B(n_752),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_742),
.B(n_643),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_753),
.B(n_643),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_781),
.B(n_547),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_753),
.B(n_646),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_767),
.B(n_646),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_758),
.B(n_612),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_733),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_770),
.B(n_547),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_694),
.B(n_616),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_752),
.B(n_665),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_704),
.B(n_620),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_704),
.B(n_631),
.Y(n_861)
);

BUFx6f_ASAP7_75t_SL g862 ( 
.A(n_733),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_713),
.B(n_634),
.Y(n_863)
);

BUFx6f_ASAP7_75t_SL g864 ( 
.A(n_773),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_763),
.A2(n_602),
.B1(n_548),
.B2(n_586),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_759),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_760),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_755),
.B(n_665),
.Y(n_868)
);

BUFx4f_ASAP7_75t_SL g869 ( 
.A(n_823),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_SL g870 ( 
.A(n_811),
.B(n_699),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_808),
.B(n_755),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_856),
.B(n_705),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_859),
.A2(n_764),
.B(n_763),
.C(n_551),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_868),
.A2(n_757),
.B1(n_687),
.B2(n_681),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_813),
.B(n_757),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_810),
.B(n_764),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_795),
.A2(n_771),
.B(n_746),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_795),
.A2(n_771),
.B(n_746),
.Y(n_878)
);

AOI21x1_ASAP7_75t_L g879 ( 
.A1(n_791),
.A2(n_761),
.B(n_751),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_831),
.B(n_708),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_830),
.B(n_746),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_818),
.B(n_762),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_L g883 ( 
.A(n_842),
.B(n_771),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_796),
.A2(n_804),
.B(n_792),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_806),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_791),
.A2(n_788),
.B(n_778),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_805),
.A2(n_687),
.B(n_681),
.C(n_641),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_792),
.A2(n_673),
.B(n_590),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_793),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_830),
.B(n_370),
.Y(n_890)
);

INVx6_ASAP7_75t_L g891 ( 
.A(n_847),
.Y(n_891)
);

NOR2xp67_ASAP7_75t_L g892 ( 
.A(n_822),
.B(n_695),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_820),
.A2(n_780),
.B(n_778),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_849),
.A2(n_502),
.B1(n_504),
.B2(n_501),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_797),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_865),
.A2(n_790),
.B(n_829),
.Y(n_896)
);

OAI321xp33_ASAP7_75t_L g897 ( 
.A1(n_809),
.A2(n_633),
.A3(n_648),
.B1(n_683),
.B2(n_627),
.C(n_551),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_801),
.A2(n_555),
.B(n_574),
.C(n_509),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_852),
.Y(n_899)
);

BUFx6f_ASAP7_75t_SL g900 ( 
.A(n_839),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_807),
.B(n_371),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_802),
.A2(n_783),
.B(n_782),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_794),
.B(n_615),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_806),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_837),
.B(n_841),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_803),
.A2(n_783),
.B(n_782),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_833),
.B(n_569),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_815),
.A2(n_786),
.B(n_784),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_819),
.A2(n_844),
.B(n_816),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_826),
.B(n_374),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_837),
.B(n_784),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_814),
.A2(n_786),
.B(n_787),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_837),
.B(n_787),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_857),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_836),
.Y(n_915)
);

OAI21xp33_ASAP7_75t_L g916 ( 
.A1(n_799),
.A2(n_633),
.B(n_555),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_817),
.A2(n_812),
.B1(n_834),
.B2(n_845),
.Y(n_917)
);

OR2x6_ASAP7_75t_L g918 ( 
.A(n_839),
.B(n_773),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_854),
.B(n_708),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_806),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_850),
.A2(n_717),
.B(n_714),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_858),
.A2(n_647),
.B(n_649),
.C(n_639),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_851),
.A2(n_721),
.B(n_717),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_839),
.Y(n_924)
);

AO22x1_ASAP7_75t_L g925 ( 
.A1(n_821),
.A2(n_609),
.B1(n_562),
.B2(n_626),
.Y(n_925)
);

INVx11_ASAP7_75t_L g926 ( 
.A(n_862),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_855),
.B(n_686),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_853),
.A2(n_380),
.B1(n_381),
.B2(n_378),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_798),
.A2(n_721),
.B(n_772),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_866),
.B(n_693),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_798),
.A2(n_777),
.B(n_693),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_832),
.A2(n_700),
.B(n_698),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_824),
.B(n_828),
.Y(n_933)
);

AO21x1_ASAP7_75t_L g934 ( 
.A1(n_835),
.A2(n_533),
.B(n_505),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_840),
.A2(n_709),
.B(n_707),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_838),
.B(n_710),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_846),
.B(n_711),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_800),
.A2(n_548),
.B1(n_586),
.B2(n_550),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_867),
.A2(n_669),
.B(n_630),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_858),
.B(n_686),
.Y(n_940)
);

AOI21xp33_ASAP7_75t_L g941 ( 
.A1(n_860),
.A2(n_773),
.B(n_669),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_860),
.B(n_382),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_861),
.A2(n_675),
.B(n_688),
.C(n_656),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_861),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_863),
.Y(n_945)
);

AO21x1_ASAP7_75t_L g946 ( 
.A1(n_863),
.A2(n_750),
.B(n_747),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_843),
.A2(n_630),
.B(n_594),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_825),
.B(n_562),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_848),
.A2(n_731),
.B(n_712),
.Y(n_949)
);

OAI21x1_ASAP7_75t_SL g950 ( 
.A1(n_946),
.A2(n_827),
.B(n_583),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_L g951 ( 
.A(n_873),
.B(n_387),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_884),
.A2(n_740),
.B(n_768),
.Y(n_952)
);

NOR2x1_ASAP7_75t_L g953 ( 
.A(n_872),
.B(n_518),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_896),
.A2(n_389),
.B(n_388),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_889),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_886),
.A2(n_584),
.B(n_580),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_907),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_879),
.A2(n_588),
.B(n_587),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_904),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_869),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_876),
.A2(n_579),
.B1(n_390),
.B2(n_392),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_914),
.B(n_609),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_895),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_875),
.B(n_692),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_888),
.A2(n_878),
.B(n_877),
.Y(n_965)
);

BUFx5_ASAP7_75t_L g966 ( 
.A(n_944),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_883),
.A2(n_610),
.B(n_606),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_882),
.B(n_945),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_908),
.A2(n_589),
.B(n_582),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_899),
.B(n_582),
.Y(n_970)
);

BUFx2_ASAP7_75t_SL g971 ( 
.A(n_880),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_933),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_887),
.A2(n_492),
.B(n_397),
.C(n_398),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_911),
.A2(n_610),
.B(n_606),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_912),
.A2(n_589),
.B(n_76),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_871),
.B(n_399),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_874),
.B(n_402),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_933),
.Y(n_978)
);

INVx4_ASAP7_75t_L g979 ( 
.A(n_904),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_898),
.A2(n_407),
.B(n_406),
.Y(n_980)
);

AO31x2_ASAP7_75t_L g981 ( 
.A1(n_894),
.A2(n_52),
.A3(n_53),
.B(n_54),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_913),
.A2(n_78),
.B(n_73),
.Y(n_982)
);

OAI21xp33_ASAP7_75t_L g983 ( 
.A1(n_916),
.A2(n_948),
.B(n_940),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_893),
.A2(n_83),
.B(n_79),
.Y(n_984)
);

NOR2x1_ASAP7_75t_SL g985 ( 
.A(n_905),
.B(n_610),
.Y(n_985)
);

OAI22x1_ASAP7_75t_L g986 ( 
.A1(n_924),
.A2(n_560),
.B1(n_864),
.B2(n_618),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_909),
.A2(n_644),
.B(n_619),
.Y(n_987)
);

AOI221x1_ASAP7_75t_L g988 ( 
.A1(n_941),
.A2(n_684),
.B1(n_657),
.B2(n_619),
.C(n_644),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_902),
.A2(n_93),
.B(n_89),
.Y(n_989)
);

AND2x2_ASAP7_75t_SL g990 ( 
.A(n_870),
.B(n_692),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_SL g991 ( 
.A(n_903),
.B(n_416),
.C(n_415),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_891),
.B(n_684),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_892),
.A2(n_512),
.B(n_423),
.C(n_431),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_930),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_881),
.A2(n_939),
.B(n_947),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_906),
.A2(n_101),
.B(n_95),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_915),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_921),
.A2(n_105),
.B(n_102),
.Y(n_998)
);

AOI221xp5_ASAP7_75t_L g999 ( 
.A1(n_897),
.A2(n_864),
.B1(n_756),
.B2(n_729),
.C(n_716),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_923),
.A2(n_110),
.B(n_106),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_938),
.A2(n_441),
.B(n_435),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_901),
.A2(n_449),
.B(n_447),
.Y(n_1002)
);

AOI21x1_ASAP7_75t_L g1003 ( 
.A1(n_936),
.A2(n_657),
.B(n_749),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_917),
.A2(n_890),
.B(n_942),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_920),
.B(n_119),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_929),
.A2(n_121),
.B(n_120),
.Y(n_1006)
);

BUFx8_ASAP7_75t_L g1007 ( 
.A(n_900),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_937),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_891),
.B(n_450),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_910),
.A2(n_541),
.B(n_542),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_931),
.A2(n_537),
.B(n_539),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_904),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_885),
.B(n_454),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_922),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_928),
.A2(n_514),
.B(n_457),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_885),
.B(n_456),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_932),
.A2(n_263),
.B(n_327),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_968),
.B(n_927),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_997),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_995),
.A2(n_949),
.B(n_935),
.Y(n_1020)
);

AO21x2_ASAP7_75t_L g1021 ( 
.A1(n_950),
.A2(n_985),
.B(n_965),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_960),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_959),
.Y(n_1023)
);

INVx5_ASAP7_75t_L g1024 ( 
.A(n_959),
.Y(n_1024)
);

INVx8_ASAP7_75t_L g1025 ( 
.A(n_959),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_958),
.A2(n_934),
.B(n_943),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_1004),
.A2(n_919),
.B(n_872),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_956),
.A2(n_270),
.B(n_321),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_975),
.A2(n_265),
.B(n_320),
.Y(n_1029)
);

AOI21xp33_ASAP7_75t_SL g1030 ( 
.A1(n_964),
.A2(n_925),
.B(n_918),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_966),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_983),
.B(n_668),
.Y(n_1032)
);

NAND2x1p5_ASAP7_75t_L g1033 ( 
.A(n_979),
.B(n_926),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_970),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_979),
.B(n_872),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_966),
.A2(n_900),
.B1(n_918),
.B2(n_522),
.Y(n_1036)
);

CKINVDCx11_ASAP7_75t_R g1037 ( 
.A(n_1007),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_969),
.A2(n_251),
.B(n_319),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_1005),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_952),
.A2(n_244),
.B(n_316),
.Y(n_1040)
);

OA21x2_ASAP7_75t_L g1041 ( 
.A1(n_988),
.A2(n_530),
.B(n_531),
.Y(n_1041)
);

OA21x2_ASAP7_75t_L g1042 ( 
.A1(n_987),
.A2(n_526),
.B(n_528),
.Y(n_1042)
);

INVx6_ASAP7_75t_L g1043 ( 
.A(n_1007),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_951),
.A2(n_543),
.B(n_466),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_998),
.A2(n_232),
.B(n_313),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_997),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_966),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_955),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_962),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_1000),
.A2(n_230),
.B(n_312),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_992),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_1005),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_SL g1053 ( 
.A(n_990),
.Y(n_1053)
);

BUFx8_ASAP7_75t_L g1054 ( 
.A(n_957),
.Y(n_1054)
);

AO21x2_ASAP7_75t_L g1055 ( 
.A1(n_980),
.A2(n_524),
.B(n_519),
.Y(n_1055)
);

OA21x2_ASAP7_75t_L g1056 ( 
.A1(n_984),
.A2(n_996),
.B(n_989),
.Y(n_1056)
);

NAND3xp33_ASAP7_75t_L g1057 ( 
.A(n_977),
.B(n_632),
.C(n_622),
.Y(n_1057)
);

BUFx12f_ASAP7_75t_L g1058 ( 
.A(n_971),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_963),
.Y(n_1059)
);

AO21x2_ASAP7_75t_L g1060 ( 
.A1(n_973),
.A2(n_517),
.B(n_516),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_1012),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_994),
.A2(n_918),
.B(n_513),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_1006),
.A2(n_210),
.B(n_311),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_966),
.B(n_468),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_994),
.B(n_1008),
.Y(n_1065)
);

AO21x2_ASAP7_75t_L g1066 ( 
.A1(n_954),
.A2(n_511),
.B(n_487),
.Y(n_1066)
);

AO31x2_ASAP7_75t_L g1067 ( 
.A1(n_1014),
.A2(n_54),
.A3(n_56),
.B(n_57),
.Y(n_1067)
);

INVx6_ASAP7_75t_L g1068 ( 
.A(n_953),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_972),
.A2(n_756),
.B1(n_486),
.B2(n_484),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1017),
.A2(n_203),
.B(n_122),
.Y(n_1070)
);

CKINVDCx16_ASAP7_75t_R g1071 ( 
.A(n_991),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_982),
.A2(n_204),
.B(n_127),
.Y(n_1072)
);

OA21x2_ASAP7_75t_L g1073 ( 
.A1(n_974),
.A2(n_483),
.B(n_482),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_1003),
.A2(n_201),
.B(n_130),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_967),
.A2(n_205),
.B(n_131),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_961),
.B(n_706),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1001),
.A2(n_475),
.B(n_471),
.Y(n_1077)
);

OA21x2_ASAP7_75t_L g1078 ( 
.A1(n_976),
.A2(n_479),
.B(n_749),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1019),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1049),
.B(n_978),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1046),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_1022),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1065),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_1029),
.A2(n_1016),
.B(n_1013),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_1024),
.Y(n_1085)
);

INVx8_ASAP7_75t_L g1086 ( 
.A(n_1025),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1065),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1038),
.A2(n_1028),
.B(n_1020),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1048),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1031),
.Y(n_1090)
);

INVxp67_ASAP7_75t_SL g1091 ( 
.A(n_1031),
.Y(n_1091)
);

AOI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_1032),
.A2(n_986),
.B1(n_999),
.B2(n_1015),
.C(n_1002),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_1039),
.B(n_1009),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1059),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1047),
.Y(n_1095)
);

INVx8_ASAP7_75t_L g1096 ( 
.A(n_1025),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1047),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1021),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1061),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1077),
.A2(n_1010),
.B1(n_981),
.B2(n_1011),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1021),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1077),
.A2(n_1057),
.B1(n_1062),
.B2(n_1018),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1023),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1018),
.B(n_981),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1039),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1052),
.A2(n_993),
.B1(n_729),
.B2(n_716),
.Y(n_1106)
);

BUFx12f_ASAP7_75t_L g1107 ( 
.A(n_1037),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1034),
.B(n_1051),
.Y(n_1108)
);

NAND2x1p5_ASAP7_75t_L g1109 ( 
.A(n_1024),
.B(n_981),
.Y(n_1109)
);

OR2x6_ASAP7_75t_L g1110 ( 
.A(n_1058),
.B(n_706),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1026),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1057),
.A2(n_56),
.B1(n_135),
.B2(n_136),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1074),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1045),
.A2(n_1050),
.B(n_1063),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1070),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1062),
.B(n_138),
.Y(n_1116)
);

AOI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1027),
.A2(n_310),
.B(n_143),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1071),
.B(n_141),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1072),
.Y(n_1119)
);

AOI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1064),
.A2(n_309),
.B(n_147),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_SL g1121 ( 
.A(n_1043),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1035),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1064),
.A2(n_303),
.B(n_148),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1067),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1030),
.B(n_145),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1067),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1040),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1054),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1054),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1033),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_1053),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1067),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_1043),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1075),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1068),
.B(n_149),
.Y(n_1135)
);

NAND2x1p5_ASAP7_75t_L g1136 ( 
.A(n_1036),
.B(n_155),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1090),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1086),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1092),
.A2(n_1071),
.B1(n_1076),
.B2(n_1055),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1083),
.B(n_1060),
.Y(n_1140)
);

OAI222xp33_ASAP7_75t_L g1141 ( 
.A1(n_1112),
.A2(n_1036),
.B1(n_1069),
.B2(n_1044),
.C1(n_1030),
.C2(n_1066),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1095),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_1086),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1091),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1104),
.B(n_1078),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1095),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1097),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1091),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1087),
.B(n_1060),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1124),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1126),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1081),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1132),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1098),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1102),
.B(n_1041),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1080),
.B(n_1041),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1079),
.B(n_1042),
.Y(n_1157)
);

OR2x2_ASAP7_75t_L g1158 ( 
.A(n_1111),
.B(n_1042),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1111),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1093),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1089),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1094),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1109),
.B(n_1073),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1125),
.B(n_1056),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1082),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_SL g1166 ( 
.A1(n_1136),
.A2(n_164),
.B(n_177),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1098),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1093),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1108),
.B(n_299),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1093),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1101),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1119),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1109),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1099),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1131),
.B(n_183),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1086),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1119),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1116),
.B(n_298),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1117),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1127),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1105),
.B(n_295),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1135),
.B(n_184),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1135),
.B(n_294),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1127),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1115),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1115),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1134),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1113),
.Y(n_1188)
);

AOI222xp33_ASAP7_75t_L g1189 ( 
.A1(n_1118),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.C1(n_196),
.C2(n_199),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1140),
.B(n_1100),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1150),
.Y(n_1191)
);

OAI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_1139),
.A2(n_1100),
.B(n_1106),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1151),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1140),
.B(n_1123),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1160),
.B(n_1122),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1142),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1153),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1153),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1149),
.B(n_1120),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1138),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1149),
.B(n_1134),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1161),
.B(n_1103),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1142),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1144),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1145),
.B(n_1103),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1144),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1146),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1137),
.Y(n_1208)
);

OAI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1166),
.A2(n_1128),
.B1(n_1129),
.B2(n_1133),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1162),
.B(n_1085),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1148),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1148),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1145),
.B(n_1084),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_L g1214 ( 
.A(n_1138),
.B(n_1133),
.Y(n_1214)
);

INVxp67_ASAP7_75t_SL g1215 ( 
.A(n_1137),
.Y(n_1215)
);

NOR2x1_ASAP7_75t_SL g1216 ( 
.A(n_1173),
.B(n_1110),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1162),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1147),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1170),
.B(n_1084),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1170),
.B(n_1088),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1189),
.A2(n_1121),
.B1(n_1107),
.B2(n_1128),
.Y(n_1221)
);

AND2x4_ASAP7_75t_SL g1222 ( 
.A(n_1176),
.B(n_1130),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1170),
.B(n_1168),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1159),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1164),
.B(n_1156),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1152),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_1165),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1159),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1154),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1155),
.B(n_1129),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1167),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1167),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1174),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1180),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1187),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1168),
.B(n_1114),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1236),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1236),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1234),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1225),
.B(n_1184),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1190),
.B(n_1184),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1190),
.B(n_1180),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1191),
.Y(n_1243)
);

BUFx2_ASAP7_75t_SL g1244 ( 
.A(n_1200),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1227),
.B(n_1175),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1233),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1193),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1234),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1230),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1201),
.B(n_1171),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1205),
.B(n_1173),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1230),
.B(n_1163),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1197),
.Y(n_1253)
);

BUFx2_ASAP7_75t_SL g1254 ( 
.A(n_1200),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1194),
.B(n_1157),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1213),
.B(n_1194),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1198),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1199),
.B(n_1172),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1199),
.B(n_1172),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1217),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1229),
.B(n_1177),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1231),
.B(n_1177),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1232),
.B(n_1219),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1235),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1204),
.B(n_1186),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1224),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1210),
.B(n_1178),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1206),
.B(n_1186),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1211),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1212),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1246),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1243),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1243),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1253),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1237),
.B(n_1220),
.Y(n_1275)
);

NOR3xp33_ASAP7_75t_SL g1276 ( 
.A(n_1245),
.B(n_1209),
.C(n_1192),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1247),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1247),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1256),
.B(n_1220),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1267),
.A2(n_1221),
.B(n_1141),
.Y(n_1280)
);

INVxp67_ASAP7_75t_L g1281 ( 
.A(n_1249),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1263),
.B(n_1216),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1252),
.B(n_1228),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1257),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1255),
.B(n_1218),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1257),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1238),
.B(n_1223),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1240),
.B(n_1215),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1240),
.B(n_1223),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1239),
.Y(n_1290)
);

OR2x6_ASAP7_75t_L g1291 ( 
.A(n_1280),
.B(n_1244),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1290),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1276),
.A2(n_1178),
.B1(n_1183),
.B2(n_1182),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1271),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1272),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1273),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1281),
.B(n_1258),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1285),
.B(n_1259),
.Y(n_1298)
);

AOI32xp33_ASAP7_75t_L g1299 ( 
.A1(n_1282),
.A2(n_1183),
.A3(n_1242),
.B1(n_1241),
.B2(n_1251),
.Y(n_1299)
);

AOI322xp5_ASAP7_75t_L g1300 ( 
.A1(n_1275),
.A2(n_1241),
.A3(n_1242),
.B1(n_1270),
.B2(n_1269),
.C1(n_1264),
.C2(n_1259),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1279),
.B(n_1283),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1293),
.A2(n_1254),
.B1(n_1288),
.B2(n_1271),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1295),
.Y(n_1303)
);

AOI21xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1291),
.A2(n_1110),
.B(n_1278),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1291),
.A2(n_1195),
.B1(n_1289),
.B2(n_1287),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1296),
.Y(n_1306)
);

AO32x1_ASAP7_75t_L g1307 ( 
.A1(n_1292),
.A2(n_1260),
.A3(n_1286),
.B1(n_1277),
.B2(n_1284),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1299),
.A2(n_1254),
.B1(n_1260),
.B2(n_1274),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1297),
.A2(n_1202),
.B1(n_1250),
.B2(n_1248),
.Y(n_1309)
);

A2O1A1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1300),
.A2(n_1214),
.B(n_1222),
.C(n_1143),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1310),
.A2(n_1298),
.B1(n_1301),
.B2(n_1294),
.Y(n_1311)
);

AOI211xp5_ASAP7_75t_SL g1312 ( 
.A1(n_1302),
.A2(n_1169),
.B(n_1181),
.C(n_1226),
.Y(n_1312)
);

OAI222xp33_ASAP7_75t_L g1313 ( 
.A1(n_1308),
.A2(n_1110),
.B1(n_1266),
.B2(n_1265),
.C1(n_1268),
.C2(n_1261),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1304),
.A2(n_1268),
.B(n_1262),
.Y(n_1314)
);

NAND2x1_ASAP7_75t_L g1315 ( 
.A(n_1305),
.B(n_1228),
.Y(n_1315)
);

NAND4xp25_ASAP7_75t_L g1316 ( 
.A(n_1309),
.B(n_1143),
.C(n_1207),
.D(n_1203),
.Y(n_1316)
);

AND4x1_ASAP7_75t_L g1317 ( 
.A(n_1312),
.B(n_1306),
.C(n_1303),
.D(n_1307),
.Y(n_1317)
);

NOR4xp25_ASAP7_75t_L g1318 ( 
.A(n_1311),
.B(n_1307),
.C(n_1196),
.D(n_1207),
.Y(n_1318)
);

O2A1O1Ixp5_ASAP7_75t_L g1319 ( 
.A1(n_1315),
.A2(n_1179),
.B(n_1203),
.C(n_1196),
.Y(n_1319)
);

NOR4xp25_ASAP7_75t_SL g1320 ( 
.A(n_1313),
.B(n_1176),
.C(n_1208),
.D(n_1130),
.Y(n_1320)
);

NAND3xp33_ASAP7_75t_L g1321 ( 
.A(n_1317),
.B(n_1316),
.C(n_1314),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1321),
.B(n_1318),
.C(n_1320),
.Y(n_1322)
);

NOR2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1322),
.B(n_1319),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1323),
.A2(n_1096),
.B1(n_1158),
.B2(n_1188),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1324),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1325),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1326),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1327),
.A2(n_1185),
.B1(n_239),
.B2(n_242),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1328),
.B(n_227),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1329),
.A2(n_252),
.B(n_262),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1330),
.B(n_275),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1331),
.A2(n_279),
.B(n_289),
.Y(n_1332)
);


endmodule