module fake_jpeg_3346_n_694 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_694);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_694;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_612;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_SL g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_60),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_58),
.Y(n_63)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_66),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_27),
.B(n_10),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_100),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_72),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_73),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_74),
.Y(n_208)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_76),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_77),
.Y(n_215)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_79),
.Y(n_216)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_81),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_85),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_86),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_88),
.Y(n_176)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g178 ( 
.A(n_89),
.Y(n_178)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_90),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_92),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_93),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_26),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_25),
.B(n_11),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_95),
.B(n_98),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_96),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_25),
.B(n_11),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_27),
.B(n_9),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_20),
.B(n_12),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_102),
.B(n_104),
.Y(n_179)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_20),
.B(n_12),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_40),
.Y(n_112)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

BUFx24_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_39),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_117),
.B(n_127),
.Y(n_190)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_33),
.Y(n_119)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_119),
.Y(n_222)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_39),
.Y(n_120)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_33),
.Y(n_121)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

INVx6_ASAP7_75t_SL g122 ( 
.A(n_23),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_33),
.Y(n_123)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_39),
.Y(n_124)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_21),
.B(n_12),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_126),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_37),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_37),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_45),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_52),
.Y(n_147)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_39),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_37),
.Y(n_130)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_21),
.B(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_131),
.B(n_132),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_38),
.B(n_7),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_102),
.B(n_55),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_141),
.B(n_154),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_104),
.A2(n_40),
.B1(n_37),
.B2(n_44),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_146),
.A2(n_165),
.B1(n_197),
.B2(n_214),
.Y(n_280)
);

BUFx4f_ASAP7_75t_SL g251 ( 
.A(n_147),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_95),
.B(n_52),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_151),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_44),
.B1(n_52),
.B2(n_41),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_153),
.A2(n_174),
.B1(n_188),
.B2(n_191),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_98),
.B(n_74),
.Y(n_154)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_63),
.Y(n_163)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_163),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_114),
.A2(n_44),
.B1(n_49),
.B2(n_46),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_69),
.A2(n_35),
.B1(n_52),
.B2(n_44),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_166),
.A2(n_92),
.B1(n_88),
.B2(n_89),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_118),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_171),
.B(n_213),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_105),
.A2(n_29),
.B1(n_24),
.B2(n_46),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_49),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_183),
.B(n_184),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_41),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_85),
.B(n_43),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_187),
.B(n_217),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_61),
.A2(n_52),
.B1(n_43),
.B2(n_54),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_109),
.A2(n_29),
.B1(n_24),
.B2(n_32),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_196),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_62),
.A2(n_35),
.B1(n_55),
.B2(n_54),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_202),
.Y(n_253)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_L g209 ( 
.A1(n_130),
.A2(n_32),
.B1(n_35),
.B2(n_59),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_220),
.B1(n_224),
.B2(n_23),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_91),
.B(n_59),
.C(n_50),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_210),
.B(n_23),
.C(n_7),
.Y(n_275)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_212),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_64),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_67),
.A2(n_32),
.B1(n_47),
.B2(n_42),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_72),
.B(n_50),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_218),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_73),
.A2(n_86),
.B1(n_101),
.B2(n_97),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_76),
.A2(n_84),
.B1(n_77),
.B2(n_93),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_107),
.B(n_42),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_0),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_113),
.B(n_47),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_228),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_79),
.A2(n_45),
.B1(n_23),
.B2(n_14),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_166),
.B1(n_214),
.B2(n_220),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_230),
.A2(n_247),
.B1(n_211),
.B2(n_176),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_232),
.A2(n_279),
.B1(n_281),
.B2(n_296),
.Y(n_321)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_137),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_234),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_235),
.Y(n_317)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_149),
.Y(n_236)
);

INVx4_ASAP7_75t_SL g370 ( 
.A(n_236),
.Y(n_370)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_150),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_237),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_178),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_239),
.B(n_248),
.Y(n_320)
);

INVx13_ASAP7_75t_L g241 ( 
.A(n_137),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_241),
.Y(n_328)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_242),
.Y(n_347)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_243),
.Y(n_373)
);

XOR2x2_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_45),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_244),
.B(n_292),
.C(n_293),
.Y(n_313)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_245),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_134),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_194),
.Y(n_250)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_250),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_252),
.B(n_258),
.Y(n_322)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_254),
.Y(n_324)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_137),
.Y(n_255)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_255),
.Y(n_331)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_150),
.Y(n_257)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_257),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_136),
.B(n_14),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_179),
.B(n_14),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_259),
.B(n_262),
.Y(n_327)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_260),
.Y(n_344)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_261),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_227),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_151),
.B(n_14),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_263),
.Y(n_336)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_209),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_265),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_267),
.Y(n_364)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_161),
.Y(n_269)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_269),
.Y(n_335)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_145),
.Y(n_270)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_270),
.Y(n_341)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_271),
.Y(n_342)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_149),
.Y(n_272)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_272),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_143),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_274),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_297),
.Y(n_314)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_139),
.Y(n_276)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_167),
.A2(n_23),
.B1(n_7),
.B2(n_15),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_167),
.A2(n_6),
.B1(n_18),
.B2(n_17),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_157),
.Y(n_282)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_282),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_135),
.B(n_5),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_283),
.B(n_294),
.Y(n_348)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_142),
.Y(n_284)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_284),
.Y(n_362)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_219),
.Y(n_285)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_285),
.Y(n_369)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_201),
.Y(n_286)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_286),
.Y(n_372)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_175),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_198),
.Y(n_288)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_144),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_289),
.B(n_295),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_223),
.A2(n_174),
.B1(n_191),
.B2(n_155),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_290),
.A2(n_180),
.B1(n_193),
.B2(n_159),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_140),
.Y(n_291)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_291),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_160),
.B(n_5),
.C(n_17),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_168),
.B(n_6),
.C(n_17),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_170),
.B(n_19),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_158),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_229),
.A2(n_4),
.B1(n_6),
.B2(n_16),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_175),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_221),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_298),
.B(n_302),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_140),
.Y(n_299)
);

INVx8_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_190),
.B(n_4),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_300),
.B(n_301),
.Y(n_365)
);

BUFx12f_ASAP7_75t_L g301 ( 
.A(n_177),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_169),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_176),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_303),
.B(n_304),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_138),
.B(n_4),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_173),
.B(n_16),
.C(n_19),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_138),
.C(n_162),
.Y(n_337)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_133),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_306),
.Y(n_315)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_222),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_307),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_147),
.B(n_19),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g345 ( 
.A(n_308),
.Y(n_345)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_133),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_310),
.Y(n_329)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_181),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_181),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_311),
.B(n_312),
.Y(n_351)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_159),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_316),
.A2(n_360),
.B1(n_279),
.B2(n_291),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_244),
.B(n_211),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_319),
.B(n_293),
.C(n_292),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_323),
.A2(n_338),
.B1(n_339),
.B2(n_358),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_280),
.A2(n_193),
.B1(n_180),
.B2(n_215),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_325),
.A2(n_251),
.B1(n_266),
.B2(n_256),
.Y(n_378)
);

AOI32xp33_ASAP7_75t_L g334 ( 
.A1(n_246),
.A2(n_240),
.A3(n_264),
.B1(n_231),
.B2(n_273),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_319),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_275),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_265),
.A2(n_152),
.B1(n_226),
.B2(n_216),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_233),
.A2(n_152),
.B1(n_226),
.B2(n_216),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_263),
.B(n_229),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_251),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_233),
.A2(n_247),
.B1(n_231),
.B2(n_230),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_232),
.A2(n_215),
.B1(n_172),
.B2(n_189),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_359),
.A2(n_375),
.B1(n_299),
.B2(n_309),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_251),
.A2(n_172),
.B1(n_204),
.B2(n_200),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_300),
.A2(n_198),
.B1(n_162),
.B2(n_206),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_366),
.A2(n_371),
.B(n_267),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_278),
.A2(n_164),
.B(n_204),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_281),
.A2(n_164),
.B1(n_200),
.B2(n_189),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_376),
.B(n_411),
.C(n_404),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_329),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_377),
.B(n_399),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_378),
.A2(n_383),
.B1(n_389),
.B2(n_397),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_379),
.B(n_365),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_380),
.A2(n_375),
.B1(n_328),
.B2(n_344),
.Y(n_429)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_329),
.Y(n_381)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_381),
.Y(n_428)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_382),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_356),
.A2(n_316),
.B1(n_325),
.B2(n_358),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_384),
.B(n_391),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_371),
.A2(n_257),
.B(n_237),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_385),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_356),
.A2(n_307),
.B1(n_260),
.B2(n_277),
.Y(n_387)
);

OAI21xp33_ASAP7_75t_SL g464 ( 
.A1(n_387),
.A2(n_393),
.B(n_364),
.Y(n_464)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_388),
.Y(n_443)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_390),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_249),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_314),
.A2(n_253),
.B1(n_310),
.B2(n_254),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_392),
.A2(n_395),
.B1(n_420),
.B2(n_350),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_394),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_314),
.A2(n_261),
.B1(n_285),
.B2(n_271),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_396),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_314),
.A2(n_156),
.B1(n_296),
.B2(n_206),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_370),
.Y(n_398)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_398),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_348),
.B(n_238),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_400),
.Y(n_461)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_342),
.Y(n_401)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_401),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_313),
.B(n_305),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_402),
.B(n_403),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_320),
.B(n_268),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_404),
.B(n_362),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_353),
.B(n_286),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_405),
.B(n_410),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_406),
.Y(n_451)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_324),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_407),
.B(n_415),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_321),
.A2(n_156),
.B1(n_269),
.B2(n_272),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_408),
.A2(n_409),
.B1(n_413),
.B2(n_414),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_313),
.A2(n_236),
.B1(n_301),
.B2(n_288),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_365),
.B(n_301),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_337),
.B(n_241),
.C(n_234),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_328),
.A2(n_255),
.B(n_1),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_412),
.A2(n_349),
.B(n_357),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_366),
.A2(n_336),
.B1(n_365),
.B2(n_327),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_322),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_332),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_318),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_416),
.B(n_418),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_315),
.B(n_2),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_421),
.Y(n_435)
);

INVx8_ASAP7_75t_L g418 ( 
.A(n_332),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_342),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_422),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_363),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_317),
.B(n_1),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_369),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_423),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_317),
.B(n_2),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_425),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_368),
.B(n_324),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_426),
.B(n_405),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_429),
.A2(n_440),
.B1(n_389),
.B2(n_386),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g431 ( 
.A(n_400),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_431),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_434),
.A2(n_424),
.B1(n_421),
.B2(n_422),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_436),
.B(n_437),
.C(n_439),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_402),
.B(n_362),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_383),
.A2(n_326),
.B1(n_355),
.B2(n_361),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_413),
.A2(n_331),
.B1(n_349),
.B2(n_370),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_445),
.A2(n_466),
.B(n_412),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_377),
.B(n_372),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_449),
.B(n_391),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_381),
.B(n_333),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_453),
.B(n_454),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_388),
.B(n_396),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_455),
.A2(n_464),
.B(n_410),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_425),
.B(n_333),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_460),
.B(n_442),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_417),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_462),
.B(n_467),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_386),
.A2(n_361),
.B1(n_355),
.B2(n_335),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_465),
.A2(n_390),
.B1(n_382),
.B2(n_419),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_397),
.A2(n_331),
.B1(n_335),
.B2(n_374),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_394),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_458),
.Y(n_468)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_458),
.Y(n_469)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_469),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_445),
.Y(n_470)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_470),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_441),
.A2(n_393),
.B(n_385),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_471),
.A2(n_473),
.B(n_474),
.Y(n_538)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_456),
.Y(n_472)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_472),
.Y(n_515)
);

OAI21xp33_ASAP7_75t_SL g474 ( 
.A1(n_426),
.A2(n_384),
.B(n_379),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_437),
.B(n_376),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_475),
.B(n_479),
.C(n_489),
.Y(n_514)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_456),
.Y(n_476)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_476),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_436),
.B(n_409),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_447),
.Y(n_480)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_480),
.Y(n_536)
);

FAx1_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_378),
.CI(n_411),
.CON(n_481),
.SN(n_481)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_481),
.A2(n_463),
.B(n_427),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_449),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_482),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_455),
.A2(n_398),
.B(n_410),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_483),
.A2(n_487),
.B(n_492),
.Y(n_522)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_444),
.Y(n_485)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_485),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_444),
.B(n_428),
.Y(n_486)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_486),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_457),
.Y(n_488)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_488),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_439),
.B(n_392),
.C(n_405),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_490),
.B(n_491),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_455),
.A2(n_398),
.B(n_408),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_457),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_495),
.Y(n_513)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_447),
.Y(n_494)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_494),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_457),
.Y(n_495)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_496),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_453),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_497),
.B(n_407),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_498),
.A2(n_499),
.B1(n_503),
.B2(n_434),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_501),
.A2(n_504),
.B1(n_466),
.B2(n_429),
.Y(n_512)
);

XOR2x2_ASAP7_75t_SL g530 ( 
.A(n_502),
.B(n_460),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_438),
.A2(n_395),
.B1(n_415),
.B2(n_416),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_438),
.A2(n_401),
.B1(n_403),
.B2(n_406),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_459),
.B(n_462),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_505),
.B(n_491),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_427),
.B(n_346),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_430),
.C(n_452),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_508),
.A2(n_509),
.B1(n_528),
.B2(n_499),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_510),
.B(n_523),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_512),
.A2(n_532),
.B1(n_482),
.B2(n_486),
.Y(n_546)
);

XOR2x2_ASAP7_75t_L g516 ( 
.A(n_479),
.B(n_454),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_516),
.B(n_435),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_517),
.B(n_518),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_475),
.B(n_459),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_484),
.B(n_430),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_520),
.B(n_446),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_484),
.B(n_428),
.C(n_443),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_521),
.B(n_531),
.C(n_535),
.Y(n_547)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_468),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_481),
.A2(n_440),
.B1(n_465),
.B2(n_443),
.Y(n_528)
);

AOI21xp33_ASAP7_75t_L g529 ( 
.A1(n_487),
.A2(n_471),
.B(n_505),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_529),
.B(n_473),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_500),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_489),
.B(n_448),
.C(n_442),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_481),
.A2(n_448),
.B1(n_461),
.B2(n_435),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g534 ( 
.A(n_478),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_534),
.B(n_537),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_506),
.B(n_452),
.C(n_467),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_486),
.Y(n_537)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_540),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_474),
.B(n_481),
.C(n_496),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_541),
.B(n_483),
.C(n_469),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_490),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_446),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_545),
.B(n_548),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_546),
.A2(n_561),
.B1(n_563),
.B2(n_564),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_518),
.B(n_502),
.Y(n_548)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_549),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_SL g550 ( 
.A(n_520),
.B(n_500),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_550),
.B(n_562),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_478),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_551),
.B(n_558),
.Y(n_589)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_507),
.Y(n_553)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_553),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_531),
.B(n_477),
.Y(n_554)
);

CKINVDCx14_ASAP7_75t_R g594 ( 
.A(n_554),
.Y(n_594)
);

INVxp33_ASAP7_75t_L g555 ( 
.A(n_524),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_555),
.B(n_575),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_556),
.B(n_578),
.Y(n_579)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_511),
.Y(n_557)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_557),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_543),
.B(n_504),
.Y(n_560)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_560),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_532),
.A2(n_498),
.B1(n_492),
.B2(n_503),
.Y(n_561)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_524),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_514),
.B(n_494),
.C(n_480),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_565),
.B(n_566),
.C(n_577),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_514),
.B(n_472),
.C(n_476),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_528),
.A2(n_470),
.B1(n_493),
.B2(n_495),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_567),
.A2(n_512),
.B1(n_522),
.B2(n_544),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_SL g569 ( 
.A(n_517),
.B(n_541),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_569),
.B(n_572),
.Y(n_583)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_519),
.Y(n_570)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_570),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_539),
.B(n_340),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_571),
.Y(n_599)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_519),
.Y(n_573)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_573),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_543),
.B(n_542),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_516),
.B(n_450),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_576),
.B(n_538),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_535),
.B(n_432),
.C(n_451),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_509),
.B(n_345),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_575),
.A2(n_522),
.B(n_555),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_584),
.B(n_588),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_577),
.Y(n_587)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_587),
.Y(n_606)
);

FAx1_ASAP7_75t_SL g588 ( 
.A(n_558),
.B(n_530),
.CI(n_509),
.CON(n_588),
.SN(n_588)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_561),
.A2(n_546),
.B1(n_560),
.B2(n_508),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_592),
.A2(n_433),
.B1(n_488),
.B2(n_406),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_559),
.B(n_523),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_595),
.B(n_596),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_574),
.A2(n_527),
.B1(n_544),
.B2(n_470),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_597),
.A2(n_567),
.B1(n_552),
.B2(n_576),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_545),
.A2(n_527),
.B1(n_513),
.B2(n_526),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_598),
.B(n_550),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_549),
.A2(n_538),
.B(n_526),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_602),
.A2(n_525),
.B(n_433),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_604),
.B(n_605),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_566),
.B(n_536),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_607),
.A2(n_616),
.B1(n_593),
.B2(n_414),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_589),
.B(n_568),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_608),
.B(n_615),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_599),
.B(n_565),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_610),
.B(n_611),
.Y(n_644)
);

CKINVDCx16_ASAP7_75t_R g611 ( 
.A(n_584),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_587),
.B(n_551),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_612),
.B(n_614),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_605),
.B(n_548),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_589),
.B(n_568),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_600),
.A2(n_569),
.B1(n_515),
.B2(n_533),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_603),
.B(n_547),
.C(n_572),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_617),
.B(n_623),
.C(n_628),
.Y(n_629)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_581),
.B(n_547),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_618),
.B(n_627),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_602),
.A2(n_525),
.B(n_432),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_619),
.B(n_625),
.Y(n_634)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_620),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_621),
.A2(n_590),
.B(n_585),
.Y(n_635)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_586),
.Y(n_622)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_622),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_603),
.B(n_583),
.C(n_581),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_579),
.A2(n_372),
.B(n_346),
.Y(n_626)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_626),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g627 ( 
.A(n_583),
.B(n_604),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_580),
.B(n_423),
.C(n_343),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_617),
.B(n_582),
.C(n_597),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_631),
.B(n_639),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_624),
.A2(n_594),
.B(n_590),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_632),
.B(n_646),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_635),
.A2(n_619),
.B1(n_613),
.B2(n_625),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_606),
.B(n_591),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_618),
.B(n_592),
.C(n_580),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_640),
.B(n_641),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_608),
.B(n_588),
.C(n_595),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_627),
.B(n_588),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_643),
.B(n_640),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_616),
.B(n_601),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_645),
.B(n_647),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_624),
.B(n_418),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_648),
.A2(n_660),
.B(n_663),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_629),
.B(n_615),
.C(n_623),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_651),
.B(n_652),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_629),
.B(n_609),
.C(n_607),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_631),
.B(n_613),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_653),
.B(n_654),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_SL g654 ( 
.A1(n_634),
.A2(n_620),
.B1(n_621),
.B2(n_593),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_656),
.B(n_659),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_636),
.B(n_622),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_657),
.B(n_658),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_644),
.B(n_628),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_641),
.B(n_609),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_642),
.A2(n_374),
.B(n_343),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_638),
.B(n_418),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_661),
.B(n_637),
.Y(n_670)
);

OR2x2_ASAP7_75t_SL g663 ( 
.A(n_635),
.B(n_423),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_649),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_666),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_SL g668 ( 
.A1(n_662),
.A2(n_634),
.B(n_646),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_SL g680 ( 
.A1(n_668),
.A2(n_656),
.B(n_630),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_670),
.B(n_671),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_652),
.B(n_633),
.Y(n_671)
);

INVx11_ASAP7_75t_L g672 ( 
.A(n_663),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_672),
.B(n_654),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_655),
.B(n_633),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_674),
.B(n_651),
.Y(n_679)
);

AO21x1_ASAP7_75t_L g675 ( 
.A1(n_662),
.A2(n_643),
.B(n_630),
.Y(n_675)
);

OAI21xp33_ASAP7_75t_L g683 ( 
.A1(n_675),
.A2(n_330),
.B(n_369),
.Y(n_683)
);

AOI21xp33_ASAP7_75t_L g685 ( 
.A1(n_676),
.A2(n_679),
.B(n_680),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_664),
.B(n_650),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_677),
.B(n_682),
.Y(n_688)
);

XOR2xp5_ASAP7_75t_L g682 ( 
.A(n_667),
.B(n_665),
.Y(n_682)
);

AOI21x1_ASAP7_75t_L g684 ( 
.A1(n_683),
.A2(n_673),
.B(n_669),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_SL g689 ( 
.A1(n_684),
.A2(n_687),
.B(n_672),
.Y(n_689)
);

NOR3xp33_ASAP7_75t_SL g686 ( 
.A(n_678),
.B(n_675),
.C(n_681),
.Y(n_686)
);

AOI321xp33_ASAP7_75t_SL g690 ( 
.A1(n_686),
.A2(n_354),
.A3(n_330),
.B1(n_357),
.B2(n_373),
.C(n_347),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_SL g687 ( 
.A1(n_683),
.A2(n_673),
.B(n_668),
.Y(n_687)
);

MAJx2_ASAP7_75t_L g691 ( 
.A(n_689),
.B(n_690),
.C(n_688),
.Y(n_691)
);

OAI211xp5_ASAP7_75t_L g692 ( 
.A1(n_691),
.A2(n_685),
.B(n_373),
.C(n_347),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_692),
.B(n_364),
.C(n_350),
.Y(n_693)
);

XNOR2xp5_ASAP7_75t_L g694 ( 
.A(n_693),
.B(n_354),
.Y(n_694)
);


endmodule