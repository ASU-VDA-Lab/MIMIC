module real_jpeg_29353_n_18 (n_17, n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx11_ASAP7_75t_L g93 ( 
.A(n_0),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_0),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g162 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_1),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_163),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_1),
.A2(n_60),
.B1(n_61),
.B2(n_163),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_1),
.A2(n_54),
.B1(n_56),
.B2(n_163),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_2),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_2),
.A2(n_60),
.B1(n_61),
.B2(n_100),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_100),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_2),
.A2(n_54),
.B1(n_56),
.B2(n_100),
.Y(n_244)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_5),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_SL g177 ( 
.A1(n_5),
.A2(n_29),
.B(n_33),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_5),
.B(n_31),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_5),
.A2(n_60),
.B(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_5),
.B(n_60),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_5),
.B(n_74),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_5),
.A2(n_90),
.B1(n_93),
.B2(n_256),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_5),
.A2(n_32),
.B(n_273),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_6),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_174),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_174),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_6),
.A2(n_54),
.B1(n_56),
.B2(n_174),
.Y(n_256)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_49),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_8),
.A2(n_49),
.B1(n_60),
.B2(n_61),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_8),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_9),
.A2(n_37),
.B1(n_60),
.B2(n_61),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_9),
.A2(n_37),
.B1(n_54),
.B2(n_56),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_10),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

OAI32xp33_ASAP7_75t_L g232 ( 
.A1(n_11),
.A2(n_56),
.A3(n_60),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_12),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_12),
.A2(n_27),
.B1(n_60),
.B2(n_61),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_12),
.A2(n_27),
.B1(n_54),
.B2(n_56),
.Y(n_125)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_32),
.B(n_68),
.C(n_71),
.Y(n_67)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_15),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_102),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g169 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_102),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_15),
.A2(n_54),
.B1(n_56),
.B2(n_102),
.Y(n_188)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_17),
.A2(n_25),
.B1(n_26),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_17),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_132),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_17),
.A2(n_54),
.B1(n_56),
.B2(n_132),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_17),
.A2(n_60),
.B1(n_61),
.B2(n_132),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_22),
.B(n_43),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_24),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_26),
.A2(n_35),
.B(n_172),
.C(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_31),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_31),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_28),
.A2(n_31),
.B1(n_99),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_28),
.A2(n_31),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_28),
.A2(n_31),
.B1(n_131),
.B2(n_203),
.Y(n_217)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_32),
.B(n_69),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g281 ( 
.A1(n_32),
.A2(n_61),
.A3(n_69),
.B1(n_274),
.B2(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_33),
.B(n_172),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_82),
.B(n_337),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_75),
.C(n_77),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_44),
.A2(n_45),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_64),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_46),
.B(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_48),
.A2(n_79),
.B1(n_81),
.B2(n_101),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_52),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_52),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_52),
.A2(n_64),
.B1(n_141),
.B2(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_58),
.B(n_63),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_53),
.A2(n_58),
.B1(n_63),
.B2(n_111),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_53),
.A2(n_58),
.B1(n_108),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_53),
.A2(n_58),
.B1(n_127),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_53),
.A2(n_58),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_53),
.A2(n_58),
.B1(n_230),
.B2(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_53),
.B(n_172),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_53),
.A2(n_58),
.B1(n_168),
.B2(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_54),
.B(n_57),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_54),
.B(n_261),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_60),
.B(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_64),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_73),
.B2(n_74),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_65),
.A2(n_66),
.B1(n_74),
.B2(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_66),
.A2(n_74),
.B1(n_117),
.B2(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_66),
.A2(n_74),
.B1(n_162),
.B2(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_66),
.A2(n_74),
.B1(n_129),
.B2(n_206),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_71),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_67),
.A2(n_71),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_67),
.A2(n_71),
.B1(n_161),
.B2(n_164),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_67),
.A2(n_71),
.B1(n_164),
.B2(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_67),
.A2(n_71),
.B1(n_186),
.B2(n_272),
.Y(n_271)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_69),
.Y(n_283)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_75),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_81),
.B1(n_98),
.B2(n_101),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_79),
.A2(n_81),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_330),
.B(n_336),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_144),
.A3(n_153),
.B1(n_328),
.B2(n_329),
.C(n_341),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_133),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_85),
.B(n_133),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_114),
.C(n_121),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_86),
.B(n_114),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_103),
.B1(n_104),
.B2(n_113),
.Y(n_86)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_96),
.B2(n_97),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_88),
.A2(n_97),
.B(n_103),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_88),
.A2(n_89),
.B1(n_105),
.B2(n_106),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_94),
.B(n_95),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_94),
.B1(n_95),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_90),
.A2(n_94),
.B1(n_125),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_90),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_90),
.A2(n_94),
.B1(n_250),
.B2(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_90),
.A2(n_94),
.B1(n_244),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_91),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_91),
.A2(n_92),
.B1(n_179),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_91),
.A2(n_180),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g245 ( 
.A(n_92),
.Y(n_245)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_94),
.Y(n_180)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_109),
.A2(n_112),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_109),
.A2(n_112),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_119),
.B(n_120),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_119),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_134),
.CI(n_143),
.CON(n_133),
.SN(n_133)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_134),
.C(n_143),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_121),
.A2(n_122),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.C(n_130),
.Y(n_122)
);

FAx1_ASAP7_75t_L g311 ( 
.A(n_123),
.B(n_128),
.CI(n_130),
.CON(n_311),
.SN(n_311)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_124),
.B(n_126),
.Y(n_213)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_133),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_142),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_136),
.B1(n_148),
.B2(n_151),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_138),
.C(n_141),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_136),
.B(n_151),
.C(n_152),
.Y(n_331)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_145),
.B(n_146),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

AOI321xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_309),
.A3(n_317),
.B1(n_322),
.B2(n_327),
.C(n_342),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_208),
.C(n_220),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_190),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_156),
.B(n_190),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_175),
.C(n_182),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_157),
.B(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_170),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_165),
.B2(n_166),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_166),
.C(n_170),
.Y(n_197)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_169),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_172),
.B(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_173),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_175),
.A2(n_182),
.B1(n_183),
.B2(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_175),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_178),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_181),
.Y(n_196)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_184),
.B(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_187),
.B(n_189),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_188),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_198),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_197),
.C(n_198),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_195),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_204),
.C(n_207),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_209),
.A2(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_210),
.B(n_211),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_213),
.B(n_214),
.C(n_219),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_215),
.B(n_217),
.C(n_218),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_303),
.B(n_308),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_289),
.B(n_302),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_267),
.B(n_288),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_246),
.B(n_266),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_225),
.B(n_235),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_227),
.B1(n_231),
.B2(n_232),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_229),
.Y(n_233)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_242),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_240),
.C(n_242),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_241),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_243),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_253),
.B(n_265),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_248),
.B(n_252),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_258),
.B(n_264),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_255),
.B(n_257),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_268),
.B(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_280),
.B1(n_286),
.B2(n_287),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_275),
.B1(n_278),
.B2(n_279),
.Y(n_270)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_279),
.C(n_287),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_277),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_280),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_284),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_290),
.B(n_291),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_298),
.C(n_300),
.Y(n_304)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_300),
.B2(n_301),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_298),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_314),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_314),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.C(n_313),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_312),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_311),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_318),
.A2(n_323),
.B(n_326),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_320),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);


endmodule