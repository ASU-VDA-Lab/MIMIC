module fake_jpeg_21793_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_18),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_16),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_35),
.B1(n_32),
.B2(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_28),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_64),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_32),
.B(n_18),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_58),
.C(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_18),
.B(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_13),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_16),
.Y(n_62)
);

OAI32xp33_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_29),
.A3(n_18),
.B1(n_17),
.B2(n_25),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_79),
.B1(n_51),
.B2(n_61),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_69),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_39),
.C(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_14),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_46),
.Y(n_76)
);

XNOR2x1_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_45),
.B1(n_43),
.B2(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_65),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_76),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_56),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_64),
.B(n_56),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_55),
.B(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_54),
.A3(n_70),
.B1(n_76),
.B2(n_68),
.C1(n_79),
.C2(n_9),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_101),
.C(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_68),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_61),
.B1(n_63),
.B2(n_45),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_102),
.A2(n_63),
.B1(n_91),
.B2(n_43),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_81),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_110),
.B1(n_113),
.B2(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_107),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_111),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_63),
.B1(n_84),
.B2(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_2),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

NAND2xp67_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_42),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_98),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_114),
.B(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_111),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_123),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_108),
.Y(n_123)
);

AOI31xp33_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_126),
.A3(n_97),
.B(n_12),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_98),
.B1(n_97),
.B2(n_99),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_124),
.A3(n_26),
.B1(n_20),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_27),
.Y(n_129)
);

AOI211xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_26),
.B(n_8),
.C(n_7),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_121),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_25),
.B(n_5),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_133),
.B1(n_129),
.B2(n_128),
.Y(n_134)
);

OAI211xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_135),
.B(n_133),
.C(n_5),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_7),
.Y(n_137)
);


endmodule