module fake_jpeg_24930_n_180 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_31),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g34 ( 
.A(n_20),
.B(n_0),
.CON(n_34),
.SN(n_34)
);

OR2x2_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_44),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_2),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_31),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_29),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_49),
.B(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_24),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_25),
.B1(n_30),
.B2(n_19),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_61),
.B1(n_75),
.B2(n_17),
.Y(n_87)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_59),
.Y(n_90)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_62),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_22),
.B1(n_25),
.B2(n_16),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_25),
.C(n_36),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_3),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_21),
.B(n_27),
.C(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_32),
.B(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_37),
.A2(n_22),
.B1(n_30),
.B2(n_18),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_23),
.B1(n_6),
.B2(n_7),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_7),
.Y(n_99)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_40),
.A2(n_26),
.B1(n_19),
.B2(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_80),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_99),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_21),
.B(n_17),
.C(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_83),
.B(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_27),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_3),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_95),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_4),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_6),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_67),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_51),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_101),
.A2(n_53),
.B1(n_67),
.B2(n_74),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_73),
.B1(n_64),
.B2(n_56),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_73),
.B1(n_64),
.B2(n_59),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_53),
.B1(n_47),
.B2(n_48),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g119 ( 
.A1(n_78),
.A2(n_70),
.B1(n_10),
.B2(n_8),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_101),
.B(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_84),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_88),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_88),
.Y(n_128)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_98),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_137),
.B(n_107),
.Y(n_145)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_135),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_114),
.B1(n_117),
.B2(n_119),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_96),
.B(n_86),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_85),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_81),
.Y(n_159)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_119),
.B(n_102),
.C(n_108),
.D(n_121),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_148),
.C(n_105),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_151),
.B(n_125),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_136),
.B1(n_132),
.B2(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_123),
.B(n_124),
.C(n_134),
.D(n_127),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_111),
.B1(n_107),
.B2(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_95),
.B1(n_122),
.B2(n_104),
.Y(n_151)
);

OAI321xp33_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_81),
.A3(n_129),
.B1(n_85),
.B2(n_82),
.C(n_100),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_161),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_126),
.C(n_129),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_147),
.C(n_144),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_143),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_166),
.C(n_158),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_146),
.B1(n_142),
.B2(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_160),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_171),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_169),
.B(n_131),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_162),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_160),
.B1(n_155),
.B2(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_173),
.A2(n_172),
.B(n_170),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_76),
.B(n_86),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_131),
.Y(n_179)
);


endmodule