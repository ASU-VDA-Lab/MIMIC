module fake_jpeg_9597_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_16),
.Y(n_63)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_54),
.Y(n_71)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_57),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_63),
.B(n_64),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_29),
.B(n_28),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_24),
.B1(n_32),
.B2(n_35),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_46),
.B1(n_38),
.B2(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_37),
.B(n_16),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_69),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_88),
.B1(n_96),
.B2(n_56),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_80),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_35),
.B1(n_32),
.B2(n_16),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_79),
.A2(n_90),
.B(n_99),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_61),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_82),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_42),
.B1(n_36),
.B2(n_46),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_83),
.A2(n_103),
.B1(n_109),
.B2(n_18),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_20),
.B(n_30),
.C(n_33),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_85),
.B(n_102),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_42),
.B1(n_46),
.B2(n_38),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_20),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_43),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_94),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_49),
.A2(n_38),
.B1(n_36),
.B2(n_32),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_35),
.B1(n_32),
.B2(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_106),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_34),
.B(n_33),
.C(n_23),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_51),
.A2(n_31),
.B1(n_19),
.B2(n_25),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_43),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_48),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_52),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_55),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_49),
.A2(n_31),
.B1(n_19),
.B2(n_25),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_115),
.B(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_0),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_123),
.B(n_102),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_26),
.B1(n_31),
.B2(n_25),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_119),
.A2(n_132),
.B1(n_18),
.B2(n_29),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_48),
.B1(n_62),
.B2(n_73),
.Y(n_164)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_133),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_105),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_43),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_55),
.B1(n_67),
.B2(n_37),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_73),
.B1(n_78),
.B2(n_89),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_26),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_87),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_37),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_138),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_74),
.B(n_48),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_126),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_95),
.B1(n_75),
.B2(n_100),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_166),
.B1(n_129),
.B2(n_120),
.Y(n_178)
);

OAI22x1_ASAP7_75t_SL g141 ( 
.A1(n_136),
.A2(n_79),
.B1(n_99),
.B2(n_90),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_152),
.B1(n_164),
.B2(n_115),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_142),
.B(n_161),
.C(n_21),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_75),
.B(n_85),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_165),
.B(n_123),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_144),
.B(n_148),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_146),
.B(n_149),
.Y(n_195)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_156),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_81),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

BUFx4f_ASAP7_75t_SL g153 ( 
.A(n_112),
.Y(n_153)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

AOI31xp33_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_98),
.A3(n_92),
.B(n_77),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_155),
.B(n_163),
.Y(n_175)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_135),
.B(n_98),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_159),
.B(n_160),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_23),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_134),
.B(n_14),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_162),
.B(n_169),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_138),
.B(n_93),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_113),
.A2(n_108),
.B1(n_62),
.B2(n_29),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_168),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_121),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_62),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_173),
.A2(n_197),
.B1(n_166),
.B2(n_164),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_174),
.B(n_198),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_176),
.A2(n_200),
.B(n_4),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_117),
.Y(n_177)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_178),
.A2(n_186),
.B1(n_190),
.B2(n_154),
.Y(n_216)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_189),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_123),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_181),
.B(n_161),
.Y(n_215)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_125),
.A3(n_117),
.B1(n_127),
.B2(n_114),
.Y(n_182)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_127),
.B(n_114),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_143),
.B(n_162),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_128),
.B1(n_133),
.B2(n_78),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_110),
.Y(n_188)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_139),
.A2(n_78),
.B1(n_28),
.B2(n_21),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_131),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_202),
.C(n_21),
.Y(n_220)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_131),
.B1(n_112),
.B2(n_28),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_82),
.Y(n_198)
);

AO22x1_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_97),
.B1(n_2),
.B2(n_3),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_145),
.B(n_82),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_204),
.B(n_3),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_173),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_145),
.B(n_153),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_185),
.B(n_200),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_187),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_216),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_140),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_220),
.C(n_221),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_179),
.B1(n_189),
.B2(n_190),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_219),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_167),
.B1(n_160),
.B2(n_153),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_217),
.A2(n_225),
.B1(n_200),
.B2(n_192),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_181),
.B(n_10),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_176),
.B(n_9),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_151),
.C(n_150),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_223),
.C(n_230),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_1),
.C(n_2),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_203),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_231),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_4),
.C(n_5),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_233),
.B(n_5),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_250),
.B1(n_232),
.B2(n_205),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_179),
.C(n_180),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_249),
.C(n_220),
.Y(n_259)
);

AND2x6_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_182),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_252),
.B(n_209),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_202),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_185),
.B1(n_175),
.B2(n_199),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_251),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_217),
.B1(n_216),
.B2(n_208),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_177),
.B1(n_199),
.B2(n_193),
.Y(n_273)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_274),
.B1(n_251),
.B2(n_236),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_235),
.A2(n_214),
.B1(n_225),
.B2(n_231),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_257),
.A2(n_269),
.B1(n_6),
.B2(n_7),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_267),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_234),
.B(n_245),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_273),
.B1(n_247),
.B2(n_250),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_254),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_270),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_206),
.C(n_219),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_265),
.C(n_267),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_221),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_177),
.C(n_227),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_239),
.A2(n_212),
.B1(n_230),
.B2(n_201),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_201),
.B(n_184),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_223),
.B1(n_193),
.B2(n_184),
.Y(n_272)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_272),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_276),
.B(n_277),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_260),
.Y(n_278)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_283),
.C(n_271),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_269),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_233),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_259),
.C(n_245),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_287),
.C(n_288),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_270),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_289),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_241),
.C(n_249),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_261),
.C(n_262),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_258),
.A2(n_248),
.B1(n_242),
.B2(n_8),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_257),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_291),
.B1(n_268),
.B2(n_275),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_265),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_296),
.C(n_300),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_287),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_301),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_299),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_268),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_278),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_285),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_295),
.A2(n_280),
.B1(n_291),
.B2(n_283),
.Y(n_310)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_284),
.B(n_13),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_314),
.C(n_313),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_12),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_313),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_14),
.Y(n_314)
);

XOR2x2_ASAP7_75t_SL g316 ( 
.A(n_310),
.B(n_304),
.Y(n_316)
);

AOI21x1_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_308),
.B(n_311),
.Y(n_322)
);

OA21x2_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_304),
.B(n_292),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_317),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_302),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_307),
.C(n_306),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_319),
.C(n_315),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_323),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_324),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_325),
.B(n_321),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_326),
.C(n_316),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_318),
.Y(n_331)
);


endmodule