module real_jpeg_30117_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_343, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_343;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_0),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_0),
.A2(n_34),
.B1(n_36),
.B2(n_157),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_0),
.A2(n_100),
.B1(n_101),
.B2(n_157),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_0),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_303)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_2),
.A2(n_34),
.B1(n_36),
.B2(n_63),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_2),
.A2(n_63),
.B1(n_100),
.B2(n_101),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_2),
.A2(n_63),
.B1(n_160),
.B2(n_161),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_3),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_3),
.A2(n_34),
.B1(n_36),
.B2(n_221),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_3),
.A2(n_100),
.B1(n_101),
.B2(n_221),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_3),
.A2(n_160),
.B1(n_161),
.B2(n_221),
.Y(n_332)
);

BUFx12_ASAP7_75t_L g136 ( 
.A(n_4),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_5),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_5),
.A2(n_34),
.B1(n_36),
.B2(n_140),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_5),
.A2(n_100),
.B1(n_101),
.B2(n_140),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_5),
.A2(n_140),
.B1(n_160),
.B2(n_161),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_6),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_6),
.A2(n_34),
.B1(n_36),
.B2(n_117),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_6),
.A2(n_100),
.B1(n_101),
.B2(n_117),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_6),
.A2(n_117),
.B1(n_160),
.B2(n_161),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_8),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_8),
.A2(n_34),
.B1(n_36),
.B2(n_202),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_8),
.A2(n_100),
.B1(n_101),
.B2(n_202),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_8),
.A2(n_160),
.B1(n_161),
.B2(n_202),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_9),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_10),
.B(n_36),
.Y(n_35)
);

A2O1A1O1Ixp25_ASAP7_75t_L g38 ( 
.A1(n_10),
.A2(n_35),
.B(n_36),
.C(n_39),
.D(n_43),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_10),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_60),
.B(n_64),
.Y(n_87)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_10),
.A2(n_100),
.B(n_102),
.C(n_103),
.D(n_107),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_10),
.B(n_100),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_10),
.B(n_134),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_10),
.A2(n_136),
.B(n_159),
.C(n_160),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_10),
.A2(n_82),
.B1(n_160),
.B2(n_161),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_11),
.A2(n_34),
.B1(n_36),
.B2(n_45),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_45),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_11),
.A2(n_45),
.B1(n_100),
.B2(n_101),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_11),
.A2(n_45),
.B1(n_160),
.B2(n_161),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_12),
.A2(n_34),
.B1(n_36),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_12),
.A2(n_56),
.B1(n_100),
.B2(n_101),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_12),
.A2(n_56),
.B1(n_160),
.B2(n_161),
.Y(n_194)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_31),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_13),
.A2(n_36),
.B(n_40),
.C(n_42),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g101 ( 
.A(n_14),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_15),
.A2(n_34),
.B1(n_36),
.B2(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_335),
.B(n_338),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_330),
.B(n_334),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_317),
.B(n_329),
.Y(n_19)
);

OAI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_281),
.A3(n_310),
.B1(n_315),
.B2(n_316),
.C(n_342),
.Y(n_20)
);

AOI321xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_231),
.A3(n_270),
.B1(n_275),
.B2(n_280),
.C(n_343),
.Y(n_21)
);

NOR3xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_181),
.C(n_227),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_148),
.B(n_180),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_123),
.B(n_147),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_95),
.B(n_122),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_69),
.B(n_94),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_47),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_28),
.B(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_38),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_29),
.B(n_38),
.Y(n_78)
);

AOI32xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.A3(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_30),
.B(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_31),
.B(n_61),
.Y(n_60)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_34),
.B(n_120),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_41),
.Y(n_40)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_36),
.A2(n_101),
.A3(n_102),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_39),
.A2(n_42),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_39),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_39),
.A2(n_42),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_39),
.A2(n_42),
.B1(n_247),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_43),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_55),
.B(n_57),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_46),
.A2(n_57),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_46),
.A2(n_144),
.B1(n_179),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_46),
.A2(n_144),
.B1(n_204),
.B2(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_46),
.A2(n_144),
.B(n_256),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_59),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_54),
.C(n_59),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_51),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_51),
.A2(n_103),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_51),
.A2(n_103),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_51),
.A2(n_103),
.B1(n_259),
.B2(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_51),
.A2(n_103),
.B(n_322),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_52),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.Y(n_104)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_55),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_64),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_60),
.A2(n_68),
.B1(n_116),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_60),
.A2(n_68),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_60),
.A2(n_201),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_60),
.A2(n_77),
.B(n_220),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_67),
.A2(n_85),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_67),
.A2(n_74),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx5_ASAP7_75t_SL g219 ( 
.A(n_67),
.Y(n_219)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_79),
.B(n_93),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_78),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_78),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_77),
.B(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_86),
.B(n_92),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_90),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_82),
.A2(n_100),
.B(n_135),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_97),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_113),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_110),
.C(n_113),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_101),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_109),
.A2(n_129),
.B(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_109),
.A2(n_189),
.B1(n_216),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_109),
.A2(n_189),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_112),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_118),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_125),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_141),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_142),
.C(n_143),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_132),
.C(n_138),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_128),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_134),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_134),
.A2(n_166),
.B1(n_194),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_134),
.A2(n_166),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_134),
.A2(n_166),
.B1(n_325),
.B2(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_134),
.A2(n_166),
.B(n_332),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_136),
.B1(n_160),
.B2(n_161),
.Y(n_167)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_139),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_150),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_164),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_152),
.B(n_153),
.C(n_164),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_158),
.B1(n_162),
.B2(n_163),
.Y(n_153)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_156),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_158),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_162),
.Y(n_185)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_172),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_174),
.C(n_177),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_168),
.B(n_169),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_166),
.B(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_166),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_170),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_178),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_182),
.A2(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_206),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_183),
.B(n_206),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_198),
.C(n_205),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_187),
.C(n_197),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_197),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B(n_191),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_192),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_195),
.B(n_196),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_195),
.A2(n_196),
.B(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_195),
.A2(n_238),
.B1(n_266),
.B2(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_195),
.A2(n_238),
.B1(n_293),
.B2(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_205),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_203),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_217),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_208),
.B(n_217),
.C(n_226),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_212),
.C(n_214),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_222),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_228),
.B(n_229),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_251),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_251),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_243),
.C(n_250),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_243),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_242),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_234),
.Y(n_242)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_240),
.C(n_242),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_241),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_249),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_249),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_249),
.A2(n_264),
.B(n_267),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_269),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_261),
.B1(n_262),
.B2(n_268),
.Y(n_252)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_257),
.B(n_260),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_257),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_260),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_260),
.A2(n_283),
.B1(n_284),
.B2(n_295),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_261),
.B(n_268),
.C(n_269),
.Y(n_311)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_271),
.A2(n_276),
.B(n_279),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_272),
.B(n_273),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_298),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_282),
.B(n_298),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_295),
.C(n_296),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_292),
.B2(n_294),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_287),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_291),
.C(n_292),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_288),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_289),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_291),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_302),
.C(n_306),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_292),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_294),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_301),
.C(n_309),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_297),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_309),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_303),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_308),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_319),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_328),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_323),
.B1(n_326),
.B2(n_327),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_321),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_323),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_327),
.C(n_328),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_333),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_331),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_337),
.B(n_340),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);


endmodule