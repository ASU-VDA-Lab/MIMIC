module fake_jpeg_6673_n_104 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_20),
.B(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_35),
.Y(n_45)
);

NOR3xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.C(n_1),
.Y(n_33)
);

AO22x1_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_13),
.B1(n_15),
.B2(n_22),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_1),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_39),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_26),
.C(n_24),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_26),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_21),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_51),
.Y(n_64)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_32),
.B1(n_30),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_32),
.B1(n_60),
.B2(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_60),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_30),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_16),
.B(n_23),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_44),
.B(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_17),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_67),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_32),
.B1(n_43),
.B2(n_28),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_37),
.B1(n_28),
.B2(n_32),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_51),
.B1(n_54),
.B2(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_70),
.Y(n_82)
);

MAJx2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_41),
.C(n_39),
.Y(n_68)
);

XOR2x2_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_53),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_41),
.B(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_56),
.B(n_57),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_76),
.B(n_68),
.Y(n_87)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_65),
.B1(n_43),
.B2(n_71),
.Y(n_84)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_27),
.B(n_25),
.C(n_22),
.D(n_35),
.Y(n_88)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_87),
.A2(n_80),
.B(n_82),
.Y(n_89)
);

OAI322xp33_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_77),
.A3(n_27),
.B1(n_25),
.B2(n_35),
.C1(n_31),
.C2(n_7),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_27),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_81),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_91),
.B(n_93),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_87),
.A2(n_82),
.B(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_91),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_3),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_9),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_100),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_8),
.Y(n_104)
);


endmodule