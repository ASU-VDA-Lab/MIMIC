module fake_jpeg_24594_n_161 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_161);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_29),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_15),
.B1(n_25),
.B2(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_32),
.B1(n_25),
.B2(n_16),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_20),
.Y(n_37)
);

AOI21xp33_ASAP7_75t_SL g32 ( 
.A1(n_15),
.A2(n_1),
.B(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_48),
.B1(n_14),
.B2(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_35),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_31),
.B1(n_30),
.B2(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_31),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

AO22x1_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_62),
.B(n_65),
.C(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_13),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_64),
.B1(n_49),
.B2(n_43),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_34),
.B1(n_35),
.B2(n_20),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_40),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_43),
.C(n_41),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_78),
.C(n_59),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_49),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_39),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_45),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_77),
.B1(n_64),
.B2(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_39),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_47),
.C(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_17),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_40),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_36),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_68),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_96),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_56),
.B1(n_58),
.B2(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_95),
.B1(n_98),
.B2(n_19),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_78),
.B(n_67),
.Y(n_110)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_72),
.C(n_66),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_13),
.B1(n_17),
.B2(n_26),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_68),
.A2(n_14),
.B1(n_23),
.B2(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_79),
.Y(n_99)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_85),
.B(n_91),
.C(n_90),
.D(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_94),
.B(n_73),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_96),
.C(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_67),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_76),
.B(n_79),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_106),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_121),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_103),
.B1(n_113),
.B2(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_105),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_99),
.B1(n_97),
.B2(n_80),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_36),
.B(n_104),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_100),
.C(n_106),
.Y(n_126)
);

NAND4xp25_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_116),
.C(n_22),
.D(n_20),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_132),
.B(n_133),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_107),
.C(n_101),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_117),
.C(n_122),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_116),
.B(n_110),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_104),
.B(n_2),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_22),
.Y(n_143)
);

AOI322xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_29),
.A3(n_51),
.B1(n_22),
.B2(n_20),
.C1(n_5),
.C2(n_6),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_115),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_120),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_137),
.C(n_140),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_118),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_139),
.B(n_143),
.Y(n_146)
);

OAI21x1_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_114),
.B(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_51),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_1),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_134),
.B(n_51),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

AOI21x1_ASAP7_75t_L g150 ( 
.A1(n_146),
.A2(n_136),
.B(n_140),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_152),
.B1(n_149),
.B2(n_9),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_22),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_3),
.C(n_6),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_157),
.B(n_8),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_149),
.Y(n_157)
);

AOI221xp5_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_160),
.B1(n_156),
.B2(n_8),
.C(n_22),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_158),
.A2(n_8),
.B(n_11),
.Y(n_160)
);


endmodule