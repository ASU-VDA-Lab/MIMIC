module fake_ariane_1181_n_111 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_38, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_111);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_111;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_106;
wire n_53;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_84;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_82;
wire n_57;
wire n_70;
wire n_85;
wire n_94;
wire n_101;
wire n_58;
wire n_65;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_87;
wire n_81;
wire n_55;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_59;
wire n_63;
wire n_99;
wire n_54;

OAI21x1_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_20),
.B(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_8),
.B(n_13),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_43),
.B1(n_42),
.B2(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_7),
.B(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx8_ASAP7_75t_SL g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_39),
.A2(n_24),
.B1(n_34),
.B2(n_4),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_0),
.B(n_37),
.Y(n_67)
);

OAI21x1_ASAP7_75t_L g68 ( 
.A1(n_2),
.A2(n_30),
.B(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_15),
.B(n_21),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_16),
.Y(n_72)
);

NOR2xp67_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_6),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_9),
.Y(n_78)
);

NOR2xp67_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_10),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_53),
.B(n_11),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_12),
.C(n_25),
.Y(n_81)
);

OR2x6_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_68),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_52),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_54),
.B1(n_66),
.B2(n_63),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_69),
.Y(n_86)
);

OAI22x1_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_53),
.B1(n_70),
.B2(n_60),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_52),
.B(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

OAI21x1_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_55),
.B(n_57),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_95),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_84),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_96),
.B1(n_99),
.B2(n_84),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_87),
.B1(n_72),
.B2(n_91),
.Y(n_104)
);

NAND4xp25_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_81),
.C(n_91),
.D(n_58),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_106),
.Y(n_107)
);

AOI222xp33_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_104),
.B1(n_65),
.B2(n_35),
.C1(n_38),
.C2(n_41),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_65),
.B1(n_29),
.B2(n_45),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_108),
.B(n_46),
.Y(n_110)
);

AO21x2_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_26),
.B(n_47),
.Y(n_111)
);


endmodule