module fake_jpeg_736_n_55 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_55);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_15;

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_19),
.B(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_23),
.Y(n_25)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_33),
.B(n_20),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_28),
.B1(n_22),
.B2(n_15),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_25),
.C(n_20),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_2),
.C(n_3),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_15),
.B1(n_28),
.B2(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_0),
.Y(n_40)
);

OA21x2_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_28),
.B(n_4),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_13),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_49),
.C(n_50),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_47),
.C(n_10),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_11),
.B(n_9),
.Y(n_53)
);

BUFx24_ASAP7_75t_SL g54 ( 
.A(n_53),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_51),
.Y(n_55)
);


endmodule