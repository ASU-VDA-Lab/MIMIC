module real_jpeg_5253_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_70;
wire n_74;
wire n_41;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_225;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx8_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_1),
.B(n_65),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_2),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_2),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_2),
.B(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_3),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_3),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_4),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_4),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_4),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_4),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_4),
.B(n_139),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_5),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_5),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_5),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_5),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_5),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_32),
.Y(n_47)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_8),
.Y(n_110)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_8),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_8),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_12),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_12),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_12),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_12),
.B(n_168),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_12),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_13),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_13),
.B(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_13),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_13),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_13),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_13),
.B(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_14),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_15),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_15),
.B(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_152),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_150),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_130),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_19),
.B(n_130),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_70),
.B2(n_129),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_45),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.C(n_41),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_23),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_24),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_135)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_29),
.Y(n_180)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_35),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_36),
.B(n_41),
.Y(n_149)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_53),
.B1(n_68),
.B2(n_69),
.Y(n_45)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B(n_52),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_48),
.Y(n_52)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_63),
.Y(n_174)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_111),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_84),
.C(n_101),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_132),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g232 ( 
.A(n_72),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_77),
.CI(n_81),
.CON(n_72),
.SN(n_72)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_77),
.C(n_81),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_76),
.Y(n_206)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_80),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_84),
.A2(n_85),
.B1(n_101),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.C(n_96),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_86),
.A2(n_87),
.B1(n_96),
.B2(n_97),
.Y(n_225)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_91),
.B(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_126),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.C(n_148),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_131),
.B(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_134),
.B(n_148),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.C(n_141),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_135),
.B(n_136),
.Y(n_218)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_141),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_142),
.B(n_146),
.Y(n_197)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21x1_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_227),
.B(n_231),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_212),
.B(n_226),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_194),
.B(n_211),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_183),
.B(n_193),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_164),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_161),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_175),
.B2(n_176),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_169),
.C(n_175),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_181),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_188),
.B(n_192),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_210),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_210),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_198),
.C(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_207),
.C(n_209),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_215),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_222),
.C(n_223),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_229),
.Y(n_231)
);


endmodule