module fake_jpeg_27138_n_288 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_11),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_26),
.B(n_27),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_24),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_19),
.B1(n_15),
.B2(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_12),
.B1(n_13),
.B2(n_21),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_34),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_27),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_52),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_25),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_26),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_43),
.B1(n_45),
.B2(n_41),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_33),
.B1(n_45),
.B2(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_68),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_32),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_33),
.B1(n_45),
.B2(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_71),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_10),
.C(n_11),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_46),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_49),
.Y(n_89)
);

AO22x2_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_37),
.B1(n_29),
.B2(n_42),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_57),
.B(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_34),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_83),
.B(n_85),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_51),
.C(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_78),
.B(n_46),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_62),
.C(n_52),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_97),
.B1(n_53),
.B2(n_67),
.Y(n_113)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_57),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_57),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_80),
.B1(n_79),
.B2(n_59),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_110),
.B1(n_111),
.B2(n_122),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_118),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_80),
.A3(n_77),
.B1(n_32),
.B2(n_42),
.Y(n_105)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_87),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_107),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_80),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_86),
.B(n_99),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_77),
.B1(n_55),
.B2(n_42),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_77),
.B1(n_82),
.B2(n_67),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_74),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_43),
.B1(n_58),
.B2(n_63),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_145),
.B(n_103),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_91),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_125),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_76),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_111),
.B1(n_104),
.B2(n_106),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_127),
.B1(n_133),
.B2(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_135),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_109),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_76),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_99),
.B1(n_101),
.B2(n_92),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_99),
.B1(n_120),
.B2(n_114),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_87),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_85),
.Y(n_144)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

AO21x1_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_109),
.B(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_167),
.B1(n_132),
.B2(n_136),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_138),
.Y(n_182)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_84),
.C(n_117),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_165),
.C(n_168),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_83),
.C(n_28),
.Y(n_156)
);

XNOR2x1_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_135),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_169),
.B1(n_170),
.B2(n_137),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_20),
.B(n_24),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_163),
.B(n_126),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_74),
.B(n_20),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_74),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_136),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_131),
.C(n_148),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_128),
.A2(n_61),
.B1(n_43),
.B2(n_63),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_35),
.C(n_61),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_43),
.B1(n_18),
.B2(n_24),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_23),
.B1(n_20),
.B2(n_18),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_179),
.A2(n_191),
.B1(n_196),
.B2(n_198),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_180),
.A2(n_189),
.B(n_160),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_153),
.C(n_165),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_184),
.C(n_164),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_194),
.B1(n_172),
.B2(n_65),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_154),
.C(n_152),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

NOR2x1_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_22),
.Y(n_187)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_134),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_56),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_162),
.B(n_10),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_190),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_16),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_162),
.B(n_174),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_193),
.A2(n_195),
.B(n_160),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_23),
.B1(n_22),
.B2(n_16),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_166),
.B(n_65),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_28),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_166),
.Y(n_197)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_197),
.B(n_163),
.C(n_159),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_28),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_178),
.C(n_189),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_184),
.A2(n_157),
.B(n_168),
.C(n_158),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_203),
.B1(n_206),
.B2(n_202),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_191),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_171),
.C(n_154),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_216),
.C(n_218),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_152),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_213),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_150),
.B1(n_171),
.B2(n_167),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_187),
.B1(n_196),
.B2(n_198),
.Y(n_226)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_35),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_56),
.C(n_35),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_176),
.C(n_189),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_213),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_212),
.B(n_180),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_220),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_233),
.C(n_221),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_218),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_204),
.B(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_226),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_R g227 ( 
.A(n_203),
.B(n_25),
.Y(n_227)
);

XOR2x2_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_25),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_207),
.B(n_22),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_228),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_56),
.B1(n_29),
.B2(n_2),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_230),
.B1(n_217),
.B2(n_200),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_215),
.A2(n_0),
.B(n_1),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_234),
.B(n_200),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_214),
.B(n_202),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_234),
.B(n_221),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_245),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_200),
.B1(n_209),
.B2(n_199),
.Y(n_243)
);

AO221x1_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_222),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_252)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_247),
.C(n_0),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_233),
.Y(n_249)
);

OAI321xp33_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_201),
.A3(n_16),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_247)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_230),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_251),
.B(n_253),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_3),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_1),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_1),
.B(n_2),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_257),
.C(n_258),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_235),
.A2(n_237),
.B(n_245),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_29),
.C(n_4),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_236),
.A2(n_244),
.B(n_4),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_5),
.C(n_6),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_269),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_29),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_268),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_29),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_29),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_264),
.B(n_250),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_271),
.Y(n_278)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_254),
.B(n_6),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_5),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_272),
.A2(n_266),
.B(n_261),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_260),
.B(n_5),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_267),
.C(n_268),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_279),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_273),
.C(n_276),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_275),
.C(n_7),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_280),
.B1(n_7),
.B2(n_8),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_6),
.C(n_7),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_9),
.C(n_261),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_9),
.Y(n_288)
);


endmodule