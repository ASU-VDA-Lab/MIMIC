module fake_ibex_1601_n_3214 (n_151, n_85, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_13, n_122, n_523, n_116, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_355, n_474, n_594, n_407, n_102, n_490, n_568, n_52, n_448, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_536, n_352, n_290, n_558, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_267, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3214);

input n_151;
input n_85;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_523;
input n_116;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_594;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_536;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_267;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3214;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2498;
wire n_1802;
wire n_2235;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3168;
wire n_884;
wire n_667;
wire n_2396;
wire n_3135;
wire n_850;
wire n_3175;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_3192;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_641;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_2995;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2846;
wire n_2685;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_605;
wire n_2373;
wire n_630;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_702;
wire n_971;
wire n_1326;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_2987;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3203;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_3117;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3091;
wire n_3006;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3055;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_3003;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_607;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2991;
wire n_2234;
wire n_847;
wire n_2699;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_615;
wire n_2905;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1539;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2352;
wire n_2212;
wire n_2263;
wire n_2716;
wire n_863;
wire n_597;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3167;
wire n_997;
wire n_2308;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2654;
wire n_2463;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_2997;
wire n_1349;
wire n_634;
wire n_991;
wire n_1223;
wire n_1331;
wire n_961;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_2862;
wire n_3100;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_604;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_636;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_3196;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_768;
wire n_839;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_2818;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3011;
wire n_1167;
wire n_818;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_1256;
wire n_2798;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3109;
wire n_1961;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_688;
wire n_3104;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_682;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1572;
wire n_1635;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_750;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_3207;
wire n_1379;
wire n_759;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_635;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_783;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3114;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2302;
wire n_3056;
wire n_2560;
wire n_2092;
wire n_3008;
wire n_1365;
wire n_1472;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_658;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_866;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_3195;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_450),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_557),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_190),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_115),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_301),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_408),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_591),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_5),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_503),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_144),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_44),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_184),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_51),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_224),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_538),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_388),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_499),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_548),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_192),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_447),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_229),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_262),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_157),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_70),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_322),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_546),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_459),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_94),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_53),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_26),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_466),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_205),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_89),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_1),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_4),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_23),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_527),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_585),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_391),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_282),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_146),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_296),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_5),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_280),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_409),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_0),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_370),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_504),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_19),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_583),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_218),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_65),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_442),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_95),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_368),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_101),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_567),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_376),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_264),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_227),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_108),
.Y(n_656)
);

CKINVDCx16_ASAP7_75t_R g657 ( 
.A(n_563),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_50),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_542),
.Y(n_659)
);

BUFx8_ASAP7_75t_SL g660 ( 
.A(n_0),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_56),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_201),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_124),
.Y(n_663)
);

CKINVDCx16_ASAP7_75t_R g664 ( 
.A(n_571),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_316),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_203),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_212),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_352),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_483),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_208),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_398),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_437),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_449),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_457),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_595),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_199),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_556),
.Y(n_677)
);

CKINVDCx16_ASAP7_75t_R g678 ( 
.A(n_164),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_510),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_258),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_412),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_246),
.Y(n_682)
);

BUFx8_ASAP7_75t_SL g683 ( 
.A(n_377),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_426),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_520),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_492),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_569),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_34),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_243),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_586),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_433),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_257),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_399),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_258),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_415),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_536),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_262),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_13),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_416),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_196),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_373),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_48),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_189),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_335),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_424),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_511),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_447),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_554),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_581),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_408),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_487),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_22),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_204),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_486),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_488),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_192),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_412),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_66),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_326),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_331),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_328),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_240),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_274),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_221),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_168),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_366),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_241),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_593),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_383),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_105),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_172),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_239),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_263),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_579),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_467),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_383),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_468),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_489),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_144),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_530),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_20),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_526),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_300),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_516),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_592),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_403),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_52),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_303),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_288),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_267),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_101),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_522),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_79),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_519),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_401),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_573),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_118),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_306),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_93),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_238),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_127),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_456),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_517),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_541),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_212),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_521),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_177),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_446),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_480),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_211),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_253),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_344),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_201),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_417),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_472),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_178),
.Y(n_776)
);

CKINVDCx16_ASAP7_75t_R g777 ( 
.A(n_16),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_51),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_52),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_587),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_391),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_500),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_195),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_37),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_555),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_244),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_167),
.Y(n_787)
);

CKINVDCx16_ASAP7_75t_R g788 ( 
.A(n_307),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_2),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_58),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_315),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_440),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_252),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_491),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_537),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_313),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_279),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_264),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_121),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_171),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_354),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_496),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_484),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_359),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_243),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_493),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_375),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_180),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_256),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_68),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_70),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_473),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_116),
.Y(n_813)
);

BUFx10_ASAP7_75t_L g814 ( 
.A(n_217),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_455),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_221),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_174),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_523),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_399),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_353),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_277),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_335),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_387),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_147),
.Y(n_824)
);

BUFx10_ASAP7_75t_L g825 ( 
.A(n_290),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_338),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_416),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_508),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_60),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_149),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_103),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_92),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_228),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_589),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_439),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_549),
.Y(n_836)
);

CKINVDCx16_ASAP7_75t_R g837 ( 
.A(n_453),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_3),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_435),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_240),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_293),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_208),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_565),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_68),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_424),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_89),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_222),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_574),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_285),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_66),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_136),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_124),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_422),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_422),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_134),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_248),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_272),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_381),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_421),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_236),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_48),
.Y(n_861)
);

BUFx10_ASAP7_75t_L g862 ( 
.A(n_359),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_340),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_478),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_207),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_346),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_228),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_281),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_580),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_207),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_518),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_375),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_173),
.Y(n_873)
);

BUFx5_ASAP7_75t_L g874 ( 
.A(n_156),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_578),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_388),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_514),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_213),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_83),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_308),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_309),
.Y(n_881)
);

HB1xp67_ASAP7_75t_SL g882 ( 
.A(n_385),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_139),
.Y(n_883)
);

BUFx10_ASAP7_75t_L g884 ( 
.A(n_122),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_296),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_566),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_395),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_104),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_588),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_332),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_30),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_474),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_338),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_111),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_560),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_17),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_524),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_131),
.Y(n_898)
);

CKINVDCx16_ASAP7_75t_R g899 ( 
.A(n_423),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_35),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_576),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_509),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_122),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_350),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_277),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_63),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_33),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_36),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_352),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_543),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_384),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_233),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_59),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_71),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_194),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_476),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_155),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_218),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_403),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_63),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_263),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_10),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_582),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_18),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_433),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_561),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_363),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_287),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_443),
.Y(n_929)
);

BUFx2_ASAP7_75t_R g930 ( 
.A(n_427),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_272),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_200),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_12),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_547),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_545),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_515),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_395),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_446),
.Y(n_938)
);

CKINVDCx14_ASAP7_75t_R g939 ( 
.A(n_223),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_287),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_360),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_465),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_326),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_490),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_105),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_257),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_195),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_436),
.Y(n_948)
);

CKINVDCx16_ASAP7_75t_R g949 ( 
.A(n_414),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_384),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_145),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_77),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_215),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_160),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_41),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_295),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_161),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_308),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_143),
.Y(n_959)
);

BUFx5_ASAP7_75t_L g960 ( 
.A(n_67),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_288),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_145),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_143),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_828),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_751),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_927),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_722),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_751),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_633),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_652),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_874),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_634),
.Y(n_972)
);

CKINVDCx16_ASAP7_75t_R g973 ( 
.A(n_678),
.Y(n_973)
);

NOR2xp67_ASAP7_75t_L g974 ( 
.A(n_820),
.B(n_2),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_777),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_831),
.B(n_3),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_814),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_788),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_814),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_715),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_764),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_766),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_802),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_709),
.B(n_4),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_939),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_837),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_899),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_657),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_634),
.Y(n_989)
);

INVxp67_ASAP7_75t_SL g990 ( 
.A(n_710),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_728),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_710),
.Y(n_992)
);

INVxp33_ASAP7_75t_SL g993 ( 
.A(n_596),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_814),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_713),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_709),
.B(n_6),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_596),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_738),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_886),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_664),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_660),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_949),
.B(n_6),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_713),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_683),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_733),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_910),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_825),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_610),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_711),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_610),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_598),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_612),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_599),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_606),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_639),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_613),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_599),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_733),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_605),
.B(n_7),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_826),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_613),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_825),
.B(n_7),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_604),
.B(n_8),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_621),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_644),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_826),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_621),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_940),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_676),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_600),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_940),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_608),
.Y(n_1032)
);

INVxp67_ASAP7_75t_SL g1033 ( 
.A(n_608),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_611),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_692),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_611),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_626),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_825),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_731),
.Y(n_1039)
);

CKINVDCx16_ASAP7_75t_R g1040 ( 
.A(n_882),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_626),
.Y(n_1041)
);

INVxp33_ASAP7_75t_SL g1042 ( 
.A(n_600),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_731),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_743),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_693),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_643),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_743),
.Y(n_1047)
);

INVxp67_ASAP7_75t_SL g1048 ( 
.A(n_746),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_746),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_601),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_761),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_695),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_698),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_601),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_R g1055 ( 
.A(n_679),
.B(n_469),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_761),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_774),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_603),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_774),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_603),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_699),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_614),
.B(n_8),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_614),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_643),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_783),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_783),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_645),
.Y(n_1067)
);

INVxp67_ASAP7_75t_SL g1068 ( 
.A(n_838),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_838),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_879),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_862),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_645),
.Y(n_1072)
);

INVxp67_ASAP7_75t_SL g1073 ( 
.A(n_879),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_707),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_771),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_669),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_894),
.Y(n_1077)
);

NOR2xp67_ASAP7_75t_L g1078 ( 
.A(n_894),
.B(n_9),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_669),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_922),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_840),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_922),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_866),
.Y(n_1083)
);

INVxp33_ASAP7_75t_SL g1084 ( 
.A(n_615),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_956),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_874),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_877),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_956),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_659),
.B(n_9),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_877),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_878),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_880),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_874),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_874),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_889),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_889),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_677),
.B(n_10),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_874),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_1006),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_1006),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_964),
.B(n_615),
.Y(n_1101)
);

AND3x2_ASAP7_75t_L g1102 ( 
.A(n_966),
.B(n_930),
.C(n_809),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_968),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_989),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_971),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_995),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1003),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1005),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_971),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1086),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_972),
.B(n_616),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1018),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_1009),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1026),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1033),
.B(n_607),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1028),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_990),
.B(n_616),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1048),
.B(n_1068),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1031),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1093),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_1094),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1073),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_969),
.B(n_602),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_992),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_967),
.B(n_962),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1020),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_970),
.B(n_622),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1098),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1009),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1009),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1009),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_981),
.B(n_602),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1032),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_996),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1034),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_1036),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1039),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1043),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_997),
.B(n_862),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_1013),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1044),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1047),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1049),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1051),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1056),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1057),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_1059),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1017),
.B(n_862),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1065),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1066),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1069),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_984),
.A2(n_864),
.B(n_690),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_982),
.B(n_618),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_983),
.B(n_864),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1070),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_1030),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_993),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_1077),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1022),
.B(n_627),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1080),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1050),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1082),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1085),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1088),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1019),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1060),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1058),
.B(n_884),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_973),
.B(n_957),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_1054),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1023),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1078),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_976),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_974),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1089),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1097),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_977),
.B(n_696),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1062),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_993),
.B(n_618),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_979),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_994),
.B(n_708),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1007),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1038),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1042),
.B(n_619),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1096),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1071),
.B(n_714),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_1011),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_1060),
.Y(n_1187)
);

OA21x2_ASAP7_75t_L g1188 ( 
.A1(n_1063),
.A2(n_744),
.B(n_742),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1008),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1055),
.B(n_754),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1002),
.B(n_629),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1042),
.B(n_619),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1095),
.Y(n_1193)
);

CKINVDCx16_ASAP7_75t_R g1194 ( 
.A(n_1040),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1010),
.Y(n_1195)
);

AND3x2_ASAP7_75t_L g1196 ( 
.A(n_1084),
.B(n_638),
.C(n_630),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1084),
.A2(n_623),
.B1(n_624),
.B2(n_620),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1012),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1016),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1063),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1021),
.Y(n_1201)
);

NAND2x1_ASAP7_75t_L g1202 ( 
.A(n_985),
.B(n_769),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1024),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_985),
.B(n_884),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1027),
.B(n_623),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1037),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1041),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1046),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1064),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1067),
.B(n_624),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1072),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_988),
.B(n_884),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1076),
.B(n_625),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1079),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_988),
.B(n_898),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1087),
.Y(n_1216)
);

INVx5_ASAP7_75t_L g1217 ( 
.A(n_1090),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1000),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_980),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_975),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_975),
.B(n_775),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1001),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_978),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_978),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_986),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_986),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_991),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_998),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_999),
.B(n_625),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1004),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_987),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_987),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1014),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1014),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1015),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1015),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1092),
.Y(n_1237)
);

INVx4_ASAP7_75t_L g1238 ( 
.A(n_1025),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1025),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1029),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1029),
.A2(n_785),
.B(n_780),
.Y(n_1241)
);

AND2x6_ASAP7_75t_L g1242 ( 
.A(n_1035),
.B(n_910),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1035),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1045),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1045),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1052),
.B(n_834),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1052),
.B(n_628),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1053),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1053),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1061),
.B(n_843),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1061),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1074),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1074),
.B(n_935),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1075),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1075),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1081),
.B(n_898),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1081),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1083),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1083),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1091),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1091),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1092),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_965),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_965),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1006),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1011),
.A2(n_932),
.B1(n_631),
.B2(n_635),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1009),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_971),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_965),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_964),
.B(n_628),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_965),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_964),
.B(n_631),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_966),
.B(n_898),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_965),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_971),
.Y(n_1275)
);

AND2x6_ASAP7_75t_L g1276 ( 
.A(n_1022),
.B(n_942),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_965),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_969),
.B(n_892),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_966),
.B(n_874),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_965),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1006),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_997),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1009),
.Y(n_1283)
);

NAND2xp33_ASAP7_75t_L g1284 ( 
.A(n_985),
.B(n_874),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_966),
.B(n_874),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_971),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_965),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_971),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_965),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_964),
.B(n_635),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_966),
.B(n_960),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_993),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_965),
.B(n_641),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1006),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1060),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_966),
.B(n_960),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_964),
.B(n_636),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_964),
.B(n_636),
.Y(n_1298)
);

NAND2xp33_ASAP7_75t_L g1299 ( 
.A(n_985),
.B(n_960),
.Y(n_1299)
);

INVxp33_ASAP7_75t_L g1300 ( 
.A(n_997),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_966),
.B(n_960),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_965),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_965),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_964),
.B(n_637),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_965),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_997),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_965),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_971),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_993),
.Y(n_1309)
);

NAND2xp33_ASAP7_75t_L g1310 ( 
.A(n_985),
.B(n_960),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1169),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1172),
.A2(n_640),
.B1(n_642),
.B2(n_637),
.Y(n_1312)
);

INVx8_ASAP7_75t_L g1313 ( 
.A(n_1276),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1103),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1134),
.B(n_711),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1294),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1294),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1177),
.A2(n_960),
.B1(n_653),
.B2(n_658),
.Y(n_1318)
);

OR2x6_ASAP7_75t_L g1319 ( 
.A(n_1219),
.B(n_647),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1294),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1100),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1136),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1263),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1136),
.Y(n_1324)
);

INVx5_ASAP7_75t_L g1325 ( 
.A(n_1136),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1264),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1186),
.Y(n_1327)
);

AND2x6_ASAP7_75t_L g1328 ( 
.A(n_1198),
.B(n_711),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1179),
.B(n_895),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1100),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1269),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1157),
.B(n_646),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1179),
.B(n_895),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1271),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_SL g1335 ( 
.A(n_1292),
.B(n_640),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1125),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1170),
.A2(n_960),
.B1(n_661),
.B2(n_665),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1118),
.B(n_960),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1274),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1136),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1124),
.B(n_1126),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1181),
.B(n_897),
.Y(n_1342)
);

NAND3xp33_ASAP7_75t_L g1343 ( 
.A(n_1197),
.B(n_646),
.C(n_642),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_1186),
.Y(n_1344)
);

AND2x2_ASAP7_75t_SL g1345 ( 
.A(n_1188),
.B(n_650),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1161),
.Y(n_1346)
);

INVxp67_ASAP7_75t_SL g1347 ( 
.A(n_1118),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1247),
.B(n_648),
.Y(n_1348)
);

INVx6_ASAP7_75t_L g1349 ( 
.A(n_1144),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1277),
.Y(n_1350)
);

BUFx4f_ASAP7_75t_L g1351 ( 
.A(n_1189),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1280),
.Y(n_1352)
);

INVx5_ASAP7_75t_L g1353 ( 
.A(n_1144),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1118),
.B(n_897),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1181),
.B(n_901),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1182),
.B(n_901),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1207),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1287),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1265),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1265),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1144),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1182),
.B(n_902),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1147),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1289),
.Y(n_1364)
);

NAND2xp33_ASAP7_75t_L g1365 ( 
.A(n_1276),
.B(n_902),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1161),
.B(n_648),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1121),
.B(n_711),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1302),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1122),
.B(n_916),
.Y(n_1369)
);

INVx5_ASAP7_75t_L g1370 ( 
.A(n_1147),
.Y(n_1370)
);

INVxp33_ASAP7_75t_L g1371 ( 
.A(n_1282),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1170),
.A2(n_667),
.B1(n_668),
.B2(n_662),
.Y(n_1372)
);

BUFx8_ASAP7_75t_SL g1373 ( 
.A(n_1262),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1198),
.B(n_916),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1147),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1149),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1207),
.B(n_672),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1174),
.B(n_923),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1300),
.B(n_651),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1303),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1174),
.B(n_923),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1305),
.Y(n_1382)
);

INVx5_ASAP7_75t_L g1383 ( 
.A(n_1149),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_1282),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1300),
.B(n_651),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1307),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1099),
.Y(n_1387)
);

AO22x2_ASAP7_75t_L g1388 ( 
.A1(n_1173),
.A2(n_674),
.B1(n_680),
.B2(n_673),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1166),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1188),
.A2(n_694),
.B1(n_717),
.B2(n_681),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1137),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1137),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1158),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1188),
.A2(n_726),
.B1(n_730),
.B2(n_720),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1158),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1293),
.B(n_926),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1306),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1121),
.B(n_711),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1162),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1162),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1165),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1111),
.B(n_926),
.Y(n_1402)
);

NAND2xp33_ASAP7_75t_R g1403 ( 
.A(n_1309),
.B(n_649),
.Y(n_1403)
);

OR2x6_ASAP7_75t_L g1404 ( 
.A(n_1219),
.B(n_732),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1162),
.Y(n_1405)
);

BUFx10_ASAP7_75t_L g1406 ( 
.A(n_1309),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1138),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1145),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1117),
.B(n_1293),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1306),
.B(n_649),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1152),
.A2(n_757),
.B1(n_760),
.B2(n_755),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1150),
.Y(n_1412)
);

BUFx4f_ASAP7_75t_L g1413 ( 
.A(n_1189),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1155),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1201),
.B(n_765),
.Y(n_1415)
);

INVx5_ASAP7_75t_L g1416 ( 
.A(n_1158),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1250),
.A2(n_656),
.B1(n_663),
.B2(n_655),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1201),
.B(n_1203),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1168),
.B(n_655),
.Y(n_1419)
);

INVxp33_ASAP7_75t_L g1420 ( 
.A(n_1266),
.Y(n_1420)
);

INVx1_ASAP7_75t_SL g1421 ( 
.A(n_1200),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1293),
.B(n_934),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1133),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1175),
.B(n_934),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1099),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1133),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1160),
.Y(n_1427)
);

INVxp33_ASAP7_75t_L g1428 ( 
.A(n_1256),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1152),
.B(n_936),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1164),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1203),
.B(n_936),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1135),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1135),
.Y(n_1433)
);

INVx5_ASAP7_75t_L g1434 ( 
.A(n_1276),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1152),
.B(n_944),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1115),
.B(n_944),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1165),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1099),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1141),
.Y(n_1439)
);

CKINVDCx16_ASAP7_75t_R g1440 ( 
.A(n_1194),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1141),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1281),
.Y(n_1442)
);

INVxp33_ASAP7_75t_L g1443 ( 
.A(n_1273),
.Y(n_1443)
);

BUFx10_ASAP7_75t_L g1444 ( 
.A(n_1278),
.Y(n_1444)
);

INVx4_ASAP7_75t_L g1445 ( 
.A(n_1189),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1142),
.Y(n_1446)
);

AND2x6_ASAP7_75t_L g1447 ( 
.A(n_1208),
.B(n_650),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1115),
.B(n_685),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1165),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1278),
.B(n_663),
.C(n_656),
.Y(n_1450)
);

INVx5_ASAP7_75t_L g1451 ( 
.A(n_1276),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1142),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1295),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1143),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1115),
.B(n_686),
.Y(n_1455)
);

XNOR2xp5_ASAP7_75t_L g1456 ( 
.A(n_1262),
.B(n_957),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1143),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1281),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1175),
.B(n_597),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1146),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1165),
.B(n_687),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1146),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_SL g1463 ( 
.A(n_1187),
.B(n_666),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1151),
.Y(n_1464)
);

BUFx4f_ASAP7_75t_L g1465 ( 
.A(n_1195),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1175),
.B(n_1180),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1163),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1175),
.B(n_706),
.Y(n_1468)
);

AND2x2_ASAP7_75t_SL g1469 ( 
.A(n_1241),
.B(n_650),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1104),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1106),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1101),
.B(n_734),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1270),
.B(n_735),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1272),
.B(n_1290),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1195),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1107),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1140),
.B(n_890),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1108),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1112),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1114),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1250),
.A2(n_876),
.B1(n_885),
.B2(n_666),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1121),
.B(n_737),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1156),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1191),
.A2(n_885),
.B1(n_887),
.B2(n_876),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1195),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1191),
.B(n_900),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1116),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1139),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1119),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1159),
.Y(n_1490)
);

BUFx10_ASAP7_75t_L g1491 ( 
.A(n_1196),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1195),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1241),
.A2(n_773),
.B1(n_778),
.B2(n_768),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1191),
.B(n_1148),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1222),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1159),
.Y(n_1496)
);

NAND2xp33_ASAP7_75t_L g1497 ( 
.A(n_1276),
.B(n_740),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1127),
.A2(n_791),
.B1(n_792),
.B2(n_789),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1113),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1120),
.B(n_1105),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1159),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1127),
.A2(n_800),
.B1(n_801),
.B2(n_793),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1120),
.B(n_745),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1105),
.B(n_1109),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1297),
.B(n_1298),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1304),
.B(n_752),
.Y(n_1506)
);

AND2x6_ASAP7_75t_L g1507 ( 
.A(n_1208),
.B(n_650),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1127),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1279),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1123),
.A2(n_807),
.B1(n_808),
.B2(n_804),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1113),
.Y(n_1511)
);

AND2x6_ASAP7_75t_L g1512 ( 
.A(n_1209),
.B(n_650),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1285),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1167),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1178),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1222),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1209),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1291),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1296),
.B(n_756),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1211),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1183),
.Y(n_1521)
);

NOR3xp33_ASAP7_75t_L g1522 ( 
.A(n_1253),
.B(n_617),
.C(n_609),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1259),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1301),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1192),
.B(n_887),
.Y(n_1525)
);

NAND2x1p5_ASAP7_75t_L g1526 ( 
.A(n_1217),
.B(n_819),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1110),
.B(n_763),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1211),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1171),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1204),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1214),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1217),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1123),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1216),
.Y(n_1534)
);

OR2x6_ASAP7_75t_L g1535 ( 
.A(n_1238),
.B(n_822),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1217),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1259),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1240),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1212),
.B(n_900),
.Y(n_1539)
);

AOI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1128),
.A2(n_841),
.B(n_833),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1113),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1180),
.B(n_632),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1132),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1132),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1216),
.B(n_782),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1113),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1153),
.A2(n_890),
.B1(n_896),
.B2(n_888),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1154),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1154),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1215),
.Y(n_1550)
);

INVx4_ASAP7_75t_L g1551 ( 
.A(n_1217),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1205),
.B(n_1210),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1268),
.Y(n_1553)
);

INVx5_ASAP7_75t_L g1554 ( 
.A(n_1267),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1241),
.A2(n_850),
.B1(n_855),
.B2(n_849),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1176),
.B(n_675),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1176),
.Y(n_1557)
);

INVx4_ASAP7_75t_L g1558 ( 
.A(n_1242),
.Y(n_1558)
);

BUFx10_ASAP7_75t_L g1559 ( 
.A(n_1242),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1213),
.B(n_928),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1185),
.B(n_794),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1185),
.B(n_795),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1284),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1275),
.Y(n_1564)
);

INVx4_ASAP7_75t_L g1565 ( 
.A(n_1242),
.Y(n_1565)
);

AO22x2_ASAP7_75t_L g1566 ( 
.A1(n_1253),
.A2(n_860),
.B1(n_861),
.B2(n_858),
.Y(n_1566)
);

INVxp33_ASAP7_75t_L g1567 ( 
.A(n_1240),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1286),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1286),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1238),
.B(n_863),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1184),
.B(n_803),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1193),
.B(n_806),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1202),
.Y(n_1573)
);

INVx5_ASAP7_75t_L g1574 ( 
.A(n_1267),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1288),
.B(n_818),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1288),
.B(n_836),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1308),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1347),
.B(n_1199),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1347),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1409),
.B(n_1206),
.Y(n_1580)
);

NAND2x1p5_ASAP7_75t_L g1581 ( 
.A(n_1434),
.B(n_1222),
.Y(n_1581)
);

BUFx8_ASAP7_75t_L g1582 ( 
.A(n_1389),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1371),
.B(n_1229),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1311),
.Y(n_1584)
);

INVxp67_ASAP7_75t_SL g1585 ( 
.A(n_1346),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1423),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1443),
.B(n_1218),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1437),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1469),
.A2(n_1242),
.B1(n_1310),
.B2(n_1299),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1437),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1557),
.B(n_1221),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1490),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1496),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1384),
.B(n_1227),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1453),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1474),
.B(n_1221),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1357),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1384),
.B(n_1228),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1483),
.B(n_1220),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1505),
.B(n_1310),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1313),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1501),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1421),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1409),
.B(n_1190),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1373),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_SL g1606 ( 
.A(n_1313),
.B(n_1406),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1403),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1346),
.A2(n_1246),
.B1(n_1224),
.B2(n_1225),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1533),
.B(n_1543),
.Y(n_1609)
);

NOR3xp33_ASAP7_75t_L g1610 ( 
.A(n_1440),
.B(n_1237),
.C(n_1243),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1397),
.B(n_1246),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1397),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1319),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1423),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1319),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1313),
.Y(n_1616)
);

BUFx5_ASAP7_75t_L g1617 ( 
.A(n_1447),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1366),
.B(n_1235),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1544),
.B(n_888),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1463),
.B(n_1230),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1321),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1335),
.Y(n_1622)
);

AO221x1_ASAP7_75t_L g1623 ( 
.A1(n_1493),
.A2(n_1244),
.B1(n_1245),
.B2(n_1239),
.C(n_1234),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1321),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1314),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1521),
.B(n_1223),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1522),
.B(n_1224),
.C(n_1223),
.Y(n_1627)
);

OR2x6_ASAP7_75t_L g1628 ( 
.A(n_1535),
.B(n_1570),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1323),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1326),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1332),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1321),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1522),
.B(n_1231),
.C(n_1226),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1331),
.Y(n_1634)
);

INVx8_ASAP7_75t_L g1635 ( 
.A(n_1535),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1387),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1429),
.A2(n_1130),
.B(n_1129),
.Y(n_1637)
);

AO22x2_ASAP7_75t_L g1638 ( 
.A1(n_1493),
.A2(n_1243),
.B1(n_1258),
.B2(n_1235),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1426),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_SL g1640 ( 
.A(n_1406),
.B(n_1102),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1354),
.B(n_896),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1466),
.A2(n_891),
.B(n_903),
.C(n_881),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1411),
.A2(n_907),
.B1(n_912),
.B2(n_906),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1354),
.B(n_904),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1319),
.Y(n_1645)
);

AO221x1_ASAP7_75t_L g1646 ( 
.A1(n_1555),
.A2(n_1244),
.B1(n_1245),
.B2(n_1239),
.C(n_1234),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1548),
.B(n_904),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1334),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1494),
.A2(n_1231),
.B1(n_1232),
.B2(n_1226),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1404),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1379),
.B(n_1232),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1385),
.B(n_1234),
.Y(n_1652)
);

NOR3xp33_ASAP7_75t_L g1653 ( 
.A(n_1343),
.B(n_1258),
.C(n_1243),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1339),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1336),
.A2(n_909),
.B1(n_911),
.B2(n_905),
.Y(n_1655)
);

OR2x6_ASAP7_75t_L g1656 ( 
.A(n_1535),
.B(n_1234),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1403),
.Y(n_1657)
);

INVx4_ASAP7_75t_L g1658 ( 
.A(n_1434),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1387),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1426),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1549),
.B(n_905),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1439),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1439),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1550),
.B(n_1233),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1327),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1486),
.B(n_1239),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_R g1667 ( 
.A(n_1344),
.B(n_1258),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1404),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1350),
.B(n_913),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1446),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1352),
.B(n_1358),
.Y(n_1671)
);

AND2x6_ASAP7_75t_SL g1672 ( 
.A(n_1570),
.B(n_1236),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1508),
.B(n_1239),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1364),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1530),
.B(n_1248),
.Y(n_1675)
);

INVx4_ASAP7_75t_L g1676 ( 
.A(n_1434),
.Y(n_1676)
);

INVx2_ASAP7_75t_SL g1677 ( 
.A(n_1404),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1451),
.B(n_848),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1436),
.B(n_913),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1477),
.B(n_1244),
.Y(n_1680)
);

INVxp67_ASAP7_75t_SL g1681 ( 
.A(n_1365),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1515),
.B(n_1249),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1368),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1436),
.B(n_917),
.Y(n_1684)
);

BUFx5_ASAP7_75t_L g1685 ( 
.A(n_1447),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1539),
.A2(n_918),
.B1(n_920),
.B2(n_917),
.Y(n_1686)
);

NOR2x1p5_ASAP7_75t_L g1687 ( 
.A(n_1410),
.B(n_1244),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1380),
.B(n_920),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1446),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1454),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1451),
.B(n_871),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1454),
.Y(n_1692)
);

OR2x6_ASAP7_75t_L g1693 ( 
.A(n_1570),
.B(n_1245),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1484),
.B(n_1245),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1451),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1312),
.B(n_1251),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1378),
.B(n_921),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1498),
.A2(n_1260),
.B1(n_1261),
.B2(n_1257),
.C(n_1254),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1457),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1560),
.B(n_1251),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1378),
.B(n_928),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1396),
.B(n_875),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1469),
.A2(n_915),
.B1(n_919),
.B2(n_914),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1457),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1419),
.B(n_1251),
.Y(n_1705)
);

AOI22x1_ASAP7_75t_L g1706 ( 
.A1(n_1563),
.A2(n_1130),
.B1(n_1131),
.B2(n_1129),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1382),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1488),
.A2(n_933),
.B1(n_938),
.B2(n_929),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1386),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1418),
.B(n_1252),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1514),
.B(n_1252),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1525),
.B(n_1428),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1418),
.B(n_1252),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1547),
.B(n_1252),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1325),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1471),
.B(n_961),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1422),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1470),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1478),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1476),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1567),
.B(n_1255),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1316),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1341),
.B(n_962),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1348),
.B(n_1255),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1341),
.B(n_933),
.Y(n_1725)
);

BUFx12f_ASAP7_75t_SL g1726 ( 
.A(n_1377),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1317),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_SL g1728 ( 
.A(n_1491),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1320),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1460),
.Y(n_1730)
);

OAI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1420),
.A2(n_941),
.B1(n_952),
.B2(n_938),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1487),
.B(n_941),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1489),
.B(n_952),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1351),
.B(n_954),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1407),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1408),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1444),
.B(n_954),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1495),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1412),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1422),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1464),
.Y(n_1741)
);

INVxp33_ASAP7_75t_L g1742 ( 
.A(n_1456),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1414),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1427),
.B(n_955),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1430),
.B(n_955),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1351),
.B(n_812),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1338),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1349),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_SL g1749 ( 
.A(n_1491),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1532),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1538),
.Y(n_1751)
);

INVx2_ASAP7_75t_SL g1752 ( 
.A(n_1516),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1338),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1411),
.B(n_670),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1444),
.B(n_671),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1498),
.B(n_682),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1479),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1349),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1413),
.B(n_869),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1552),
.B(n_684),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1480),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1555),
.A2(n_1566),
.B1(n_1415),
.B2(n_1513),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1573),
.B(n_924),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1502),
.B(n_688),
.Y(n_1764)
);

INVxp67_ASAP7_75t_SL g1765 ( 
.A(n_1497),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1391),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1566),
.A2(n_931),
.B1(n_937),
.B2(n_925),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_L g1768 ( 
.A(n_1325),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1502),
.B(n_689),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1349),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1381),
.B(n_691),
.Y(n_1771)
);

AO22x1_ASAP7_75t_L g1772 ( 
.A1(n_1523),
.A2(n_1537),
.B1(n_1565),
.B2(n_1558),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1413),
.B(n_697),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1415),
.B(n_700),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1432),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1532),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1392),
.Y(n_1777)
);

NAND2xp33_ASAP7_75t_SL g1778 ( 
.A(n_1558),
.B(n_702),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1318),
.B(n_1390),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1369),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1536),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1318),
.B(n_703),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1433),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1566),
.A2(n_943),
.B1(n_946),
.B2(n_945),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1325),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_L g1786 ( 
.A(n_1390),
.B(n_705),
.C(n_704),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1441),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1509),
.B(n_712),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1399),
.Y(n_1789)
);

INVxp67_ASAP7_75t_L g1790 ( 
.A(n_1369),
.Y(n_1790)
);

NOR3xp33_ASAP7_75t_L g1791 ( 
.A(n_1417),
.B(n_1481),
.C(n_1450),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1400),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1394),
.B(n_716),
.Y(n_1793)
);

A2O1A1Ixp33_ASAP7_75t_L g1794 ( 
.A1(n_1466),
.A2(n_1435),
.B(n_1429),
.C(n_1452),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1465),
.B(n_718),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1518),
.B(n_719),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1485),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1405),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1517),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1524),
.B(n_721),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1462),
.B(n_723),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1465),
.B(n_724),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1467),
.B(n_727),
.Y(n_1803)
);

BUFx5_ASAP7_75t_L g1804 ( 
.A(n_1447),
.Y(n_1804)
);

NAND2xp33_ASAP7_75t_L g1805 ( 
.A(n_1526),
.B(n_729),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1517),
.B(n_736),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1345),
.A2(n_1377),
.B1(n_1449),
.B2(n_1401),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1425),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1520),
.B(n_739),
.Y(n_1809)
);

AO22x1_ASAP7_75t_L g1810 ( 
.A1(n_1565),
.A2(n_741),
.B1(n_748),
.B2(n_747),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1342),
.B(n_1355),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1424),
.B(n_749),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1438),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1528),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1472),
.B(n_750),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1528),
.B(n_753),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1531),
.B(n_758),
.Y(n_1817)
);

NOR3xp33_ASAP7_75t_L g1818 ( 
.A(n_1473),
.B(n_767),
.C(n_654),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1556),
.A2(n_762),
.B1(n_770),
.B2(n_759),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1531),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_1534),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1534),
.Y(n_1822)
);

NAND2x1p5_ASAP7_75t_L g1823 ( 
.A(n_1445),
.B(n_947),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1325),
.Y(n_1824)
);

NAND2xp33_ASAP7_75t_L g1825 ( 
.A(n_1526),
.B(n_772),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1506),
.B(n_779),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1337),
.B(n_781),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1448),
.B(n_776),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1353),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1506),
.B(n_784),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1448),
.B(n_786),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1337),
.B(n_787),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1553),
.Y(n_1833)
);

INVxp67_ASAP7_75t_L g1834 ( 
.A(n_1355),
.Y(n_1834)
);

AOI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1556),
.A2(n_797),
.B1(n_799),
.B2(n_798),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1402),
.B(n_1362),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1492),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1362),
.B(n_1372),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1372),
.B(n_805),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1388),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1388),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1388),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1345),
.A2(n_950),
.B1(n_953),
.B2(n_948),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1455),
.B(n_810),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1529),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1564),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1461),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1571),
.B(n_811),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1561),
.B(n_813),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1572),
.B(n_815),
.Y(n_1850)
);

BUFx2_ASAP7_75t_L g1851 ( 
.A(n_1475),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1540),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1461),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1568),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1510),
.B(n_816),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1510),
.B(n_817),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1500),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1569),
.Y(n_1858)
);

OAI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1561),
.A2(n_821),
.B1(n_824),
.B2(n_823),
.Y(n_1859)
);

OA22x2_ASAP7_75t_L g1860 ( 
.A1(n_1475),
.A2(n_865),
.B1(n_893),
.B2(n_796),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1459),
.B(n_1542),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1500),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1459),
.B(n_827),
.Y(n_1863)
);

INVxp67_ASAP7_75t_L g1864 ( 
.A(n_1329),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1542),
.B(n_1577),
.Y(n_1865)
);

BUFx5_ASAP7_75t_L g1866 ( 
.A(n_1447),
.Y(n_1866)
);

OR2x6_ASAP7_75t_L g1867 ( 
.A(n_1374),
.B(n_958),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1504),
.A2(n_1283),
.B(n_1267),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1482),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1468),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1575),
.B(n_829),
.Y(n_1871)
);

BUFx3_ASAP7_75t_L g1872 ( 
.A(n_1353),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1562),
.B(n_830),
.Y(n_1873)
);

OAI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1315),
.A2(n_959),
.B(n_951),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1353),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1600),
.A2(n_1576),
.B(n_1575),
.Y(n_1876)
);

BUFx6f_ASAP7_75t_L g1877 ( 
.A(n_1715),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1596),
.B(n_1519),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1596),
.B(n_1591),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1794),
.A2(n_1315),
.B(n_1367),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1591),
.B(n_1519),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1585),
.B(n_1333),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1612),
.B(n_1559),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1609),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1579),
.B(n_1356),
.Y(n_1885)
);

O2A1O1Ixp33_ASAP7_75t_SL g1886 ( 
.A1(n_1861),
.A2(n_1398),
.B(n_1367),
.C(n_1527),
.Y(n_1886)
);

CKINVDCx10_ASAP7_75t_R g1887 ( 
.A(n_1728),
.Y(n_1887)
);

NAND2x1p5_ASAP7_75t_L g1888 ( 
.A(n_1616),
.B(n_1536),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1611),
.B(n_1578),
.Y(n_1889)
);

O2A1O1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1836),
.A2(n_1431),
.B(n_1503),
.C(n_1545),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1603),
.Y(n_1891)
);

A2O1A1Ixp33_ASAP7_75t_L g1892 ( 
.A1(n_1836),
.A2(n_1359),
.B(n_1360),
.C(n_1330),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1762),
.A2(n_1458),
.B1(n_1442),
.B2(n_1551),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1578),
.B(n_1503),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1628),
.A2(n_1527),
.B1(n_1551),
.B2(n_1458),
.Y(n_1895)
);

INVx1_ASAP7_75t_SL g1896 ( 
.A(n_1628),
.Y(n_1896)
);

AO21x1_ASAP7_75t_L g1897 ( 
.A1(n_1840),
.A2(n_1398),
.B(n_1376),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1671),
.B(n_1442),
.Y(n_1898)
);

OAI21xp33_ASAP7_75t_SL g1899 ( 
.A1(n_1628),
.A2(n_1324),
.B(n_1322),
.Y(n_1899)
);

NOR2x1_ASAP7_75t_L g1900 ( 
.A(n_1656),
.B(n_1322),
.Y(n_1900)
);

OAI21x1_ASAP7_75t_L g1901 ( 
.A1(n_1868),
.A2(n_1637),
.B(n_1852),
.Y(n_1901)
);

NOR3xp33_ASAP7_75t_L g1902 ( 
.A(n_1698),
.B(n_835),
.C(n_832),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1625),
.Y(n_1903)
);

OR2x6_ASAP7_75t_SL g1904 ( 
.A(n_1605),
.B(n_1751),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1726),
.B(n_1442),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1629),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1584),
.B(n_1559),
.Y(n_1907)
);

OAI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1779),
.A2(n_1395),
.B(n_1393),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1767),
.A2(n_725),
.B1(n_790),
.B2(n_701),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1630),
.B(n_1634),
.Y(n_1910)
);

OAI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1779),
.A2(n_1340),
.B(n_1324),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1717),
.B(n_839),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1780),
.B(n_844),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1838),
.A2(n_1363),
.B(n_1361),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1740),
.B(n_845),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1790),
.B(n_846),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1648),
.Y(n_1917)
);

BUFx4f_ASAP7_75t_L g1918 ( 
.A(n_1635),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1865),
.A2(n_1375),
.B(n_1370),
.Y(n_1919)
);

BUFx4f_ASAP7_75t_L g1920 ( 
.A(n_1635),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1654),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1631),
.B(n_847),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1650),
.B(n_851),
.Y(n_1923)
);

BUFx6f_ASAP7_75t_L g1924 ( 
.A(n_1715),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1580),
.B(n_852),
.Y(n_1925)
);

A2O1A1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1853),
.A2(n_1370),
.B(n_1383),
.C(n_1353),
.Y(n_1926)
);

O2A1O1Ixp33_ASAP7_75t_L g1927 ( 
.A1(n_1838),
.A2(n_854),
.B(n_856),
.C(n_853),
.Y(n_1927)
);

INVx4_ASAP7_75t_L g1928 ( 
.A(n_1635),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1613),
.B(n_1615),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1674),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1651),
.B(n_857),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1645),
.B(n_1370),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1683),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1707),
.B(n_859),
.Y(n_1934)
);

BUFx6f_ASAP7_75t_L g1935 ( 
.A(n_1715),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1668),
.B(n_867),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1709),
.B(n_868),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1747),
.A2(n_1328),
.B(n_1447),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1712),
.B(n_870),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1718),
.B(n_872),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1720),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1735),
.B(n_873),
.Y(n_1942)
);

OAI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1753),
.A2(n_1328),
.B(n_1507),
.Y(n_1943)
);

A2O1A1Ixp33_ASAP7_75t_L g1944 ( 
.A1(n_1811),
.A2(n_1416),
.B(n_1383),
.C(n_725),
.Y(n_1944)
);

NOR2x1p5_ASAP7_75t_SL g1945 ( 
.A(n_1617),
.B(n_1507),
.Y(n_1945)
);

BUFx3_ASAP7_75t_L g1946 ( 
.A(n_1582),
.Y(n_1946)
);

AO21x1_ASAP7_75t_L g1947 ( 
.A1(n_1841),
.A2(n_1328),
.B(n_1507),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1768),
.Y(n_1948)
);

O2A1O1Ixp33_ASAP7_75t_L g1949 ( 
.A1(n_1642),
.A2(n_1507),
.B(n_1512),
.C(n_1328),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1677),
.B(n_1383),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1736),
.B(n_1739),
.Y(n_1951)
);

CKINVDCx10_ASAP7_75t_R g1952 ( 
.A(n_1728),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1743),
.B(n_1383),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1757),
.Y(n_1954)
);

AOI22xp33_ASAP7_75t_L g1955 ( 
.A1(n_1791),
.A2(n_1512),
.B1(n_1416),
.B2(n_725),
.Y(n_1955)
);

NOR3xp33_ASAP7_75t_L g1956 ( 
.A(n_1610),
.B(n_1512),
.C(n_1416),
.Y(n_1956)
);

NOR2xp67_ASAP7_75t_L g1957 ( 
.A(n_1622),
.B(n_11),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1595),
.B(n_1416),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1834),
.A2(n_725),
.B(n_790),
.C(n_701),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1828),
.B(n_12),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1604),
.A2(n_1511),
.B(n_1499),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1619),
.B(n_1512),
.Y(n_1962)
);

A2O1A1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1604),
.A2(n_725),
.B(n_790),
.C(n_701),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1643),
.A2(n_1512),
.B(n_1554),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1619),
.B(n_790),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1647),
.B(n_790),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1583),
.B(n_1599),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1647),
.B(n_1661),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_SL g1969 ( 
.A1(n_1681),
.A2(n_1546),
.B(n_1541),
.Y(n_1969)
);

BUFx3_ASAP7_75t_L g1970 ( 
.A(n_1582),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1606),
.B(n_1554),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1661),
.B(n_842),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1616),
.B(n_1554),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_L g1974 ( 
.A(n_1768),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1775),
.Y(n_1975)
);

BUFx12f_ASAP7_75t_L g1976 ( 
.A(n_1665),
.Y(n_1976)
);

BUFx3_ASAP7_75t_L g1977 ( 
.A(n_1597),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1607),
.B(n_1554),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1761),
.Y(n_1979)
);

BUFx2_ASAP7_75t_L g1980 ( 
.A(n_1656),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1669),
.B(n_842),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1669),
.B(n_842),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1688),
.B(n_842),
.Y(n_1983)
);

OAI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1643),
.A2(n_1574),
.B(n_1546),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1845),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1768),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1842),
.Y(n_1987)
);

A2O1A1Ixp33_ASAP7_75t_L g1988 ( 
.A1(n_1771),
.A2(n_908),
.B(n_963),
.C(n_883),
.Y(n_1988)
);

AOI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1694),
.A2(n_908),
.B1(n_963),
.B2(n_883),
.Y(n_1989)
);

AOI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1871),
.A2(n_1546),
.B(n_1541),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1688),
.B(n_1732),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1601),
.B(n_1574),
.Y(n_1992)
);

INVx3_ASAP7_75t_L g1993 ( 
.A(n_1785),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1784),
.A2(n_1703),
.B1(n_1843),
.B2(n_1807),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1783),
.Y(n_1995)
);

INVxp67_ASAP7_75t_L g1996 ( 
.A(n_1656),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1732),
.B(n_883),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1601),
.B(n_883),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1601),
.B(n_883),
.Y(n_1999)
);

A2O1A1Ixp33_ASAP7_75t_L g2000 ( 
.A1(n_1627),
.A2(n_1633),
.B(n_1847),
.C(n_1724),
.Y(n_2000)
);

AOI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1801),
.A2(n_963),
.B(n_908),
.Y(n_2001)
);

OAI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1786),
.A2(n_963),
.B(n_908),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1787),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1618),
.B(n_14),
.Y(n_2004)
);

AOI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1801),
.A2(n_471),
.B(n_470),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1733),
.B(n_15),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1626),
.B(n_16),
.Y(n_2007)
);

AOI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1803),
.A2(n_477),
.B(n_475),
.Y(n_2008)
);

O2A1O1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1793),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_2009)
);

AOI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1803),
.A2(n_481),
.B(n_479),
.Y(n_2010)
);

BUFx4f_ASAP7_75t_L g2011 ( 
.A(n_1693),
.Y(n_2011)
);

OAI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1857),
.A2(n_20),
.B(n_21),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1592),
.Y(n_2013)
);

INVxp67_ASAP7_75t_L g2014 ( 
.A(n_1693),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1815),
.A2(n_485),
.B(n_482),
.Y(n_2015)
);

BUFx2_ASAP7_75t_L g2016 ( 
.A(n_1693),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1733),
.B(n_21),
.Y(n_2017)
);

O2A1O1Ixp33_ASAP7_75t_L g2018 ( 
.A1(n_1697),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_2018)
);

CKINVDCx10_ASAP7_75t_R g2019 ( 
.A(n_1749),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_SL g2020 ( 
.A(n_1617),
.B(n_494),
.Y(n_2020)
);

AOI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1682),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_2021)
);

A2O1A1Ixp33_ASAP7_75t_L g2022 ( 
.A1(n_1874),
.A2(n_28),
.B(n_25),
.C(n_27),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1608),
.B(n_27),
.Y(n_2023)
);

INVx1_ASAP7_75t_SL g2024 ( 
.A(n_1823),
.Y(n_2024)
);

AOI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_1826),
.A2(n_497),
.B(n_495),
.Y(n_2025)
);

AOI21x1_ASAP7_75t_L g2026 ( 
.A1(n_1638),
.A2(n_501),
.B(n_498),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1593),
.Y(n_2027)
);

AOI21xp5_ASAP7_75t_L g2028 ( 
.A1(n_1830),
.A2(n_505),
.B(n_502),
.Y(n_2028)
);

AOI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_1716),
.A2(n_507),
.B(n_506),
.Y(n_2029)
);

AOI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1716),
.A2(n_513),
.B(n_512),
.Y(n_2030)
);

OAI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_1862),
.A2(n_28),
.B(n_29),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1666),
.B(n_29),
.Y(n_2032)
);

INVx3_ASAP7_75t_L g2033 ( 
.A(n_1785),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1594),
.A2(n_528),
.B(n_525),
.Y(n_2034)
);

AO21x1_ASAP7_75t_L g2035 ( 
.A1(n_1765),
.A2(n_531),
.B(n_529),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1744),
.B(n_31),
.Y(n_2036)
);

BUFx12f_ASAP7_75t_L g2037 ( 
.A(n_1672),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_1598),
.A2(n_533),
.B(n_532),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1744),
.B(n_1745),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1602),
.Y(n_2040)
);

A2O1A1Ixp33_ASAP7_75t_L g2041 ( 
.A1(n_1874),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1745),
.B(n_32),
.Y(n_2042)
);

AOI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1587),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2043)
);

NOR2xp67_ASAP7_75t_L g2044 ( 
.A(n_1655),
.B(n_37),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1723),
.B(n_38),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1652),
.Y(n_2046)
);

O2A1O1Ixp33_ASAP7_75t_L g2047 ( 
.A1(n_1701),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1723),
.B(n_39),
.Y(n_2048)
);

AOI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_1831),
.A2(n_535),
.B(n_534),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1725),
.B(n_40),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1686),
.B(n_41),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_1823),
.Y(n_2052)
);

BUFx4f_ASAP7_75t_L g2053 ( 
.A(n_1581),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1785),
.Y(n_2054)
);

AOI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_1702),
.A2(n_540),
.B(n_539),
.Y(n_2055)
);

O2A1O1Ixp33_ASAP7_75t_L g2056 ( 
.A1(n_1818),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1700),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1725),
.B(n_42),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1737),
.B(n_45),
.Y(n_2059)
);

OAI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1754),
.A2(n_45),
.B(n_46),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1680),
.B(n_46),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1714),
.B(n_47),
.Y(n_2062)
);

A2O1A1Ixp33_ASAP7_75t_L g2063 ( 
.A1(n_1719),
.A2(n_50),
.B(n_47),
.C(n_49),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1849),
.A2(n_550),
.B(n_544),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1808),
.Y(n_2065)
);

O2A1O1Ixp33_ASAP7_75t_L g2066 ( 
.A1(n_1855),
.A2(n_54),
.B(n_49),
.C(n_53),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1696),
.B(n_1839),
.Y(n_2067)
);

INVx1_ASAP7_75t_SL g2068 ( 
.A(n_1851),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1673),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1869),
.B(n_54),
.Y(n_2070)
);

NAND2xp33_ASAP7_75t_L g2071 ( 
.A(n_1617),
.B(n_551),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1774),
.B(n_55),
.Y(n_2072)
);

AND2x2_ASAP7_75t_SL g2073 ( 
.A(n_1805),
.B(n_55),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1839),
.B(n_56),
.Y(n_2074)
);

AOI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_1844),
.A2(n_553),
.B(n_552),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_1687),
.B(n_1738),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1855),
.B(n_57),
.Y(n_2077)
);

OAI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_1589),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1856),
.B(n_60),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_1752),
.B(n_61),
.Y(n_2080)
);

AOI21xp5_ASAP7_75t_L g2081 ( 
.A1(n_1766),
.A2(n_559),
.B(n_558),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_1870),
.A2(n_64),
.B1(n_61),
.B2(n_62),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1856),
.B(n_62),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_1875),
.B(n_64),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1641),
.B(n_65),
.Y(n_2085)
);

INVx3_ASAP7_75t_L g2086 ( 
.A(n_1824),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1813),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1644),
.B(n_69),
.Y(n_2088)
);

AOI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_1777),
.A2(n_564),
.B(n_562),
.Y(n_2089)
);

NOR2xp67_ASAP7_75t_L g2090 ( 
.A(n_1657),
.B(n_72),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1673),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_1705),
.B(n_73),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1756),
.B(n_73),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_1749),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1588),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1756),
.B(n_74),
.Y(n_2096)
);

AOI21xp5_ASAP7_75t_L g2097 ( 
.A1(n_1789),
.A2(n_570),
.B(n_568),
.Y(n_2097)
);

INVx3_ASAP7_75t_L g2098 ( 
.A(n_1824),
.Y(n_2098)
);

HB1xp67_ASAP7_75t_L g2099 ( 
.A(n_1667),
.Y(n_2099)
);

AND2x6_ASAP7_75t_L g2100 ( 
.A(n_1695),
.B(n_74),
.Y(n_2100)
);

INVx5_ASAP7_75t_L g2101 ( 
.A(n_1824),
.Y(n_2101)
);

O2A1O1Ixp33_ASAP7_75t_L g2102 ( 
.A1(n_1800),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1763),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1792),
.B(n_75),
.Y(n_2104)
);

AND2x2_ASAP7_75t_SL g2105 ( 
.A(n_1825),
.B(n_1640),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1798),
.B(n_76),
.Y(n_2106)
);

AOI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_1664),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_2107)
);

NOR2xp67_ASAP7_75t_L g2108 ( 
.A(n_1708),
.B(n_78),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1800),
.B(n_80),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1679),
.B(n_1684),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_1721),
.B(n_81),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_1812),
.A2(n_575),
.B(n_572),
.Y(n_2112)
);

BUFx6f_ASAP7_75t_L g2113 ( 
.A(n_1829),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1649),
.B(n_81),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1764),
.B(n_82),
.Y(n_2115)
);

AND2x4_ASAP7_75t_SL g2116 ( 
.A(n_1829),
.B(n_84),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1763),
.Y(n_2117)
);

OAI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_1827),
.A2(n_1832),
.B(n_1782),
.Y(n_2118)
);

A2O1A1Ixp33_ASAP7_75t_L g2119 ( 
.A1(n_1675),
.A2(n_1788),
.B(n_1796),
.C(n_1863),
.Y(n_2119)
);

NAND2x1p5_ASAP7_75t_L g2120 ( 
.A(n_1829),
.B(n_1875),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_R g2121 ( 
.A(n_1778),
.B(n_85),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_L g2122 ( 
.A(n_1755),
.B(n_85),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1875),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1859),
.B(n_86),
.Y(n_2124)
);

INVx3_ASAP7_75t_L g2125 ( 
.A(n_1658),
.Y(n_2125)
);

BUFx8_ASAP7_75t_L g2126 ( 
.A(n_1797),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1590),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1863),
.A2(n_584),
.B(n_577),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1769),
.B(n_1774),
.Y(n_2129)
);

NAND2x1p5_ASAP7_75t_L g2130 ( 
.A(n_1658),
.B(n_87),
.Y(n_2130)
);

O2A1O1Ixp33_ASAP7_75t_L g2131 ( 
.A1(n_1731),
.A2(n_91),
.B(n_88),
.C(n_90),
.Y(n_2131)
);

INVx4_ASAP7_75t_L g2132 ( 
.A(n_1695),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1806),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_1581),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1864),
.B(n_90),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1799),
.B(n_91),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1814),
.B(n_92),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1806),
.Y(n_2138)
);

OAI21xp5_ASAP7_75t_L g2139 ( 
.A1(n_1827),
.A2(n_93),
.B(n_94),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1809),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1820),
.B(n_95),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1833),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_SL g2143 ( 
.A(n_1695),
.B(n_96),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_1676),
.Y(n_2144)
);

OAI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_1832),
.A2(n_96),
.B(n_97),
.Y(n_2145)
);

AOI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_1846),
.A2(n_590),
.B(n_594),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1782),
.B(n_97),
.Y(n_2147)
);

OAI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_1730),
.A2(n_98),
.B(n_99),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1809),
.Y(n_2149)
);

AOI21xp5_ASAP7_75t_L g2150 ( 
.A1(n_1854),
.A2(n_98),
.B(n_99),
.Y(n_2150)
);

AOI21xp5_ASAP7_75t_L g2151 ( 
.A1(n_1858),
.A2(n_100),
.B(n_102),
.Y(n_2151)
);

OAI21xp5_ASAP7_75t_L g2152 ( 
.A1(n_1741),
.A2(n_1727),
.B(n_1722),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1816),
.B(n_100),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1816),
.B(n_102),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1817),
.B(n_103),
.Y(n_2155)
);

CKINVDCx6p67_ASAP7_75t_R g2156 ( 
.A(n_1867),
.Y(n_2156)
);

AOI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_1586),
.A2(n_106),
.B(n_107),
.Y(n_2157)
);

OAI22xp5_ASAP7_75t_L g2158 ( 
.A1(n_1860),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1760),
.B(n_109),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1729),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1710),
.Y(n_2161)
);

AO21x1_ASAP7_75t_L g2162 ( 
.A1(n_1713),
.A2(n_109),
.B(n_110),
.Y(n_2162)
);

INVx3_ASAP7_75t_L g2163 ( 
.A(n_1676),
.Y(n_2163)
);

AOI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_1653),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_2164)
);

A2O1A1Ixp33_ASAP7_75t_L g2165 ( 
.A1(n_1711),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_2165)
);

OR2x2_ASAP7_75t_L g2166 ( 
.A(n_1819),
.B(n_114),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1867),
.B(n_116),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1867),
.B(n_117),
.Y(n_2168)
);

AOI21xp5_ASAP7_75t_L g2169 ( 
.A1(n_1614),
.A2(n_119),
.B(n_120),
.Y(n_2169)
);

AOI21x1_ASAP7_75t_L g2170 ( 
.A1(n_1620),
.A2(n_120),
.B(n_121),
.Y(n_2170)
);

BUFx4f_ASAP7_75t_L g2171 ( 
.A(n_1636),
.Y(n_2171)
);

AOI21xp5_ASAP7_75t_L g2172 ( 
.A1(n_1639),
.A2(n_123),
.B(n_125),
.Y(n_2172)
);

AOI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_1660),
.A2(n_123),
.B(n_125),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_1662),
.A2(n_126),
.B(n_127),
.Y(n_2174)
);

OAI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_1663),
.A2(n_126),
.B(n_128),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_1632),
.B(n_1837),
.Y(n_2176)
);

AOI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_1670),
.A2(n_128),
.B(n_129),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1632),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_1632),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1835),
.B(n_129),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_1872),
.B(n_130),
.Y(n_2181)
);

AOI21xp5_ASAP7_75t_L g2182 ( 
.A1(n_1689),
.A2(n_130),
.B(n_131),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_1623),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_2183)
);

OAI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_1690),
.A2(n_132),
.B(n_133),
.Y(n_2184)
);

A2O1A1Ixp33_ASAP7_75t_L g2185 ( 
.A1(n_1692),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1699),
.Y(n_2186)
);

AND2x2_ASAP7_75t_SL g2187 ( 
.A(n_1646),
.B(n_135),
.Y(n_2187)
);

AOI21xp5_ASAP7_75t_L g2188 ( 
.A1(n_1704),
.A2(n_137),
.B(n_138),
.Y(n_2188)
);

AO21x1_ASAP7_75t_L g2189 ( 
.A1(n_1746),
.A2(n_138),
.B(n_139),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1821),
.Y(n_2190)
);

AOI21xp5_ASAP7_75t_L g2191 ( 
.A1(n_1822),
.A2(n_140),
.B(n_141),
.Y(n_2191)
);

BUFx4f_ASAP7_75t_L g2192 ( 
.A(n_1636),
.Y(n_2192)
);

A2O1A1Ixp33_ASAP7_75t_L g2193 ( 
.A1(n_1873),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_2193)
);

AOI21xp33_ASAP7_75t_L g2194 ( 
.A1(n_1621),
.A2(n_142),
.B(n_146),
.Y(n_2194)
);

AOI21xp5_ASAP7_75t_L g2195 ( 
.A1(n_1678),
.A2(n_147),
.B(n_148),
.Y(n_2195)
);

AOI21xp5_ASAP7_75t_L g2196 ( 
.A1(n_1691),
.A2(n_148),
.B(n_149),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1734),
.Y(n_2197)
);

OAI21xp5_ASAP7_75t_L g2198 ( 
.A1(n_1706),
.A2(n_150),
.B(n_151),
.Y(n_2198)
);

A2O1A1Ixp33_ASAP7_75t_L g2199 ( 
.A1(n_1848),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_1742),
.B(n_152),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1659),
.Y(n_2201)
);

AND2x4_ASAP7_75t_L g2202 ( 
.A(n_1659),
.B(n_153),
.Y(n_2202)
);

NAND2xp33_ASAP7_75t_L g2203 ( 
.A(n_1866),
.B(n_153),
.Y(n_2203)
);

AOI21xp5_ASAP7_75t_L g2204 ( 
.A1(n_1748),
.A2(n_154),
.B(n_155),
.Y(n_2204)
);

A2O1A1Ixp33_ASAP7_75t_L g2205 ( 
.A1(n_1850),
.A2(n_158),
.B(n_154),
.C(n_157),
.Y(n_2205)
);

AO21x1_ASAP7_75t_L g2206 ( 
.A1(n_1759),
.A2(n_1795),
.B(n_1773),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_1750),
.B(n_159),
.Y(n_2207)
);

INVxp67_ASAP7_75t_L g2208 ( 
.A(n_1810),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_1776),
.B(n_159),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1772),
.B(n_160),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1879),
.B(n_1802),
.Y(n_2211)
);

BUFx6f_ASAP7_75t_L g2212 ( 
.A(n_2101),
.Y(n_2212)
);

AO21x2_ASAP7_75t_L g2213 ( 
.A1(n_1911),
.A2(n_1770),
.B(n_1758),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1884),
.B(n_1781),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_2011),
.B(n_1617),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1889),
.B(n_1781),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_1967),
.B(n_161),
.Y(n_2217)
);

OAI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_1898),
.A2(n_1621),
.B1(n_1624),
.B2(n_1617),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1878),
.B(n_1624),
.Y(n_2219)
);

OAI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_1898),
.A2(n_1685),
.B1(n_1804),
.B2(n_1617),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2156),
.B(n_162),
.Y(n_2221)
);

O2A1O1Ixp33_ASAP7_75t_L g2222 ( 
.A1(n_2119),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1881),
.B(n_1968),
.Y(n_2223)
);

NOR3xp33_ASAP7_75t_SL g2224 ( 
.A(n_2094),
.B(n_163),
.C(n_165),
.Y(n_2224)
);

BUFx2_ASAP7_75t_L g2225 ( 
.A(n_1918),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1991),
.B(n_165),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2039),
.B(n_166),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2129),
.B(n_167),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2110),
.B(n_168),
.Y(n_2229)
);

NAND3xp33_ASAP7_75t_L g2230 ( 
.A(n_2183),
.B(n_1804),
.C(n_1685),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2110),
.B(n_169),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1921),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_2011),
.B(n_1685),
.Y(n_2233)
);

AND2x4_ASAP7_75t_L g2234 ( 
.A(n_1928),
.B(n_169),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2133),
.B(n_170),
.Y(n_2235)
);

BUFx8_ASAP7_75t_SL g2236 ( 
.A(n_1976),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_1896),
.B(n_170),
.Y(n_2237)
);

BUFx2_ASAP7_75t_R g2238 ( 
.A(n_1904),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1930),
.Y(n_2239)
);

BUFx3_ASAP7_75t_L g2240 ( 
.A(n_2126),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1933),
.Y(n_2241)
);

CKINVDCx20_ASAP7_75t_R g2242 ( 
.A(n_1946),
.Y(n_2242)
);

O2A1O1Ixp33_ASAP7_75t_L g2243 ( 
.A1(n_2056),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_2243)
);

AO221x2_ASAP7_75t_L g2244 ( 
.A1(n_2158),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.C(n_177),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_2073),
.B(n_2024),
.Y(n_2245)
);

HB1xp67_ASAP7_75t_L g2246 ( 
.A(n_1891),
.Y(n_2246)
);

INVx3_ASAP7_75t_L g2247 ( 
.A(n_2053),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_1939),
.B(n_175),
.Y(n_2248)
);

NAND3xp33_ASAP7_75t_SL g2249 ( 
.A(n_2121),
.B(n_2158),
.C(n_2043),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2138),
.B(n_176),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_1876),
.A2(n_1866),
.B(n_178),
.Y(n_2251)
);

BUFx2_ASAP7_75t_L g2252 ( 
.A(n_1918),
.Y(n_2252)
);

OAI22xp5_ASAP7_75t_SL g2253 ( 
.A1(n_2105),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_2253)
);

O2A1O1Ixp33_ASAP7_75t_L g2254 ( 
.A1(n_2159),
.A2(n_185),
.B(n_182),
.C(n_183),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_1920),
.Y(n_2255)
);

NAND2xp33_ASAP7_75t_SL g2256 ( 
.A(n_1928),
.B(n_182),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2140),
.B(n_183),
.Y(n_2257)
);

BUFx3_ASAP7_75t_L g2258 ( 
.A(n_2126),
.Y(n_2258)
);

A2O1A1Ixp33_ASAP7_75t_L g2259 ( 
.A1(n_1890),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_2259)
);

OAI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_2004),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2149),
.B(n_188),
.Y(n_2261)
);

INVx2_ASAP7_75t_SL g2262 ( 
.A(n_1920),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2053),
.B(n_189),
.Y(n_2263)
);

OAI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_1960),
.A2(n_193),
.B1(n_190),
.B2(n_191),
.Y(n_2264)
);

AOI21x1_ASAP7_75t_L g2265 ( 
.A1(n_2026),
.A2(n_191),
.B(n_193),
.Y(n_2265)
);

NAND3xp33_ASAP7_75t_L g2266 ( 
.A(n_1988),
.B(n_194),
.C(n_196),
.Y(n_2266)
);

AOI21xp5_ASAP7_75t_L g2267 ( 
.A1(n_1990),
.A2(n_197),
.B(n_198),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1910),
.B(n_197),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_1912),
.B(n_198),
.Y(n_2269)
);

AOI33xp33_ASAP7_75t_L g2270 ( 
.A1(n_2051),
.A2(n_199),
.A3(n_202),
.B1(n_203),
.B2(n_204),
.B3(n_205),
.Y(n_2270)
);

NOR2xp33_ASAP7_75t_SL g2271 ( 
.A(n_2020),
.B(n_202),
.Y(n_2271)
);

A2O1A1Ixp33_ASAP7_75t_L g2272 ( 
.A1(n_2059),
.A2(n_210),
.B(n_206),
.C(n_209),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1941),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1903),
.Y(n_2274)
);

BUFx6f_ASAP7_75t_L g2275 ( 
.A(n_2101),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1910),
.B(n_210),
.Y(n_2276)
);

AOI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2023),
.A2(n_214),
.B1(n_211),
.B2(n_213),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1906),
.Y(n_2278)
);

BUFx6f_ASAP7_75t_L g2279 ( 
.A(n_2101),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1917),
.Y(n_2280)
);

NOR2xp33_ASAP7_75t_L g2281 ( 
.A(n_1915),
.B(n_214),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_2101),
.B(n_216),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2052),
.B(n_216),
.Y(n_2283)
);

AOI33xp33_ASAP7_75t_L g2284 ( 
.A1(n_1985),
.A2(n_217),
.A3(n_219),
.B1(n_220),
.B2(n_222),
.B3(n_223),
.Y(n_2284)
);

O2A1O1Ixp33_ASAP7_75t_L g2285 ( 
.A1(n_1902),
.A2(n_224),
.B(n_219),
.C(n_220),
.Y(n_2285)
);

O2A1O1Ixp33_ASAP7_75t_L g2286 ( 
.A1(n_1927),
.A2(n_227),
.B(n_225),
.C(n_226),
.Y(n_2286)
);

AOI21xp5_ASAP7_75t_L g2287 ( 
.A1(n_1961),
.A2(n_225),
.B(n_226),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1954),
.Y(n_2288)
);

A2O1A1Ixp33_ASAP7_75t_L g2289 ( 
.A1(n_2122),
.A2(n_231),
.B(n_229),
.C(n_230),
.Y(n_2289)
);

AOI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_1994),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1979),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_1887),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_1886),
.A2(n_232),
.B(n_233),
.Y(n_2293)
);

NAND3xp33_ASAP7_75t_SL g2294 ( 
.A(n_2107),
.B(n_234),
.C(n_235),
.Y(n_2294)
);

BUFx3_ASAP7_75t_L g2295 ( 
.A(n_1970),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2208),
.B(n_1923),
.Y(n_2296)
);

O2A1O1Ixp5_ASAP7_75t_L g2297 ( 
.A1(n_2002),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1951),
.B(n_237),
.Y(n_2298)
);

CKINVDCx16_ASAP7_75t_R g2299 ( 
.A(n_2037),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_2068),
.B(n_241),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_1929),
.B(n_242),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2068),
.B(n_245),
.Y(n_2302)
);

BUFx6f_ASAP7_75t_L g2303 ( 
.A(n_1877),
.Y(n_2303)
);

BUFx12f_ASAP7_75t_L g2304 ( 
.A(n_1977),
.Y(n_2304)
);

HB1xp67_ASAP7_75t_L g2305 ( 
.A(n_2181),
.Y(n_2305)
);

BUFx3_ASAP7_75t_L g2306 ( 
.A(n_2181),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2127),
.Y(n_2307)
);

NAND2xp33_ASAP7_75t_L g2308 ( 
.A(n_2100),
.B(n_245),
.Y(n_2308)
);

OR2x6_ASAP7_75t_L g2309 ( 
.A(n_2202),
.B(n_246),
.Y(n_2309)
);

AO32x1_ASAP7_75t_L g2310 ( 
.A1(n_2078),
.A2(n_1893),
.A3(n_2082),
.B1(n_1909),
.B2(n_1987),
.Y(n_2310)
);

AOI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_1880),
.A2(n_247),
.B(n_248),
.Y(n_2311)
);

NAND2xp33_ASAP7_75t_L g2312 ( 
.A(n_2100),
.B(n_247),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_1975),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2095),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2202),
.B(n_249),
.Y(n_2315)
);

OR2x2_ASAP7_75t_L g2316 ( 
.A(n_1922),
.B(n_250),
.Y(n_2316)
);

OAI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_2092),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1995),
.Y(n_2318)
);

OAI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_2114),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_1877),
.B(n_254),
.Y(n_2320)
);

OAI22xp5_ASAP7_75t_L g2321 ( 
.A1(n_2114),
.A2(n_2130),
.B1(n_2067),
.B2(n_2070),
.Y(n_2321)
);

O2A1O1Ixp33_ASAP7_75t_L g2322 ( 
.A1(n_2167),
.A2(n_255),
.B(n_256),
.C(n_259),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2104),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2057),
.B(n_255),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_SL g2325 ( 
.A(n_1877),
.B(n_259),
.Y(n_2325)
);

OAI22xp5_ASAP7_75t_L g2326 ( 
.A1(n_2130),
.A2(n_260),
.B1(n_261),
.B2(n_265),
.Y(n_2326)
);

AOI22xp33_ASAP7_75t_L g2327 ( 
.A1(n_1994),
.A2(n_260),
.B1(n_261),
.B2(n_265),
.Y(n_2327)
);

A2O1A1Ixp33_ASAP7_75t_L g2328 ( 
.A1(n_2131),
.A2(n_266),
.B(n_268),
.C(n_269),
.Y(n_2328)
);

INVx3_ASAP7_75t_L g2329 ( 
.A(n_1973),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2046),
.B(n_266),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_SL g2331 ( 
.A(n_1924),
.B(n_268),
.Y(n_2331)
);

INVx3_ASAP7_75t_SL g2332 ( 
.A(n_2100),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2013),
.B(n_2027),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_L g2334 ( 
.A(n_1929),
.B(n_269),
.Y(n_2334)
);

O2A1O1Ixp33_ASAP7_75t_SL g2335 ( 
.A1(n_1944),
.A2(n_1964),
.B(n_1926),
.C(n_2000),
.Y(n_2335)
);

AOI21xp5_ASAP7_75t_L g2336 ( 
.A1(n_1965),
.A2(n_270),
.B(n_271),
.Y(n_2336)
);

INVx2_ASAP7_75t_SL g2337 ( 
.A(n_1952),
.Y(n_2337)
);

O2A1O1Ixp33_ASAP7_75t_L g2338 ( 
.A1(n_2168),
.A2(n_270),
.B(n_271),
.C(n_273),
.Y(n_2338)
);

A2O1A1Ixp33_ASAP7_75t_L g2339 ( 
.A1(n_2060),
.A2(n_273),
.B(n_274),
.C(n_275),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2040),
.B(n_275),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2072),
.B(n_276),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2103),
.B(n_276),
.Y(n_2342)
);

INVx4_ASAP7_75t_L g2343 ( 
.A(n_2100),
.Y(n_2343)
);

AOI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_1966),
.A2(n_278),
.B(n_279),
.Y(n_2344)
);

INVx3_ASAP7_75t_L g2345 ( 
.A(n_1973),
.Y(n_2345)
);

AOI21xp5_ASAP7_75t_L g2346 ( 
.A1(n_1972),
.A2(n_278),
.B(n_280),
.Y(n_2346)
);

INVxp67_ASAP7_75t_L g2347 ( 
.A(n_2080),
.Y(n_2347)
);

OAI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_2109),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2117),
.B(n_283),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2007),
.B(n_1925),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_L g2351 ( 
.A(n_1936),
.B(n_284),
.Y(n_2351)
);

AOI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_2044),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2080),
.B(n_286),
.Y(n_2353)
);

INVx2_ASAP7_75t_SL g2354 ( 
.A(n_2019),
.Y(n_2354)
);

INVx5_ASAP7_75t_L g2355 ( 
.A(n_1924),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2070),
.B(n_289),
.Y(n_2356)
);

NAND2x1p5_ASAP7_75t_L g2357 ( 
.A(n_2171),
.B(n_289),
.Y(n_2357)
);

BUFx6f_ASAP7_75t_L g2358 ( 
.A(n_1924),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_1931),
.B(n_290),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_1935),
.Y(n_2360)
);

INVx3_ASAP7_75t_L g2361 ( 
.A(n_1888),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2104),
.Y(n_2362)
);

INVxp67_ASAP7_75t_L g2363 ( 
.A(n_2108),
.Y(n_2363)
);

OA22x2_ASAP7_75t_L g2364 ( 
.A1(n_2082),
.A2(n_2116),
.B1(n_2021),
.B2(n_2148),
.Y(n_2364)
);

AOI21xp5_ASAP7_75t_L g2365 ( 
.A1(n_1981),
.A2(n_291),
.B(n_292),
.Y(n_2365)
);

BUFx3_ASAP7_75t_L g2366 ( 
.A(n_2120),
.Y(n_2366)
);

NOR2x1_ASAP7_75t_L g2367 ( 
.A(n_2175),
.B(n_2184),
.Y(n_2367)
);

AOI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2166),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_2368)
);

AOI21xp5_ASAP7_75t_L g2369 ( 
.A1(n_1982),
.A2(n_294),
.B(n_297),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_L g2370 ( 
.A(n_2200),
.B(n_294),
.Y(n_2370)
);

AO31x2_ASAP7_75t_L g2371 ( 
.A1(n_1897),
.A2(n_297),
.A3(n_298),
.B(n_299),
.Y(n_2371)
);

NOR3xp33_ASAP7_75t_SL g2372 ( 
.A(n_2199),
.B(n_298),
.C(n_299),
.Y(n_2372)
);

AOI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_1983),
.A2(n_300),
.B(n_301),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2003),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2109),
.B(n_1894),
.Y(n_2375)
);

BUFx2_ASAP7_75t_L g2376 ( 
.A(n_1980),
.Y(n_2376)
);

INVx4_ASAP7_75t_L g2377 ( 
.A(n_1935),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_1913),
.B(n_302),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2106),
.Y(n_2379)
);

OAI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_1984),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_2380)
);

O2A1O1Ixp33_ASAP7_75t_L g2381 ( 
.A1(n_2180),
.A2(n_304),
.B(n_305),
.C(n_307),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_R g2382 ( 
.A(n_2203),
.B(n_309),
.Y(n_2382)
);

INVx8_ASAP7_75t_L g2383 ( 
.A(n_1935),
.Y(n_2383)
);

AOI21xp5_ASAP7_75t_L g2384 ( 
.A1(n_1997),
.A2(n_310),
.B(n_311),
.Y(n_2384)
);

AND2x4_ASAP7_75t_L g2385 ( 
.A(n_2134),
.B(n_310),
.Y(n_2385)
);

OAI22xp5_ASAP7_75t_L g2386 ( 
.A1(n_1984),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2106),
.Y(n_2387)
);

OR2x6_ASAP7_75t_L g2388 ( 
.A(n_2016),
.B(n_314),
.Y(n_2388)
);

OAI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_2115),
.A2(n_1893),
.B1(n_2078),
.B2(n_1909),
.Y(n_2389)
);

NOR2xp67_ASAP7_75t_SL g2390 ( 
.A(n_2099),
.B(n_315),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2136),
.Y(n_2391)
);

NAND3xp33_ASAP7_75t_L g2392 ( 
.A(n_1963),
.B(n_316),
.C(n_317),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2061),
.B(n_317),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2142),
.Y(n_2394)
);

INVx3_ASAP7_75t_SL g2395 ( 
.A(n_2076),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_1916),
.B(n_318),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2032),
.B(n_318),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2065),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2006),
.B(n_319),
.Y(n_2399)
);

BUFx12f_ASAP7_75t_L g2400 ( 
.A(n_2076),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_SL g2401 ( 
.A(n_2020),
.B(n_319),
.Y(n_2401)
);

INVx2_ASAP7_75t_SL g2402 ( 
.A(n_2171),
.Y(n_2402)
);

NOR2xp33_ASAP7_75t_SL g2403 ( 
.A(n_1964),
.B(n_320),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2087),
.Y(n_2404)
);

O2A1O1Ixp33_ASAP7_75t_L g2405 ( 
.A1(n_2205),
.A2(n_321),
.B(n_322),
.C(n_323),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2017),
.B(n_321),
.Y(n_2406)
);

AOI21xp5_ASAP7_75t_L g2407 ( 
.A1(n_2118),
.A2(n_323),
.B(n_324),
.Y(n_2407)
);

INVx2_ASAP7_75t_SL g2408 ( 
.A(n_2192),
.Y(n_2408)
);

NOR3xp33_ASAP7_75t_SL g2409 ( 
.A(n_2193),
.B(n_324),
.C(n_325),
.Y(n_2409)
);

NOR3xp33_ASAP7_75t_SL g2410 ( 
.A(n_2135),
.B(n_325),
.C(n_327),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2036),
.B(n_327),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2042),
.B(n_328),
.Y(n_2412)
);

AOI21xp5_ASAP7_75t_L g2413 ( 
.A1(n_1908),
.A2(n_329),
.B(n_330),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2136),
.Y(n_2414)
);

O2A1O1Ixp33_ASAP7_75t_L g2415 ( 
.A1(n_2124),
.A2(n_329),
.B(n_330),
.C(n_331),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2137),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_SL g2417 ( 
.A(n_1948),
.B(n_332),
.Y(n_2417)
);

OAI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_2115),
.A2(n_333),
.B1(n_334),
.B2(n_336),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2137),
.Y(n_2419)
);

INVx3_ASAP7_75t_L g2420 ( 
.A(n_1888),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2160),
.Y(n_2421)
);

OAI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2045),
.A2(n_333),
.B1(n_334),
.B2(n_336),
.Y(n_2422)
);

O2A1O1Ixp33_ASAP7_75t_L g2423 ( 
.A1(n_2048),
.A2(n_337),
.B(n_339),
.C(n_340),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_1996),
.B(n_337),
.Y(n_2424)
);

AND2x4_ASAP7_75t_L g2425 ( 
.A(n_2132),
.B(n_339),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2141),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2141),
.Y(n_2427)
);

BUFx2_ASAP7_75t_L g2428 ( 
.A(n_2120),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_SL g2429 ( 
.A(n_1948),
.B(n_341),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_SL g2430 ( 
.A(n_1948),
.B(n_342),
.Y(n_2430)
);

CKINVDCx5p33_ASAP7_75t_R g2431 ( 
.A(n_1905),
.Y(n_2431)
);

BUFx6f_ASAP7_75t_L g2432 ( 
.A(n_1974),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2186),
.Y(n_2433)
);

OAI21xp5_ASAP7_75t_L g2434 ( 
.A1(n_2147),
.A2(n_343),
.B(n_344),
.Y(n_2434)
);

NAND2x1p5_ASAP7_75t_L g2435 ( 
.A(n_2192),
.B(n_345),
.Y(n_2435)
);

BUFx2_ASAP7_75t_L g2436 ( 
.A(n_1993),
.Y(n_2436)
);

O2A1O1Ixp33_ASAP7_75t_L g2437 ( 
.A1(n_2050),
.A2(n_346),
.B(n_347),
.C(n_348),
.Y(n_2437)
);

NOR2xp33_ASAP7_75t_L g2438 ( 
.A(n_2014),
.B(n_347),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_1885),
.B(n_348),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_L g2440 ( 
.A(n_1934),
.B(n_349),
.Y(n_2440)
);

AOI22xp33_ASAP7_75t_L g2441 ( 
.A1(n_2111),
.A2(n_350),
.B1(n_351),
.B2(n_353),
.Y(n_2441)
);

BUFx6f_ASAP7_75t_L g2442 ( 
.A(n_1974),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_SL g2443 ( 
.A(n_1974),
.B(n_351),
.Y(n_2443)
);

AOI22xp33_ASAP7_75t_L g2444 ( 
.A1(n_2077),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_2444)
);

INVx3_ASAP7_75t_SL g2445 ( 
.A(n_1986),
.Y(n_2445)
);

BUFx3_ASAP7_75t_L g2446 ( 
.A(n_1986),
.Y(n_2446)
);

O2A1O1Ixp33_ASAP7_75t_L g2447 ( 
.A1(n_2058),
.A2(n_357),
.B(n_358),
.C(n_360),
.Y(n_2447)
);

A2O1A1Ixp33_ASAP7_75t_L g2448 ( 
.A1(n_2060),
.A2(n_357),
.B(n_358),
.C(n_361),
.Y(n_2448)
);

OAI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_2147),
.A2(n_361),
.B1(n_362),
.B2(n_363),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2209),
.Y(n_2450)
);

BUFx2_ASAP7_75t_L g2451 ( 
.A(n_1993),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_1986),
.B(n_2054),
.Y(n_2452)
);

NOR2xp33_ASAP7_75t_R g2453 ( 
.A(n_2054),
.B(n_362),
.Y(n_2453)
);

CKINVDCx6p67_ASAP7_75t_R g2454 ( 
.A(n_2054),
.Y(n_2454)
);

NAND2xp33_ASAP7_75t_L g2455 ( 
.A(n_2113),
.B(n_364),
.Y(n_2455)
);

AO21x1_ASAP7_75t_L g2456 ( 
.A1(n_2198),
.A2(n_364),
.B(n_365),
.Y(n_2456)
);

AOI21xp5_ASAP7_75t_L g2457 ( 
.A1(n_1901),
.A2(n_365),
.B(n_366),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_1937),
.B(n_367),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_1940),
.B(n_367),
.Y(n_2459)
);

AOI21xp5_ASAP7_75t_L g2460 ( 
.A1(n_1914),
.A2(n_368),
.B(n_369),
.Y(n_2460)
);

INVx2_ASAP7_75t_SL g2461 ( 
.A(n_2113),
.Y(n_2461)
);

AOI21xp5_ASAP7_75t_L g2462 ( 
.A1(n_1914),
.A2(n_371),
.B(n_372),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_2113),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_1942),
.B(n_372),
.Y(n_2464)
);

OAI22xp5_ASAP7_75t_L g2465 ( 
.A1(n_2079),
.A2(n_373),
.B1(n_374),
.B2(n_376),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2083),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_1882),
.B(n_374),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2093),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2085),
.B(n_378),
.Y(n_2469)
);

BUFx8_ASAP7_75t_L g2470 ( 
.A(n_2197),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2096),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_SL g2472 ( 
.A(n_2123),
.B(n_2187),
.Y(n_2472)
);

AOI21xp5_ASAP7_75t_L g2473 ( 
.A1(n_2001),
.A2(n_379),
.B(n_380),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2069),
.B(n_379),
.Y(n_2474)
);

AOI21xp33_ASAP7_75t_L g2475 ( 
.A1(n_1899),
.A2(n_380),
.B(n_381),
.Y(n_2475)
);

O2A1O1Ixp5_ASAP7_75t_L g2476 ( 
.A1(n_2002),
.A2(n_382),
.B(n_385),
.C(n_386),
.Y(n_2476)
);

INVx5_ASAP7_75t_L g2477 ( 
.A(n_2123),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2074),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_SL g2479 ( 
.A(n_2178),
.B(n_387),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2088),
.B(n_389),
.Y(n_2480)
);

BUFx2_ASAP7_75t_L g2481 ( 
.A(n_2033),
.Y(n_2481)
);

INVx4_ASAP7_75t_L g2482 ( 
.A(n_2132),
.Y(n_2482)
);

BUFx6f_ASAP7_75t_L g2483 ( 
.A(n_2212),
.Y(n_2483)
);

NAND3xp33_ASAP7_75t_SL g2484 ( 
.A(n_2453),
.B(n_2031),
.C(n_2012),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2307),
.Y(n_2485)
);

AOI221x1_ASAP7_75t_L g2486 ( 
.A1(n_2253),
.A2(n_2012),
.B1(n_2031),
.B2(n_2148),
.C(n_2145),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2274),
.Y(n_2487)
);

NOR2xp33_ASAP7_75t_L g2488 ( 
.A(n_2363),
.B(n_2190),
.Y(n_2488)
);

AOI21xp5_ASAP7_75t_L g2489 ( 
.A1(n_2271),
.A2(n_2071),
.B(n_1969),
.Y(n_2489)
);

AOI21xp5_ASAP7_75t_L g2490 ( 
.A1(n_2271),
.A2(n_2035),
.B(n_2128),
.Y(n_2490)
);

INVx5_ASAP7_75t_L g2491 ( 
.A(n_2212),
.Y(n_2491)
);

AOI21xp5_ASAP7_75t_L g2492 ( 
.A1(n_2401),
.A2(n_1943),
.B(n_1938),
.Y(n_2492)
);

INVx5_ASAP7_75t_L g2493 ( 
.A(n_2212),
.Y(n_2493)
);

CKINVDCx6p67_ASAP7_75t_R g2494 ( 
.A(n_2240),
.Y(n_2494)
);

OR2x2_ASAP7_75t_SL g2495 ( 
.A(n_2299),
.B(n_2210),
.Y(n_2495)
);

OA21x2_ASAP7_75t_L g2496 ( 
.A1(n_2293),
.A2(n_2198),
.B(n_2145),
.Y(n_2496)
);

INVx1_ASAP7_75t_SL g2497 ( 
.A(n_2395),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2223),
.B(n_2091),
.Y(n_2498)
);

NAND2x1p5_ASAP7_75t_L g2499 ( 
.A(n_2258),
.B(n_2247),
.Y(n_2499)
);

AOI221x1_ASAP7_75t_L g2500 ( 
.A1(n_2253),
.A2(n_2139),
.B1(n_2175),
.B2(n_2184),
.C(n_2194),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2217),
.B(n_2153),
.Y(n_2501)
);

AO32x2_ASAP7_75t_L g2502 ( 
.A1(n_2380),
.A2(n_2139),
.A3(n_2162),
.B1(n_2066),
.B2(n_2194),
.Y(n_2502)
);

BUFx6f_ASAP7_75t_L g2503 ( 
.A(n_2275),
.Y(n_2503)
);

AOI221x1_ASAP7_75t_L g2504 ( 
.A1(n_2386),
.A2(n_2165),
.B1(n_2185),
.B2(n_2063),
.C(n_1959),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2278),
.B(n_2154),
.Y(n_2505)
);

INVx5_ASAP7_75t_L g2506 ( 
.A(n_2275),
.Y(n_2506)
);

AOI21xp5_ASAP7_75t_L g2507 ( 
.A1(n_2335),
.A2(n_2321),
.B(n_2403),
.Y(n_2507)
);

AO21x1_ASAP7_75t_L g2508 ( 
.A1(n_2403),
.A2(n_2009),
.B(n_2102),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2280),
.B(n_2155),
.Y(n_2509)
);

AOI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_2321),
.A2(n_2008),
.B(n_2005),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2333),
.B(n_2161),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2353),
.B(n_1957),
.Y(n_2512)
);

A2O1A1Ixp33_ASAP7_75t_L g2513 ( 
.A1(n_2256),
.A2(n_2018),
.B(n_2047),
.C(n_2041),
.Y(n_2513)
);

AOI22xp5_ASAP7_75t_L g2514 ( 
.A1(n_2309),
.A2(n_2164),
.B1(n_2207),
.B2(n_2090),
.Y(n_2514)
);

OAI21xp5_ASAP7_75t_L g2515 ( 
.A1(n_2440),
.A2(n_2022),
.B(n_2062),
.Y(n_2515)
);

AO31x2_ASAP7_75t_L g2516 ( 
.A1(n_2389),
.A2(n_1947),
.A3(n_2189),
.B(n_2010),
.Y(n_2516)
);

O2A1O1Ixp5_ASAP7_75t_L g2517 ( 
.A1(n_2245),
.A2(n_1971),
.B(n_2084),
.C(n_2143),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2288),
.Y(n_2518)
);

INVx2_ASAP7_75t_SL g2519 ( 
.A(n_2247),
.Y(n_2519)
);

OAI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2309),
.A2(n_1895),
.B1(n_1955),
.B2(n_1962),
.Y(n_2520)
);

AO31x2_ASAP7_75t_L g2521 ( 
.A1(n_2389),
.A2(n_2456),
.A3(n_2218),
.B(n_2220),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2291),
.Y(n_2522)
);

AOI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_2308),
.A2(n_2030),
.B(n_2029),
.Y(n_2523)
);

AOI221x1_ASAP7_75t_L g2524 ( 
.A1(n_2386),
.A2(n_2151),
.B1(n_2150),
.B2(n_2204),
.C(n_2182),
.Y(n_2524)
);

A2O1A1Ixp33_ASAP7_75t_L g2525 ( 
.A1(n_2285),
.A2(n_2191),
.B(n_1949),
.C(n_2195),
.Y(n_2525)
);

A2O1A1Ixp33_ASAP7_75t_L g2526 ( 
.A1(n_2243),
.A2(n_2222),
.B(n_2312),
.C(n_2286),
.Y(n_2526)
);

AOI21xp5_ASAP7_75t_SL g2527 ( 
.A1(n_2343),
.A2(n_2179),
.B(n_2178),
.Y(n_2527)
);

AO22x2_ASAP7_75t_L g2528 ( 
.A1(n_2343),
.A2(n_1958),
.B1(n_2098),
.B2(n_2033),
.Y(n_2528)
);

A2O1A1Ixp33_ASAP7_75t_L g2529 ( 
.A1(n_2405),
.A2(n_2196),
.B(n_2169),
.C(n_2173),
.Y(n_2529)
);

HB1xp67_ASAP7_75t_L g2530 ( 
.A(n_2309),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2323),
.B(n_2206),
.Y(n_2531)
);

AO32x2_ASAP7_75t_L g2532 ( 
.A1(n_2418),
.A2(n_2326),
.A3(n_2319),
.B1(n_2449),
.B2(n_2264),
.Y(n_2532)
);

OAI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2332),
.A2(n_1900),
.B1(n_1989),
.B2(n_1953),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2225),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2248),
.B(n_389),
.Y(n_2535)
);

OAI21xp5_ASAP7_75t_L g2536 ( 
.A1(n_2367),
.A2(n_1892),
.B(n_2174),
.Y(n_2536)
);

AOI21xp5_ASAP7_75t_L g2537 ( 
.A1(n_2375),
.A2(n_2064),
.B(n_2075),
.Y(n_2537)
);

A2O1A1Ixp33_ASAP7_75t_L g2538 ( 
.A1(n_2372),
.A2(n_2157),
.B(n_2188),
.C(n_2172),
.Y(n_2538)
);

OA21x2_ASAP7_75t_L g2539 ( 
.A1(n_2265),
.A2(n_2170),
.B(n_2089),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2314),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2362),
.B(n_1950),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2232),
.Y(n_2542)
);

AOI21xp5_ASAP7_75t_L g2543 ( 
.A1(n_2251),
.A2(n_2097),
.B(n_2081),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_2385),
.B(n_2356),
.Y(n_2544)
);

INVx1_ASAP7_75t_SL g2545 ( 
.A(n_2431),
.Y(n_2545)
);

AOI21xp5_ASAP7_75t_L g2546 ( 
.A1(n_2452),
.A2(n_2146),
.B(n_2152),
.Y(n_2546)
);

AND2x4_ASAP7_75t_L g2547 ( 
.A(n_2361),
.B(n_2420),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2239),
.Y(n_2548)
);

AOI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_2249),
.A2(n_1932),
.B1(n_2201),
.B2(n_1907),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_SL g2550 ( 
.A(n_2238),
.B(n_2086),
.Y(n_2550)
);

INVx6_ASAP7_75t_L g2551 ( 
.A(n_2304),
.Y(n_2551)
);

CKINVDCx6p67_ASAP7_75t_R g2552 ( 
.A(n_2242),
.Y(n_2552)
);

CKINVDCx20_ASAP7_75t_R g2553 ( 
.A(n_2236),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_2382),
.B(n_2086),
.Y(n_2554)
);

OAI21xp5_ASAP7_75t_L g2555 ( 
.A1(n_2297),
.A2(n_2476),
.B(n_2396),
.Y(n_2555)
);

AOI31xp67_ASAP7_75t_L g2556 ( 
.A1(n_2364),
.A2(n_1998),
.A3(n_1999),
.B(n_2176),
.Y(n_2556)
);

AOI21xp5_ASAP7_75t_L g2557 ( 
.A1(n_2466),
.A2(n_2152),
.B(n_1919),
.Y(n_2557)
);

INVxp67_ASAP7_75t_SL g2558 ( 
.A(n_2306),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2379),
.B(n_2387),
.Y(n_2559)
);

A2O1A1Ixp33_ASAP7_75t_L g2560 ( 
.A1(n_2409),
.A2(n_2177),
.B(n_1945),
.C(n_2015),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2241),
.B(n_2098),
.Y(n_2561)
);

OAI21x1_ASAP7_75t_L g2562 ( 
.A1(n_2457),
.A2(n_2112),
.B(n_2055),
.Y(n_2562)
);

OR2x2_ASAP7_75t_L g2563 ( 
.A(n_2273),
.B(n_2125),
.Y(n_2563)
);

INVx5_ASAP7_75t_L g2564 ( 
.A(n_2275),
.Y(n_2564)
);

AOI21xp5_ASAP7_75t_L g2565 ( 
.A1(n_2468),
.A2(n_2034),
.B(n_2038),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2313),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2318),
.Y(n_2567)
);

BUFx6f_ASAP7_75t_L g2568 ( 
.A(n_2279),
.Y(n_2568)
);

AOI221x1_ASAP7_75t_L g2569 ( 
.A1(n_2326),
.A2(n_1956),
.B1(n_2025),
.B2(n_2028),
.C(n_2049),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2374),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2211),
.B(n_2125),
.Y(n_2571)
);

O2A1O1Ixp33_ASAP7_75t_SL g2572 ( 
.A1(n_2339),
.A2(n_1992),
.B(n_1978),
.C(n_1883),
.Y(n_2572)
);

AOI21xp5_ASAP7_75t_L g2573 ( 
.A1(n_2471),
.A2(n_2163),
.B(n_2144),
.Y(n_2573)
);

HB1xp67_ASAP7_75t_L g2574 ( 
.A(n_2246),
.Y(n_2574)
);

BUFx3_ASAP7_75t_L g2575 ( 
.A(n_2295),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_2292),
.Y(n_2576)
);

INVx5_ASAP7_75t_L g2577 ( 
.A(n_2279),
.Y(n_2577)
);

AOI21x1_ASAP7_75t_L g2578 ( 
.A1(n_2472),
.A2(n_2163),
.B(n_2144),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2229),
.B(n_464),
.Y(n_2579)
);

INVx3_ASAP7_75t_L g2580 ( 
.A(n_2252),
.Y(n_2580)
);

AO31x2_ASAP7_75t_L g2581 ( 
.A1(n_2448),
.A2(n_390),
.A3(n_392),
.B(n_393),
.Y(n_2581)
);

AOI21xp5_ASAP7_75t_L g2582 ( 
.A1(n_2478),
.A2(n_390),
.B(n_392),
.Y(n_2582)
);

INVx2_ASAP7_75t_SL g2583 ( 
.A(n_2255),
.Y(n_2583)
);

A2O1A1Ixp33_ASAP7_75t_L g2584 ( 
.A1(n_2270),
.A2(n_393),
.B(n_394),
.C(n_396),
.Y(n_2584)
);

AOI21xp5_ASAP7_75t_L g2585 ( 
.A1(n_2213),
.A2(n_394),
.B(n_396),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2231),
.B(n_463),
.Y(n_2586)
);

AO31x2_ASAP7_75t_L g2587 ( 
.A1(n_2413),
.A2(n_397),
.A3(n_398),
.B(n_400),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2394),
.Y(n_2588)
);

INVxp67_ASAP7_75t_SL g2589 ( 
.A(n_2305),
.Y(n_2589)
);

NAND3xp33_ASAP7_75t_SL g2590 ( 
.A(n_2352),
.B(n_401),
.C(n_402),
.Y(n_2590)
);

AO32x2_ASAP7_75t_L g2591 ( 
.A1(n_2418),
.A2(n_2348),
.A3(n_2317),
.B1(n_2260),
.B2(n_2422),
.Y(n_2591)
);

O2A1O1Ixp33_ASAP7_75t_SL g2592 ( 
.A1(n_2289),
.A2(n_402),
.B(n_404),
.C(n_405),
.Y(n_2592)
);

AOI21xp5_ASAP7_75t_L g2593 ( 
.A1(n_2213),
.A2(n_404),
.B(n_405),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2296),
.B(n_406),
.Y(n_2594)
);

AOI21xp33_ASAP7_75t_L g2595 ( 
.A1(n_2350),
.A2(n_406),
.B(n_407),
.Y(n_2595)
);

AOI21xp5_ASAP7_75t_L g2596 ( 
.A1(n_2391),
.A2(n_407),
.B(n_409),
.Y(n_2596)
);

AO22x2_ASAP7_75t_L g2597 ( 
.A1(n_2385),
.A2(n_410),
.B1(n_411),
.B2(n_413),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2414),
.B(n_463),
.Y(n_2598)
);

AO21x2_ASAP7_75t_L g2599 ( 
.A1(n_2230),
.A2(n_410),
.B(n_411),
.Y(n_2599)
);

OAI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2378),
.A2(n_413),
.B(n_414),
.Y(n_2600)
);

A2O1A1Ixp33_ASAP7_75t_L g2601 ( 
.A1(n_2352),
.A2(n_415),
.B(n_417),
.C(n_418),
.Y(n_2601)
);

O2A1O1Ixp33_ASAP7_75t_L g2602 ( 
.A1(n_2328),
.A2(n_418),
.B(n_419),
.C(n_420),
.Y(n_2602)
);

AOI21xp5_ASAP7_75t_L g2603 ( 
.A1(n_2416),
.A2(n_419),
.B(n_420),
.Y(n_2603)
);

AO21x2_ASAP7_75t_L g2604 ( 
.A1(n_2230),
.A2(n_421),
.B(n_423),
.Y(n_2604)
);

A2O1A1Ixp33_ASAP7_75t_L g2605 ( 
.A1(n_2269),
.A2(n_425),
.B(n_426),
.C(n_427),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2419),
.B(n_462),
.Y(n_2606)
);

OA21x2_ASAP7_75t_L g2607 ( 
.A1(n_2460),
.A2(n_425),
.B(n_428),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2426),
.B(n_428),
.Y(n_2608)
);

AOI21xp5_ASAP7_75t_L g2609 ( 
.A1(n_2427),
.A2(n_429),
.B(n_430),
.Y(n_2609)
);

AND2x4_ASAP7_75t_L g2610 ( 
.A(n_2361),
.B(n_429),
.Y(n_2610)
);

AND2x4_ASAP7_75t_L g2611 ( 
.A(n_2420),
.B(n_430),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2398),
.Y(n_2612)
);

BUFx3_ASAP7_75t_L g2613 ( 
.A(n_2400),
.Y(n_2613)
);

AOI21xp5_ASAP7_75t_L g2614 ( 
.A1(n_2310),
.A2(n_431),
.B(n_432),
.Y(n_2614)
);

AOI21xp5_ASAP7_75t_L g2615 ( 
.A1(n_2310),
.A2(n_2455),
.B(n_2228),
.Y(n_2615)
);

NOR2x1_ASAP7_75t_R g2616 ( 
.A(n_2337),
.B(n_431),
.Y(n_2616)
);

INVx1_ASAP7_75t_SL g2617 ( 
.A(n_2445),
.Y(n_2617)
);

AND2x4_ASAP7_75t_L g2618 ( 
.A(n_2329),
.B(n_2345),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2268),
.B(n_432),
.Y(n_2619)
);

AO31x2_ASAP7_75t_L g2620 ( 
.A1(n_2259),
.A2(n_434),
.A3(n_435),
.B(n_437),
.Y(n_2620)
);

AOI21xp5_ASAP7_75t_L g2621 ( 
.A1(n_2310),
.A2(n_434),
.B(n_438),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2404),
.Y(n_2622)
);

INVx5_ASAP7_75t_L g2623 ( 
.A(n_2279),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2276),
.B(n_440),
.Y(n_2624)
);

INVx3_ASAP7_75t_L g2625 ( 
.A(n_2482),
.Y(n_2625)
);

AOI221x1_ASAP7_75t_L g2626 ( 
.A1(n_2475),
.A2(n_441),
.B1(n_443),
.B2(n_444),
.C(n_445),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2421),
.Y(n_2627)
);

AOI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2399),
.A2(n_444),
.B(n_445),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2347),
.B(n_448),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2226),
.B(n_448),
.Y(n_2630)
);

OA21x2_ASAP7_75t_L g2631 ( 
.A1(n_2462),
.A2(n_449),
.B(n_450),
.Y(n_2631)
);

OAI21x1_ASAP7_75t_L g2632 ( 
.A1(n_2267),
.A2(n_451),
.B(n_452),
.Y(n_2632)
);

AOI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2281),
.A2(n_451),
.B1(n_452),
.B2(n_453),
.Y(n_2633)
);

OA21x2_ASAP7_75t_L g2634 ( 
.A1(n_2311),
.A2(n_2434),
.B(n_2392),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_2262),
.B(n_454),
.Y(n_2635)
);

BUFx6f_ASAP7_75t_L g2636 ( 
.A(n_2454),
.Y(n_2636)
);

BUFx2_ASAP7_75t_L g2637 ( 
.A(n_2303),
.Y(n_2637)
);

AOI221x1_ASAP7_75t_L g2638 ( 
.A1(n_2407),
.A2(n_458),
.B1(n_459),
.B2(n_460),
.C(n_461),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2433),
.Y(n_2639)
);

AND2x4_ASAP7_75t_L g2640 ( 
.A(n_2329),
.B(n_462),
.Y(n_2640)
);

INVx2_ASAP7_75t_SL g2641 ( 
.A(n_2234),
.Y(n_2641)
);

AOI21xp5_ASAP7_75t_L g2642 ( 
.A1(n_2406),
.A2(n_2411),
.B(n_2412),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2219),
.Y(n_2643)
);

OAI21x1_ASAP7_75t_L g2644 ( 
.A1(n_2287),
.A2(n_2233),
.B(n_2215),
.Y(n_2644)
);

NOR2x1_ASAP7_75t_SL g2645 ( 
.A(n_2388),
.B(n_2482),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2227),
.B(n_2298),
.Y(n_2646)
);

AND2x4_ASAP7_75t_L g2647 ( 
.A(n_2345),
.B(n_2355),
.Y(n_2647)
);

AOI21xp5_ASAP7_75t_L g2648 ( 
.A1(n_2469),
.A2(n_2480),
.B(n_2450),
.Y(n_2648)
);

NOR2xp33_ASAP7_75t_L g2649 ( 
.A(n_2351),
.B(n_2316),
.Y(n_2649)
);

CKINVDCx9p33_ASAP7_75t_R g2650 ( 
.A(n_2301),
.Y(n_2650)
);

AOI21xp5_ASAP7_75t_L g2651 ( 
.A1(n_2214),
.A2(n_2216),
.B(n_2467),
.Y(n_2651)
);

OAI21x1_ASAP7_75t_L g2652 ( 
.A1(n_2473),
.A2(n_2479),
.B(n_2434),
.Y(n_2652)
);

AOI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2370),
.A2(n_2334),
.B1(n_2388),
.B2(n_2234),
.Y(n_2653)
);

NOR2xp33_ASAP7_75t_R g2654 ( 
.A(n_2354),
.B(n_2402),
.Y(n_2654)
);

NOR2xp67_ASAP7_75t_SL g2655 ( 
.A(n_2355),
.B(n_2477),
.Y(n_2655)
);

BUFx10_ASAP7_75t_L g2656 ( 
.A(n_2388),
.Y(n_2656)
);

OAI22x1_ASAP7_75t_L g2657 ( 
.A1(n_2357),
.A2(n_2435),
.B1(n_2277),
.B2(n_2221),
.Y(n_2657)
);

NOR2x1_ASAP7_75t_SL g2658 ( 
.A(n_2554),
.B(n_2355),
.Y(n_2658)
);

INVx6_ASAP7_75t_L g2659 ( 
.A(n_2636),
.Y(n_2659)
);

BUFx10_ASAP7_75t_L g2660 ( 
.A(n_2551),
.Y(n_2660)
);

BUFx3_ASAP7_75t_L g2661 ( 
.A(n_2575),
.Y(n_2661)
);

AOI22xp33_ASAP7_75t_L g2662 ( 
.A1(n_2657),
.A2(n_2244),
.B1(n_2484),
.B2(n_2590),
.Y(n_2662)
);

INVxp67_ASAP7_75t_SL g2663 ( 
.A(n_2530),
.Y(n_2663)
);

AOI22xp33_ASAP7_75t_L g2664 ( 
.A1(n_2649),
.A2(n_2244),
.B1(n_2294),
.B2(n_2315),
.Y(n_2664)
);

AOI22xp33_ASAP7_75t_SL g2665 ( 
.A1(n_2645),
.A2(n_2597),
.B1(n_2641),
.B2(n_2656),
.Y(n_2665)
);

CKINVDCx11_ASAP7_75t_R g2666 ( 
.A(n_2553),
.Y(n_2666)
);

BUFx12f_ASAP7_75t_L g2667 ( 
.A(n_2576),
.Y(n_2667)
);

OAI21xp33_ASAP7_75t_L g2668 ( 
.A1(n_2597),
.A2(n_2277),
.B(n_2284),
.Y(n_2668)
);

BUFx3_ASAP7_75t_L g2669 ( 
.A(n_2494),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2544),
.B(n_2302),
.Y(n_2670)
);

AOI22xp33_ASAP7_75t_L g2671 ( 
.A1(n_2594),
.A2(n_2390),
.B1(n_2237),
.B2(n_2368),
.Y(n_2671)
);

AOI22xp5_ASAP7_75t_L g2672 ( 
.A1(n_2653),
.A2(n_2290),
.B1(n_2327),
.B2(n_2465),
.Y(n_2672)
);

AOI22xp5_ASAP7_75t_L g2673 ( 
.A1(n_2646),
.A2(n_2501),
.B1(n_2633),
.B2(n_2600),
.Y(n_2673)
);

AOI22xp33_ASAP7_75t_L g2674 ( 
.A1(n_2515),
.A2(n_2425),
.B1(n_2300),
.B2(n_2357),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_L g2675 ( 
.A1(n_2512),
.A2(n_2425),
.B1(n_2435),
.B2(n_2441),
.Y(n_2675)
);

INVxp67_ASAP7_75t_SL g2676 ( 
.A(n_2574),
.Y(n_2676)
);

OR2x2_ASAP7_75t_L g2677 ( 
.A(n_2540),
.B(n_2376),
.Y(n_2677)
);

BUFx8_ASAP7_75t_L g2678 ( 
.A(n_2613),
.Y(n_2678)
);

INVx6_ASAP7_75t_L g2679 ( 
.A(n_2636),
.Y(n_2679)
);

INVx1_ASAP7_75t_SL g2680 ( 
.A(n_2637),
.Y(n_2680)
);

INVx4_ASAP7_75t_SL g2681 ( 
.A(n_2551),
.Y(n_2681)
);

HB1xp67_ASAP7_75t_L g2682 ( 
.A(n_2589),
.Y(n_2682)
);

OR2x2_ASAP7_75t_L g2683 ( 
.A(n_2542),
.B(n_2283),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2559),
.B(n_2474),
.Y(n_2684)
);

BUFx3_ASAP7_75t_L g2685 ( 
.A(n_2552),
.Y(n_2685)
);

NAND2x1p5_ASAP7_75t_L g2686 ( 
.A(n_2655),
.B(n_2477),
.Y(n_2686)
);

NAND2x1p5_ASAP7_75t_L g2687 ( 
.A(n_2491),
.B(n_2477),
.Y(n_2687)
);

BUFx2_ASAP7_75t_L g2688 ( 
.A(n_2625),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2485),
.Y(n_2689)
);

AOI22xp33_ASAP7_75t_SL g2690 ( 
.A1(n_2610),
.A2(n_2266),
.B1(n_2392),
.B2(n_2428),
.Y(n_2690)
);

AOI22xp33_ASAP7_75t_SL g2691 ( 
.A1(n_2610),
.A2(n_2266),
.B1(n_2470),
.B2(n_2366),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2487),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2518),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2522),
.B(n_2410),
.Y(n_2694)
);

CKINVDCx20_ASAP7_75t_R g2695 ( 
.A(n_2654),
.Y(n_2695)
);

AOI22xp33_ASAP7_75t_L g2696 ( 
.A1(n_2640),
.A2(n_2535),
.B1(n_2520),
.B2(n_2595),
.Y(n_2696)
);

AOI22xp33_ASAP7_75t_L g2697 ( 
.A1(n_2640),
.A2(n_2438),
.B1(n_2424),
.B2(n_2263),
.Y(n_2697)
);

INVx1_ASAP7_75t_SL g2698 ( 
.A(n_2637),
.Y(n_2698)
);

BUFx12f_ASAP7_75t_L g2699 ( 
.A(n_2499),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2548),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2566),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2567),
.Y(n_2702)
);

BUFx3_ASAP7_75t_L g2703 ( 
.A(n_2617),
.Y(n_2703)
);

CKINVDCx20_ASAP7_75t_R g2704 ( 
.A(n_2497),
.Y(n_2704)
);

INVx3_ASAP7_75t_SL g2705 ( 
.A(n_2545),
.Y(n_2705)
);

BUFx8_ASAP7_75t_L g2706 ( 
.A(n_2583),
.Y(n_2706)
);

INVx6_ASAP7_75t_L g2707 ( 
.A(n_2491),
.Y(n_2707)
);

OAI22xp5_ASAP7_75t_L g2708 ( 
.A1(n_2601),
.A2(n_2272),
.B1(n_2444),
.B2(n_2224),
.Y(n_2708)
);

INVx3_ASAP7_75t_L g2709 ( 
.A(n_2491),
.Y(n_2709)
);

BUFx6f_ASAP7_75t_L g2710 ( 
.A(n_2493),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2570),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2498),
.B(n_2340),
.Y(n_2712)
);

INVx4_ASAP7_75t_L g2713 ( 
.A(n_2493),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2588),
.Y(n_2714)
);

OAI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2514),
.A2(n_2495),
.B1(n_2584),
.B2(n_2605),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2612),
.B(n_2235),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2627),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2639),
.Y(n_2718)
);

BUFx2_ASAP7_75t_L g2719 ( 
.A(n_2483),
.Y(n_2719)
);

AOI22xp33_ASAP7_75t_SL g2720 ( 
.A1(n_2611),
.A2(n_2470),
.B1(n_2481),
.B2(n_2451),
.Y(n_2720)
);

OAI22xp5_ASAP7_75t_L g2721 ( 
.A1(n_2611),
.A2(n_2393),
.B1(n_2397),
.B2(n_2282),
.Y(n_2721)
);

INVx6_ASAP7_75t_L g2722 ( 
.A(n_2493),
.Y(n_2722)
);

AOI22xp33_ASAP7_75t_SL g2723 ( 
.A1(n_2550),
.A2(n_2436),
.B1(n_2383),
.B2(n_2408),
.Y(n_2723)
);

OAI22xp5_ASAP7_75t_L g2724 ( 
.A1(n_2526),
.A2(n_2558),
.B1(n_2507),
.B2(n_2513),
.Y(n_2724)
);

BUFx10_ASAP7_75t_L g2725 ( 
.A(n_2547),
.Y(n_2725)
);

OAI22xp5_ASAP7_75t_SL g2726 ( 
.A1(n_2616),
.A2(n_2250),
.B1(n_2257),
.B2(n_2261),
.Y(n_2726)
);

AOI22xp33_ASAP7_75t_L g2727 ( 
.A1(n_2643),
.A2(n_2359),
.B1(n_2459),
.B2(n_2458),
.Y(n_2727)
);

AOI22xp5_ASAP7_75t_L g2728 ( 
.A1(n_2541),
.A2(n_2464),
.B1(n_2341),
.B2(n_2439),
.Y(n_2728)
);

AOI22xp33_ASAP7_75t_L g2729 ( 
.A1(n_2508),
.A2(n_2430),
.B1(n_2443),
.B2(n_2429),
.Y(n_2729)
);

OAI22xp5_ASAP7_75t_L g2730 ( 
.A1(n_2549),
.A2(n_2331),
.B1(n_2417),
.B2(n_2325),
.Y(n_2730)
);

INVx6_ASAP7_75t_L g2731 ( 
.A(n_2506),
.Y(n_2731)
);

OAI22xp5_ASAP7_75t_L g2732 ( 
.A1(n_2571),
.A2(n_2320),
.B1(n_2338),
.B2(n_2322),
.Y(n_2732)
);

INVx6_ASAP7_75t_L g2733 ( 
.A(n_2506),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_2650),
.Y(n_2734)
);

CKINVDCx5p33_ASAP7_75t_R g2735 ( 
.A(n_2506),
.Y(n_2735)
);

BUFx8_ASAP7_75t_SL g2736 ( 
.A(n_2534),
.Y(n_2736)
);

OAI22xp5_ASAP7_75t_L g2737 ( 
.A1(n_2580),
.A2(n_2423),
.B1(n_2437),
.B2(n_2447),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2622),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2563),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2511),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2561),
.Y(n_2741)
);

AOI22xp33_ASAP7_75t_SL g2742 ( 
.A1(n_2533),
.A2(n_2383),
.B1(n_2377),
.B2(n_2446),
.Y(n_2742)
);

INVx1_ASAP7_75t_SL g2743 ( 
.A(n_2483),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2505),
.B(n_2330),
.Y(n_2744)
);

AOI22xp33_ASAP7_75t_SL g2745 ( 
.A1(n_2528),
.A2(n_2383),
.B1(n_2377),
.B2(n_2303),
.Y(n_2745)
);

CKINVDCx6p67_ASAP7_75t_R g2746 ( 
.A(n_2564),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_SL g2747 ( 
.A1(n_2528),
.A2(n_2463),
.B1(n_2360),
.B2(n_2303),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2509),
.B(n_2324),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2531),
.Y(n_2749)
);

AOI22xp33_ASAP7_75t_L g2750 ( 
.A1(n_2642),
.A2(n_2369),
.B1(n_2365),
.B2(n_2336),
.Y(n_2750)
);

OAI22xp33_ASAP7_75t_L g2751 ( 
.A1(n_2486),
.A2(n_2349),
.B1(n_2342),
.B2(n_2373),
.Y(n_2751)
);

AOI22xp33_ASAP7_75t_L g2752 ( 
.A1(n_2648),
.A2(n_2384),
.B1(n_2344),
.B2(n_2346),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2598),
.Y(n_2753)
);

OAI22xp5_ASAP7_75t_L g2754 ( 
.A1(n_2492),
.A2(n_2381),
.B1(n_2254),
.B2(n_2415),
.Y(n_2754)
);

CKINVDCx11_ASAP7_75t_R g2755 ( 
.A(n_2503),
.Y(n_2755)
);

CKINVDCx11_ASAP7_75t_R g2756 ( 
.A(n_2503),
.Y(n_2756)
);

AOI22xp5_ASAP7_75t_SL g2757 ( 
.A1(n_2547),
.A2(n_2461),
.B1(n_2358),
.B2(n_2360),
.Y(n_2757)
);

INVx4_ASAP7_75t_L g2758 ( 
.A(n_2564),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2606),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2608),
.Y(n_2760)
);

CKINVDCx11_ASAP7_75t_R g2761 ( 
.A(n_2568),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2587),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2618),
.B(n_2371),
.Y(n_2763)
);

BUFx12f_ASAP7_75t_L g2764 ( 
.A(n_2564),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2568),
.Y(n_2765)
);

INVx5_ASAP7_75t_L g2766 ( 
.A(n_2577),
.Y(n_2766)
);

AOI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2579),
.A2(n_2358),
.B1(n_2432),
.B2(n_2442),
.Y(n_2767)
);

AOI22xp33_ASAP7_75t_L g2768 ( 
.A1(n_2628),
.A2(n_2432),
.B1(n_2442),
.B2(n_2463),
.Y(n_2768)
);

OAI21xp5_ASAP7_75t_SL g2769 ( 
.A1(n_2500),
.A2(n_2602),
.B(n_2489),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2582),
.A2(n_2371),
.B1(n_2635),
.B2(n_2630),
.Y(n_2770)
);

INVx8_ASAP7_75t_L g2771 ( 
.A(n_2577),
.Y(n_2771)
);

OAI22xp5_ASAP7_75t_L g2772 ( 
.A1(n_2651),
.A2(n_2371),
.B1(n_2586),
.B2(n_2619),
.Y(n_2772)
);

BUFx6f_ASAP7_75t_L g2773 ( 
.A(n_2577),
.Y(n_2773)
);

BUFx3_ASAP7_75t_L g2774 ( 
.A(n_2623),
.Y(n_2774)
);

BUFx8_ASAP7_75t_L g2775 ( 
.A(n_2519),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2623),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2618),
.B(n_2624),
.Y(n_2777)
);

AOI22x1_ASAP7_75t_SL g2778 ( 
.A1(n_2532),
.A2(n_2591),
.B1(n_2623),
.B2(n_2638),
.Y(n_2778)
);

BUFx3_ASAP7_75t_L g2779 ( 
.A(n_2647),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2488),
.B(n_2647),
.Y(n_2780)
);

AOI22xp33_ASAP7_75t_L g2781 ( 
.A1(n_2596),
.A2(n_2603),
.B1(n_2609),
.B2(n_2555),
.Y(n_2781)
);

HB1xp67_ASAP7_75t_L g2782 ( 
.A(n_2682),
.Y(n_2782)
);

BUFx2_ASAP7_75t_L g2783 ( 
.A(n_2680),
.Y(n_2783)
);

AO21x1_ASAP7_75t_L g2784 ( 
.A1(n_2724),
.A2(n_2614),
.B(n_2621),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2762),
.Y(n_2785)
);

INVx2_ASAP7_75t_SL g2786 ( 
.A(n_2771),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2749),
.B(n_2521),
.Y(n_2787)
);

AO21x2_ASAP7_75t_L g2788 ( 
.A1(n_2769),
.A2(n_2615),
.B(n_2536),
.Y(n_2788)
);

INVxp33_ASAP7_75t_L g2789 ( 
.A(n_2736),
.Y(n_2789)
);

INVxp67_ASAP7_75t_L g2790 ( 
.A(n_2688),
.Y(n_2790)
);

AOI22xp33_ASAP7_75t_SL g2791 ( 
.A1(n_2778),
.A2(n_2634),
.B1(n_2607),
.B2(n_2631),
.Y(n_2791)
);

HB1xp67_ASAP7_75t_L g2792 ( 
.A(n_2676),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2740),
.B(n_2629),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2689),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2692),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2693),
.B(n_2521),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2739),
.B(n_2581),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2701),
.B(n_2581),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2700),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2702),
.Y(n_2800)
);

AO21x2_ASAP7_75t_L g2801 ( 
.A1(n_2769),
.A2(n_2557),
.B(n_2510),
.Y(n_2801)
);

BUFx4f_ASAP7_75t_SL g2802 ( 
.A(n_2695),
.Y(n_2802)
);

O2A1O1Ixp5_ASAP7_75t_L g2803 ( 
.A1(n_2713),
.A2(n_2585),
.B(n_2593),
.C(n_2578),
.Y(n_2803)
);

AO21x2_ASAP7_75t_L g2804 ( 
.A1(n_2772),
.A2(n_2490),
.B(n_2604),
.Y(n_2804)
);

OR2x6_ASAP7_75t_L g2805 ( 
.A(n_2771),
.B(n_2527),
.Y(n_2805)
);

HB1xp67_ASAP7_75t_L g2806 ( 
.A(n_2680),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2711),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2714),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2717),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2718),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2763),
.B(n_2634),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2738),
.Y(n_2812)
);

AO21x1_ASAP7_75t_SL g2813 ( 
.A1(n_2767),
.A2(n_2556),
.B(n_2532),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2741),
.B(n_2620),
.Y(n_2814)
);

INVxp67_ASAP7_75t_L g2815 ( 
.A(n_2706),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2698),
.Y(n_2816)
);

BUFx2_ASAP7_75t_L g2817 ( 
.A(n_2698),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2716),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2765),
.Y(n_2819)
);

INVx3_ASAP7_75t_L g2820 ( 
.A(n_2713),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2663),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2753),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2759),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2760),
.Y(n_2824)
);

HB1xp67_ASAP7_75t_L g2825 ( 
.A(n_2677),
.Y(n_2825)
);

INVx2_ASAP7_75t_SL g2826 ( 
.A(n_2771),
.Y(n_2826)
);

OAI21x1_ASAP7_75t_L g2827 ( 
.A1(n_2768),
.A2(n_2546),
.B(n_2523),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2757),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2757),
.Y(n_2829)
);

INVx3_ASAP7_75t_L g2830 ( 
.A(n_2758),
.Y(n_2830)
);

INVx2_ASAP7_75t_SL g2831 ( 
.A(n_2766),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2694),
.Y(n_2832)
);

AND2x4_ASAP7_75t_L g2833 ( 
.A(n_2779),
.B(n_2644),
.Y(n_2833)
);

AOI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2754),
.A2(n_2572),
.B(n_2543),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2683),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2719),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2743),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2747),
.Y(n_2838)
);

INVx2_ASAP7_75t_SL g2839 ( 
.A(n_2766),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2744),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2670),
.B(n_2516),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2748),
.Y(n_2842)
);

INVx3_ASAP7_75t_L g2843 ( 
.A(n_2758),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2780),
.B(n_2516),
.Y(n_2844)
);

AOI21xp5_ASAP7_75t_L g2845 ( 
.A1(n_2754),
.A2(n_2537),
.B(n_2496),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2662),
.B(n_2607),
.Y(n_2846)
);

AOI22xp33_ASAP7_75t_L g2847 ( 
.A1(n_2668),
.A2(n_2631),
.B1(n_2599),
.B2(n_2573),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2684),
.B(n_2712),
.Y(n_2848)
);

BUFx6f_ASAP7_75t_L g2849 ( 
.A(n_2710),
.Y(n_2849)
);

INVx5_ASAP7_75t_SL g2850 ( 
.A(n_2746),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2745),
.Y(n_2851)
);

AOI21x1_ASAP7_75t_L g2852 ( 
.A1(n_2730),
.A2(n_2539),
.B(n_2496),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2777),
.B(n_2532),
.Y(n_2853)
);

INVx5_ASAP7_75t_L g2854 ( 
.A(n_2710),
.Y(n_2854)
);

BUFx2_ASAP7_75t_L g2855 ( 
.A(n_2820),
.Y(n_2855)
);

OR2x2_ASAP7_75t_L g2856 ( 
.A(n_2782),
.B(n_2703),
.Y(n_2856)
);

OAI21xp5_ASAP7_75t_L g2857 ( 
.A1(n_2846),
.A2(n_2665),
.B(n_2715),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2794),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2844),
.B(n_2770),
.Y(n_2859)
);

AND2x2_ASAP7_75t_L g2860 ( 
.A(n_2844),
.B(n_2841),
.Y(n_2860)
);

OAI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2846),
.A2(n_2668),
.B(n_2691),
.Y(n_2861)
);

AND2x2_ASAP7_75t_L g2862 ( 
.A(n_2841),
.B(n_2696),
.Y(n_2862)
);

NOR2x1_ASAP7_75t_SL g2863 ( 
.A(n_2805),
.B(n_2764),
.Y(n_2863)
);

AND2x6_ASAP7_75t_L g2864 ( 
.A(n_2828),
.B(n_2710),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2785),
.Y(n_2865)
);

A2O1A1Ixp33_ASAP7_75t_L g2866 ( 
.A1(n_2786),
.A2(n_2664),
.B(n_2720),
.C(n_2674),
.Y(n_2866)
);

OR2x2_ASAP7_75t_L g2867 ( 
.A(n_2792),
.B(n_2705),
.Y(n_2867)
);

AO32x2_ASAP7_75t_L g2868 ( 
.A1(n_2831),
.A2(n_2732),
.A3(n_2737),
.B1(n_2726),
.B2(n_2721),
.Y(n_2868)
);

AND2x4_ASAP7_75t_L g2869 ( 
.A(n_2833),
.B(n_2766),
.Y(n_2869)
);

INVx1_ASAP7_75t_SL g2870 ( 
.A(n_2802),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2811),
.B(n_2620),
.Y(n_2871)
);

AND2x2_ASAP7_75t_L g2872 ( 
.A(n_2811),
.B(n_2620),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2785),
.Y(n_2873)
);

OR2x2_ASAP7_75t_L g2874 ( 
.A(n_2835),
.B(n_2661),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2796),
.B(n_2781),
.Y(n_2875)
);

OR2x6_ASAP7_75t_L g2876 ( 
.A(n_2805),
.B(n_2828),
.Y(n_2876)
);

INVxp67_ASAP7_75t_L g2877 ( 
.A(n_2832),
.Y(n_2877)
);

NAND3xp33_ASAP7_75t_L g2878 ( 
.A(n_2851),
.B(n_2706),
.C(n_2690),
.Y(n_2878)
);

AND2x4_ASAP7_75t_L g2879 ( 
.A(n_2833),
.B(n_2709),
.Y(n_2879)
);

AOI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2832),
.A2(n_2726),
.B1(n_2673),
.B2(n_2671),
.Y(n_2880)
);

A2O1A1Ixp33_ASAP7_75t_L g2881 ( 
.A1(n_2786),
.A2(n_2675),
.B(n_2673),
.C(n_2742),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2794),
.Y(n_2882)
);

OR2x2_ASAP7_75t_L g2883 ( 
.A(n_2835),
.B(n_2743),
.Y(n_2883)
);

NAND2xp33_ASAP7_75t_L g2884 ( 
.A(n_2826),
.B(n_2734),
.Y(n_2884)
);

AND2x2_ASAP7_75t_L g2885 ( 
.A(n_2796),
.B(n_2652),
.Y(n_2885)
);

AND2x2_ASAP7_75t_L g2886 ( 
.A(n_2825),
.B(n_2776),
.Y(n_2886)
);

AOI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2853),
.A2(n_2708),
.B1(n_2672),
.B2(n_2728),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2853),
.B(n_2728),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2787),
.B(n_2502),
.Y(n_2889)
);

AOI22xp33_ASAP7_75t_L g2890 ( 
.A1(n_2840),
.A2(n_2672),
.B1(n_2727),
.B2(n_2697),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2836),
.B(n_2709),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2836),
.B(n_2840),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2842),
.B(n_2790),
.Y(n_2893)
);

INVxp67_ASAP7_75t_L g2894 ( 
.A(n_2842),
.Y(n_2894)
);

AND2x2_ASAP7_75t_L g2895 ( 
.A(n_2787),
.B(n_2788),
.Y(n_2895)
);

INVx5_ASAP7_75t_SL g2896 ( 
.A(n_2805),
.Y(n_2896)
);

OR2x2_ASAP7_75t_L g2897 ( 
.A(n_2821),
.B(n_2774),
.Y(n_2897)
);

AND2x2_ASAP7_75t_L g2898 ( 
.A(n_2788),
.B(n_2502),
.Y(n_2898)
);

AND2x2_ASAP7_75t_L g2899 ( 
.A(n_2788),
.B(n_2502),
.Y(n_2899)
);

OR2x6_ASAP7_75t_L g2900 ( 
.A(n_2805),
.B(n_2686),
.Y(n_2900)
);

OAI21xp5_ASAP7_75t_L g2901 ( 
.A1(n_2834),
.A2(n_2729),
.B(n_2626),
.Y(n_2901)
);

OAI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2851),
.A2(n_2517),
.B(n_2723),
.Y(n_2902)
);

INVxp67_ASAP7_75t_L g2903 ( 
.A(n_2806),
.Y(n_2903)
);

OR2x6_ASAP7_75t_L g2904 ( 
.A(n_2876),
.B(n_2829),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2865),
.Y(n_2905)
);

AND2x2_ASAP7_75t_L g2906 ( 
.A(n_2860),
.B(n_2801),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2858),
.Y(n_2907)
);

HB1xp67_ASAP7_75t_L g2908 ( 
.A(n_2903),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2882),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2889),
.B(n_2823),
.Y(n_2910)
);

INVxp67_ASAP7_75t_SL g2911 ( 
.A(n_2867),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2865),
.Y(n_2912)
);

BUFx3_ASAP7_75t_L g2913 ( 
.A(n_2855),
.Y(n_2913)
);

NOR2xp33_ASAP7_75t_L g2914 ( 
.A(n_2870),
.B(n_2815),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2873),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_R g2916 ( 
.A(n_2884),
.B(n_2666),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2860),
.B(n_2801),
.Y(n_2917)
);

BUFx2_ASAP7_75t_L g2918 ( 
.A(n_2869),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2873),
.Y(n_2919)
);

INVxp67_ASAP7_75t_SL g2920 ( 
.A(n_2856),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2892),
.Y(n_2921)
);

NOR2xp67_ASAP7_75t_L g2922 ( 
.A(n_2878),
.B(n_2820),
.Y(n_2922)
);

AND2x2_ASAP7_75t_L g2923 ( 
.A(n_2895),
.B(n_2801),
.Y(n_2923)
);

AND2x2_ASAP7_75t_L g2924 ( 
.A(n_2895),
.B(n_2885),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2885),
.B(n_2804),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2875),
.B(n_2804),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2894),
.Y(n_2927)
);

HB1xp67_ASAP7_75t_L g2928 ( 
.A(n_2874),
.Y(n_2928)
);

INVx2_ASAP7_75t_SL g2929 ( 
.A(n_2869),
.Y(n_2929)
);

INVx1_ASAP7_75t_SL g2930 ( 
.A(n_2897),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2871),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2877),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2883),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2889),
.B(n_2823),
.Y(n_2934)
);

INVx1_ASAP7_75t_SL g2935 ( 
.A(n_2886),
.Y(n_2935)
);

NOR2xp33_ASAP7_75t_L g2936 ( 
.A(n_2893),
.B(n_2789),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2875),
.Y(n_2937)
);

AOI21xp5_ASAP7_75t_SL g2938 ( 
.A1(n_2863),
.A2(n_2826),
.B(n_2831),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2888),
.B(n_2824),
.Y(n_2939)
);

AOI22xp33_ASAP7_75t_L g2940 ( 
.A1(n_2890),
.A2(n_2818),
.B1(n_2848),
.B2(n_2838),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2871),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2872),
.B(n_2804),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2905),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2924),
.B(n_2859),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2924),
.B(n_2906),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2924),
.B(n_2859),
.Y(n_2946)
);

NOR3xp33_ASAP7_75t_L g2947 ( 
.A(n_2914),
.B(n_2866),
.C(n_2881),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2906),
.B(n_2862),
.Y(n_2948)
);

AOI221xp5_ASAP7_75t_L g2949 ( 
.A1(n_2926),
.A2(n_2866),
.B1(n_2890),
.B2(n_2857),
.C(n_2881),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2905),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2905),
.Y(n_2951)
);

AOI221xp5_ASAP7_75t_L g2952 ( 
.A1(n_2926),
.A2(n_2861),
.B1(n_2887),
.B2(n_2880),
.C(n_2862),
.Y(n_2952)
);

AO21x2_ASAP7_75t_L g2953 ( 
.A1(n_2926),
.A2(n_2845),
.B(n_2901),
.Y(n_2953)
);

AOI22xp33_ASAP7_75t_L g2954 ( 
.A1(n_2937),
.A2(n_2838),
.B1(n_2876),
.B2(n_2829),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2919),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2919),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2912),
.Y(n_2957)
);

OR2x2_ASAP7_75t_L g2958 ( 
.A(n_2937),
.B(n_2872),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2942),
.B(n_2898),
.Y(n_2959)
);

OR2x2_ASAP7_75t_L g2960 ( 
.A(n_2931),
.B(n_2821),
.Y(n_2960)
);

OR2x2_ASAP7_75t_L g2961 ( 
.A(n_2931),
.B(n_2783),
.Y(n_2961)
);

AOI22xp33_ASAP7_75t_L g2962 ( 
.A1(n_2940),
.A2(n_2876),
.B1(n_2902),
.B2(n_2899),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2912),
.Y(n_2963)
);

INVx3_ASAP7_75t_SL g2964 ( 
.A(n_2904),
.Y(n_2964)
);

AO21x2_ASAP7_75t_L g2965 ( 
.A1(n_2923),
.A2(n_2899),
.B(n_2898),
.Y(n_2965)
);

NOR2xp33_ASAP7_75t_L g2966 ( 
.A(n_2936),
.B(n_2685),
.Y(n_2966)
);

NAND2x1p5_ASAP7_75t_L g2967 ( 
.A(n_2913),
.B(n_2820),
.Y(n_2967)
);

AOI33xp33_ASAP7_75t_L g2968 ( 
.A1(n_2940),
.A2(n_2818),
.A3(n_2822),
.B1(n_2791),
.B2(n_2824),
.B3(n_2809),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2912),
.Y(n_2969)
);

OAI21xp5_ASAP7_75t_L g2970 ( 
.A1(n_2938),
.A2(n_2922),
.B(n_2884),
.Y(n_2970)
);

AND2x4_ASAP7_75t_SL g2971 ( 
.A(n_2928),
.B(n_2900),
.Y(n_2971)
);

AO21x2_ASAP7_75t_L g2972 ( 
.A1(n_2923),
.A2(n_2852),
.B(n_2827),
.Y(n_2972)
);

AND2x4_ASAP7_75t_L g2973 ( 
.A(n_2904),
.B(n_2879),
.Y(n_2973)
);

AND2x2_ASAP7_75t_L g2974 ( 
.A(n_2906),
.B(n_2891),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2915),
.Y(n_2975)
);

BUFx2_ASAP7_75t_L g2976 ( 
.A(n_2913),
.Y(n_2976)
);

OAI22xp5_ASAP7_75t_SL g2977 ( 
.A1(n_2916),
.A2(n_2704),
.B1(n_2900),
.B2(n_2669),
.Y(n_2977)
);

AND2x4_ASAP7_75t_L g2978 ( 
.A(n_2904),
.B(n_2879),
.Y(n_2978)
);

HB1xp67_ASAP7_75t_L g2979 ( 
.A(n_2928),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2917),
.B(n_2783),
.Y(n_2980)
);

AOI22xp33_ASAP7_75t_L g2981 ( 
.A1(n_2917),
.A2(n_2864),
.B1(n_2813),
.B2(n_2900),
.Y(n_2981)
);

AOI33xp33_ASAP7_75t_L g2982 ( 
.A1(n_2923),
.A2(n_2822),
.A3(n_2795),
.B1(n_2799),
.B2(n_2808),
.B3(n_2810),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2945),
.B(n_2917),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2952),
.B(n_2925),
.Y(n_2984)
);

AND2x4_ASAP7_75t_L g2985 ( 
.A(n_2973),
.B(n_2904),
.Y(n_2985)
);

OR2x2_ASAP7_75t_L g2986 ( 
.A(n_2959),
.B(n_2910),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2960),
.Y(n_2987)
);

OR2x2_ASAP7_75t_L g2988 ( 
.A(n_2959),
.B(n_2960),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2955),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2945),
.B(n_2925),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2955),
.Y(n_2991)
);

HB1xp67_ASAP7_75t_L g2992 ( 
.A(n_2979),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_SL g2993 ( 
.A(n_2970),
.B(n_2922),
.Y(n_2993)
);

AND2x2_ASAP7_75t_L g2994 ( 
.A(n_2944),
.B(n_2925),
.Y(n_2994)
);

OR2x2_ASAP7_75t_L g2995 ( 
.A(n_2979),
.B(n_2965),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2943),
.Y(n_2996)
);

NAND5xp2_ASAP7_75t_L g2997 ( 
.A(n_2949),
.B(n_2847),
.C(n_2868),
.D(n_2911),
.E(n_2750),
.Y(n_2997)
);

OR2x2_ASAP7_75t_L g2998 ( 
.A(n_2965),
.B(n_2910),
.Y(n_2998)
);

AND2x2_ASAP7_75t_L g2999 ( 
.A(n_2944),
.B(n_2946),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2952),
.B(n_2942),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2943),
.Y(n_3001)
);

BUFx2_ASAP7_75t_L g3002 ( 
.A(n_2970),
.Y(n_3002)
);

INVx3_ASAP7_75t_L g3003 ( 
.A(n_2967),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2956),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_3000),
.B(n_2949),
.Y(n_3005)
);

AND2x2_ASAP7_75t_L g3006 ( 
.A(n_2999),
.B(n_2946),
.Y(n_3006)
);

AOI322xp5_ASAP7_75t_L g3007 ( 
.A1(n_2984),
.A2(n_2947),
.A3(n_2962),
.B1(n_2948),
.B2(n_2911),
.C1(n_2954),
.C2(n_2973),
.Y(n_3007)
);

INVx1_ASAP7_75t_SL g3008 ( 
.A(n_3002),
.Y(n_3008)
);

OR2x2_ASAP7_75t_L g3009 ( 
.A(n_2998),
.B(n_2965),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2999),
.B(n_2968),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2996),
.Y(n_3011)
);

AND2x2_ASAP7_75t_L g3012 ( 
.A(n_3002),
.B(n_2965),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2989),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2989),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2987),
.B(n_2982),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2987),
.B(n_2948),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2992),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2996),
.Y(n_3018)
);

AOI211xp5_ASAP7_75t_L g3019 ( 
.A1(n_2997),
.A2(n_2977),
.B(n_2947),
.C(n_2964),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2991),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_SL g3021 ( 
.A(n_3003),
.B(n_2977),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2994),
.B(n_2964),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2991),
.Y(n_3023)
);

OR2x2_ASAP7_75t_L g3024 ( 
.A(n_2998),
.B(n_2988),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_3004),
.Y(n_3025)
);

AND2x2_ASAP7_75t_L g3026 ( 
.A(n_2994),
.B(n_2964),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2996),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_3004),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_3005),
.B(n_2988),
.Y(n_3029)
);

OR2x2_ASAP7_75t_L g3030 ( 
.A(n_3024),
.B(n_2986),
.Y(n_3030)
);

AND2x4_ASAP7_75t_SL g3031 ( 
.A(n_3017),
.B(n_2660),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_3006),
.B(n_2985),
.Y(n_3032)
);

OR2x2_ASAP7_75t_L g3033 ( 
.A(n_3024),
.B(n_2986),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_3008),
.B(n_2995),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_3015),
.B(n_3001),
.Y(n_3035)
);

NOR2xp67_ASAP7_75t_L g3036 ( 
.A(n_3009),
.B(n_2993),
.Y(n_3036)
);

AND2x2_ASAP7_75t_L g3037 ( 
.A(n_3006),
.B(n_2985),
.Y(n_3037)
);

AND2x2_ASAP7_75t_L g3038 ( 
.A(n_3022),
.B(n_2985),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_3013),
.Y(n_3039)
);

OR2x2_ASAP7_75t_L g3040 ( 
.A(n_3016),
.B(n_2995),
.Y(n_3040)
);

OAI21xp5_ASAP7_75t_L g3041 ( 
.A1(n_3019),
.A2(n_3003),
.B(n_2976),
.Y(n_3041)
);

OR2x2_ASAP7_75t_L g3042 ( 
.A(n_3010),
.B(n_3009),
.Y(n_3042)
);

AND2x4_ASAP7_75t_L g3043 ( 
.A(n_3022),
.B(n_2985),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_3021),
.B(n_2983),
.Y(n_3044)
);

AND2x2_ASAP7_75t_L g3045 ( 
.A(n_3026),
.B(n_2983),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_3026),
.B(n_2990),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_3029),
.B(n_3007),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_3032),
.B(n_3012),
.Y(n_3048)
);

INVx1_ASAP7_75t_SL g3049 ( 
.A(n_3031),
.Y(n_3049)
);

AOI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_3029),
.A2(n_3012),
.B1(n_3003),
.B2(n_2953),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_3036),
.B(n_3023),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_3030),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_3037),
.B(n_2990),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_3045),
.B(n_3046),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_3033),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_3034),
.Y(n_3056)
);

AND2x2_ASAP7_75t_L g3057 ( 
.A(n_3038),
.B(n_3041),
.Y(n_3057)
);

OR2x2_ASAP7_75t_L g3058 ( 
.A(n_3042),
.B(n_3025),
.Y(n_3058)
);

O2A1O1Ixp33_ASAP7_75t_L g3059 ( 
.A1(n_3041),
.A2(n_3003),
.B(n_2976),
.C(n_2908),
.Y(n_3059)
);

NOR4xp25_ASAP7_75t_L g3060 ( 
.A(n_3035),
.B(n_3028),
.C(n_3013),
.D(n_3020),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_3039),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_3038),
.B(n_3014),
.Y(n_3062)
);

OAI322xp33_ASAP7_75t_L g3063 ( 
.A1(n_3047),
.A2(n_3035),
.A3(n_3040),
.B1(n_3044),
.B2(n_2966),
.C1(n_3014),
.C2(n_3028),
.Y(n_3063)
);

AND2x2_ASAP7_75t_L g3064 ( 
.A(n_3054),
.B(n_3043),
.Y(n_3064)
);

OAI21xp5_ASAP7_75t_L g3065 ( 
.A1(n_3049),
.A2(n_3056),
.B(n_3059),
.Y(n_3065)
);

AOI321xp33_ASAP7_75t_L g3066 ( 
.A1(n_3057),
.A2(n_3043),
.A3(n_2920),
.B1(n_2981),
.B2(n_2868),
.C(n_3020),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_3054),
.B(n_3043),
.Y(n_3067)
);

AOI22xp5_ASAP7_75t_L g3068 ( 
.A1(n_3057),
.A2(n_3031),
.B1(n_2953),
.B2(n_2920),
.Y(n_3068)
);

AOI321xp33_ASAP7_75t_L g3069 ( 
.A1(n_3060),
.A2(n_2868),
.A3(n_3027),
.B1(n_3018),
.B2(n_3011),
.C(n_2973),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_3062),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_3052),
.B(n_2953),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_3055),
.B(n_3011),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_3062),
.B(n_2953),
.Y(n_3073)
);

OAI21xp33_ASAP7_75t_L g3074 ( 
.A1(n_3051),
.A2(n_2971),
.B(n_3018),
.Y(n_3074)
);

HB1xp67_ASAP7_75t_L g3075 ( 
.A(n_3061),
.Y(n_3075)
);

AND2x2_ASAP7_75t_L g3076 ( 
.A(n_3053),
.B(n_2973),
.Y(n_3076)
);

AOI22xp5_ASAP7_75t_L g3077 ( 
.A1(n_3048),
.A2(n_2971),
.B1(n_2908),
.B2(n_2978),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_3053),
.B(n_2978),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_3058),
.Y(n_3079)
);

OR2x2_ASAP7_75t_L g3080 ( 
.A(n_3072),
.B(n_3048),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_3075),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_SL g3082 ( 
.A(n_3065),
.B(n_3061),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_3064),
.B(n_3050),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_3072),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_3079),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_3067),
.Y(n_3086)
);

INVxp67_ASAP7_75t_L g3087 ( 
.A(n_3065),
.Y(n_3087)
);

O2A1O1Ixp33_ASAP7_75t_L g3088 ( 
.A1(n_3063),
.A2(n_2678),
.B(n_3027),
.C(n_2660),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_3076),
.B(n_2978),
.Y(n_3089)
);

AOI21xp33_ASAP7_75t_SL g3090 ( 
.A1(n_3074),
.A2(n_2678),
.B(n_2967),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_3070),
.B(n_3001),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_3078),
.B(n_2978),
.Y(n_3092)
);

XOR2x2_ASAP7_75t_L g3093 ( 
.A(n_3077),
.B(n_2667),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_3071),
.Y(n_3094)
);

NAND2x1p5_ASAP7_75t_L g3095 ( 
.A(n_3068),
.B(n_2681),
.Y(n_3095)
);

NAND3xp33_ASAP7_75t_L g3096 ( 
.A(n_3069),
.B(n_2775),
.C(n_2927),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_3073),
.Y(n_3097)
);

NAND2x1p5_ASAP7_75t_L g3098 ( 
.A(n_3066),
.B(n_2681),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_3064),
.B(n_2971),
.Y(n_3099)
);

A2O1A1Ixp33_ASAP7_75t_L g3100 ( 
.A1(n_3088),
.A2(n_2913),
.B(n_3001),
.C(n_2839),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_3087),
.B(n_2659),
.Y(n_3101)
);

O2A1O1Ixp33_ASAP7_75t_L g3102 ( 
.A1(n_3087),
.A2(n_2592),
.B(n_2967),
.C(n_2904),
.Y(n_3102)
);

NOR2xp33_ASAP7_75t_L g3103 ( 
.A(n_3096),
.B(n_2659),
.Y(n_3103)
);

NAND3xp33_ASAP7_75t_SL g3104 ( 
.A(n_3088),
.B(n_2735),
.C(n_2687),
.Y(n_3104)
);

NOR4xp75_ASAP7_75t_L g3105 ( 
.A(n_3082),
.B(n_2868),
.C(n_2929),
.D(n_2793),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_3081),
.Y(n_3106)
);

NOR2xp33_ASAP7_75t_L g3107 ( 
.A(n_3080),
.B(n_2679),
.Y(n_3107)
);

NOR3xp33_ASAP7_75t_L g3108 ( 
.A(n_3082),
.B(n_2761),
.C(n_2756),
.Y(n_3108)
);

OAI21xp33_ASAP7_75t_SL g3109 ( 
.A1(n_3083),
.A2(n_2904),
.B(n_2980),
.Y(n_3109)
);

INVxp67_ASAP7_75t_L g3110 ( 
.A(n_3084),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_3086),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_3098),
.B(n_2927),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_3091),
.Y(n_3113)
);

NAND2xp33_ASAP7_75t_SL g3114 ( 
.A(n_3085),
.B(n_2773),
.Y(n_3114)
);

OR2x2_ASAP7_75t_L g3115 ( 
.A(n_3091),
.B(n_2935),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_3097),
.Y(n_3116)
);

O2A1O1Ixp33_ASAP7_75t_SL g3117 ( 
.A1(n_3090),
.A2(n_3094),
.B(n_3093),
.C(n_3095),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_SL g3118 ( 
.A(n_3108),
.B(n_3095),
.Y(n_3118)
);

OAI211xp5_ASAP7_75t_L g3119 ( 
.A1(n_3110),
.A2(n_3099),
.B(n_3089),
.C(n_3092),
.Y(n_3119)
);

OAI211xp5_ASAP7_75t_L g3120 ( 
.A1(n_3111),
.A2(n_3098),
.B(n_2755),
.C(n_2918),
.Y(n_3120)
);

AOI21xp5_ASAP7_75t_L g3121 ( 
.A1(n_3117),
.A2(n_2930),
.B(n_2932),
.Y(n_3121)
);

AOI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_3104),
.A2(n_2679),
.B1(n_2699),
.B2(n_2850),
.Y(n_3122)
);

OAI321xp33_ASAP7_75t_L g3123 ( 
.A1(n_3106),
.A2(n_2918),
.A3(n_2839),
.B1(n_2932),
.B2(n_2929),
.C(n_2773),
.Y(n_3123)
);

OAI221xp5_ASAP7_75t_L g3124 ( 
.A1(n_3103),
.A2(n_2731),
.B1(n_2733),
.B2(n_2707),
.C(n_2722),
.Y(n_3124)
);

OAI211xp5_ASAP7_75t_L g3125 ( 
.A1(n_3101),
.A2(n_3116),
.B(n_3113),
.C(n_3107),
.Y(n_3125)
);

NAND4xp25_ASAP7_75t_L g3126 ( 
.A(n_3100),
.B(n_2850),
.C(n_2775),
.D(n_2980),
.Y(n_3126)
);

AND2x2_ASAP7_75t_L g3127 ( 
.A(n_3115),
.B(n_2935),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_3112),
.B(n_3102),
.Y(n_3128)
);

NAND3xp33_ASAP7_75t_SL g3129 ( 
.A(n_3105),
.B(n_2930),
.C(n_2850),
.Y(n_3129)
);

AOI211xp5_ASAP7_75t_L g3130 ( 
.A1(n_3109),
.A2(n_2773),
.B(n_2751),
.C(n_2850),
.Y(n_3130)
);

AOI211xp5_ASAP7_75t_L g3131 ( 
.A1(n_3125),
.A2(n_3114),
.B(n_2929),
.C(n_2961),
.Y(n_3131)
);

NOR4xp25_ASAP7_75t_L g3132 ( 
.A(n_3119),
.B(n_2956),
.C(n_2957),
.D(n_2963),
.Y(n_3132)
);

XNOR2xp5_ASAP7_75t_L g3133 ( 
.A(n_3122),
.B(n_2933),
.Y(n_3133)
);

O2A1O1Ixp33_ASAP7_75t_L g3134 ( 
.A1(n_3118),
.A2(n_2830),
.B(n_2843),
.C(n_2538),
.Y(n_3134)
);

AOI22xp5_ASAP7_75t_L g3135 ( 
.A1(n_3120),
.A2(n_2864),
.B1(n_2733),
.B2(n_2722),
.Y(n_3135)
);

AOI22xp5_ASAP7_75t_L g3136 ( 
.A1(n_3126),
.A2(n_2864),
.B1(n_2707),
.B2(n_2731),
.Y(n_3136)
);

AOI211xp5_ASAP7_75t_L g3137 ( 
.A1(n_3128),
.A2(n_2961),
.B(n_2942),
.C(n_2632),
.Y(n_3137)
);

OR3x1_ASAP7_75t_L g3138 ( 
.A(n_3123),
.B(n_2933),
.C(n_2921),
.Y(n_3138)
);

AOI211xp5_ASAP7_75t_L g3139 ( 
.A1(n_3121),
.A2(n_3130),
.B(n_3124),
.C(n_3127),
.Y(n_3139)
);

HB1xp67_ASAP7_75t_L g3140 ( 
.A(n_3129),
.Y(n_3140)
);

A2O1A1Ixp33_ASAP7_75t_L g3141 ( 
.A1(n_3121),
.A2(n_2830),
.B(n_2843),
.C(n_2803),
.Y(n_3141)
);

OAI22xp5_ASAP7_75t_L g3142 ( 
.A1(n_3120),
.A2(n_2896),
.B1(n_2830),
.B2(n_2843),
.Y(n_3142)
);

OAI211xp5_ASAP7_75t_L g3143 ( 
.A1(n_3125),
.A2(n_2854),
.B(n_2752),
.C(n_2504),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_3119),
.Y(n_3144)
);

AOI22xp33_ASAP7_75t_SL g3145 ( 
.A1(n_3144),
.A2(n_2896),
.B1(n_2658),
.B2(n_2864),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_3133),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_3140),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_3138),
.Y(n_3148)
);

OR2x2_ASAP7_75t_L g3149 ( 
.A(n_3132),
.B(n_2972),
.Y(n_3149)
);

NOR2x1_ASAP7_75t_L g3150 ( 
.A(n_3143),
.B(n_2972),
.Y(n_3150)
);

NAND4xp75_ASAP7_75t_L g3151 ( 
.A(n_3135),
.B(n_2974),
.C(n_2569),
.D(n_2784),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3131),
.Y(n_3152)
);

OAI221xp5_ASAP7_75t_L g3153 ( 
.A1(n_3139),
.A2(n_2854),
.B1(n_2525),
.B2(n_2849),
.C(n_2958),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3134),
.Y(n_3154)
);

NOR3xp33_ASAP7_75t_L g3155 ( 
.A(n_3142),
.B(n_2939),
.C(n_2974),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3137),
.Y(n_3156)
);

XNOR2xp5_ASAP7_75t_L g3157 ( 
.A(n_3136),
.B(n_2879),
.Y(n_3157)
);

NOR3xp33_ASAP7_75t_L g3158 ( 
.A(n_3141),
.B(n_2939),
.C(n_2797),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_3140),
.Y(n_3159)
);

NOR2x1_ASAP7_75t_L g3160 ( 
.A(n_3144),
.B(n_2972),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_3144),
.B(n_2972),
.Y(n_3161)
);

INVx1_ASAP7_75t_SL g3162 ( 
.A(n_3159),
.Y(n_3162)
);

NAND3xp33_ASAP7_75t_SL g3163 ( 
.A(n_3147),
.B(n_2958),
.C(n_2784),
.Y(n_3163)
);

NOR2xp67_ASAP7_75t_L g3164 ( 
.A(n_3152),
.B(n_2854),
.Y(n_3164)
);

AOI21xp5_ASAP7_75t_L g3165 ( 
.A1(n_3154),
.A2(n_2565),
.B(n_2854),
.Y(n_3165)
);

NAND3xp33_ASAP7_75t_L g3166 ( 
.A(n_3146),
.B(n_3148),
.C(n_3156),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_SL g3167 ( 
.A(n_3161),
.B(n_2854),
.Y(n_3167)
);

NOR4xp75_ASAP7_75t_L g3168 ( 
.A(n_3161),
.B(n_2934),
.C(n_2798),
.D(n_2814),
.Y(n_3168)
);

AND2x2_ASAP7_75t_SL g3169 ( 
.A(n_3149),
.B(n_2849),
.Y(n_3169)
);

NAND4xp75_ASAP7_75t_L g3170 ( 
.A(n_3160),
.B(n_2524),
.C(n_2957),
.D(n_2963),
.Y(n_3170)
);

OAI221xp5_ASAP7_75t_L g3171 ( 
.A1(n_3153),
.A2(n_2854),
.B1(n_2849),
.B2(n_2529),
.C(n_2560),
.Y(n_3171)
);

NAND2x2_ASAP7_75t_L g3172 ( 
.A(n_3157),
.B(n_2934),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_3150),
.Y(n_3173)
);

NOR3xp33_ASAP7_75t_L g3174 ( 
.A(n_3145),
.B(n_2837),
.C(n_2869),
.Y(n_3174)
);

O2A1O1Ixp33_ASAP7_75t_L g3175 ( 
.A1(n_3158),
.A2(n_2975),
.B(n_2969),
.C(n_2951),
.Y(n_3175)
);

AOI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_3162),
.A2(n_3155),
.B1(n_3151),
.B2(n_2864),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_3169),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3166),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3164),
.Y(n_3179)
);

OAI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_3167),
.A2(n_2975),
.B(n_2969),
.Y(n_3180)
);

AOI21xp5_ASAP7_75t_L g3181 ( 
.A1(n_3173),
.A2(n_2975),
.B(n_2943),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_3170),
.Y(n_3182)
);

AOI22x1_ASAP7_75t_L g3183 ( 
.A1(n_3165),
.A2(n_2849),
.B1(n_2951),
.B2(n_2950),
.Y(n_3183)
);

AOI21x1_ASAP7_75t_L g3184 ( 
.A1(n_3172),
.A2(n_2969),
.B(n_2951),
.Y(n_3184)
);

NAND3xp33_ASAP7_75t_SL g3185 ( 
.A(n_3171),
.B(n_2950),
.C(n_2921),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_3174),
.Y(n_3186)
);

AND3x1_ASAP7_75t_L g3187 ( 
.A(n_3175),
.B(n_2950),
.C(n_2941),
.Y(n_3187)
);

AOI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_3178),
.A2(n_3163),
.B1(n_3168),
.B2(n_2896),
.Y(n_3188)
);

OAI22xp5_ASAP7_75t_L g3189 ( 
.A1(n_3176),
.A2(n_2849),
.B1(n_2837),
.B2(n_2941),
.Y(n_3189)
);

BUFx6f_ASAP7_75t_L g3190 ( 
.A(n_3177),
.Y(n_3190)
);

AO22x2_ASAP7_75t_L g3191 ( 
.A1(n_3186),
.A2(n_2795),
.B1(n_2799),
.B2(n_2808),
.Y(n_3191)
);

OAI22x1_ASAP7_75t_L g3192 ( 
.A1(n_3182),
.A2(n_2941),
.B1(n_2931),
.B2(n_2810),
.Y(n_3192)
);

AOI22xp5_ASAP7_75t_L g3193 ( 
.A1(n_3176),
.A2(n_2725),
.B1(n_2800),
.B2(n_2807),
.Y(n_3193)
);

INVxp67_ASAP7_75t_SL g3194 ( 
.A(n_3179),
.Y(n_3194)
);

AOI22xp5_ASAP7_75t_L g3195 ( 
.A1(n_3185),
.A2(n_2725),
.B1(n_2800),
.B2(n_2807),
.Y(n_3195)
);

AO22x2_ASAP7_75t_L g3196 ( 
.A1(n_3181),
.A2(n_2909),
.B1(n_2907),
.B2(n_2819),
.Y(n_3196)
);

HB1xp67_ASAP7_75t_L g3197 ( 
.A(n_3190),
.Y(n_3197)
);

OAI22x1_ASAP7_75t_SL g3198 ( 
.A1(n_3194),
.A2(n_3184),
.B1(n_3183),
.B2(n_3187),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3188),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_3191),
.Y(n_3200)
);

OAI22xp5_ASAP7_75t_SL g3201 ( 
.A1(n_3193),
.A2(n_3180),
.B1(n_2909),
.B2(n_2907),
.Y(n_3201)
);

OR2x2_ASAP7_75t_L g3202 ( 
.A(n_3189),
.B(n_3195),
.Y(n_3202)
);

CKINVDCx20_ASAP7_75t_R g3203 ( 
.A(n_3197),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_3199),
.Y(n_3204)
);

OAI22x1_ASAP7_75t_L g3205 ( 
.A1(n_3200),
.A2(n_3196),
.B1(n_3192),
.B2(n_2817),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3198),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_3204),
.B(n_3202),
.Y(n_3207)
);

AO21x1_ASAP7_75t_L g3208 ( 
.A1(n_3206),
.A2(n_3201),
.B(n_2812),
.Y(n_3208)
);

OA21x2_ASAP7_75t_L g3209 ( 
.A1(n_3207),
.A2(n_3203),
.B(n_3205),
.Y(n_3209)
);

OA21x2_ASAP7_75t_L g3210 ( 
.A1(n_3209),
.A2(n_3208),
.B(n_2562),
.Y(n_3210)
);

AOI22x1_ASAP7_75t_L g3211 ( 
.A1(n_3210),
.A2(n_2817),
.B1(n_2915),
.B2(n_2819),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3210),
.Y(n_3212)
);

OAI221xp5_ASAP7_75t_R g3213 ( 
.A1(n_3212),
.A2(n_2813),
.B1(n_2833),
.B2(n_2915),
.C(n_2816),
.Y(n_3213)
);

AOI211xp5_ASAP7_75t_L g3214 ( 
.A1(n_3213),
.A2(n_3211),
.B(n_2816),
.C(n_2812),
.Y(n_3214)
);


endmodule