module fake_jpeg_26901_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_0),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_25),
.B(n_1),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_1),
.B(n_2),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_44),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_20),
.B1(n_13),
.B2(n_22),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_13),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_17),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_18),
.B1(n_22),
.B2(n_19),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_24),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_53),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_21),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_35),
.B1(n_34),
.B2(n_43),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_17),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_30),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_57),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_48),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_73),
.C(n_64),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_69),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_45),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_55),
.B1(n_38),
.B2(n_43),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_84),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_87),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_86),
.Y(n_95)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_56),
.B1(n_40),
.B2(n_46),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_70),
.B(n_61),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_74),
.B(n_70),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_96),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_88),
.C(n_78),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_94),
.C(n_97),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_71),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_21),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_28),
.C(n_30),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_75),
.B(n_2),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_23),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_105),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_85),
.C(n_87),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_104),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_83),
.B(n_82),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_108),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_103),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_3),
.B(n_7),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_100),
.C(n_26),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_113),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_95),
.B(n_10),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_77),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_115),
.A2(n_60),
.B1(n_62),
.B2(n_14),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_118),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_79),
.C(n_16),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_14),
.C(n_16),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_120),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_14),
.C(n_16),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_8),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_12),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_12),
.C(n_125),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_8),
.B(n_10),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_128),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_123),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_129),
.Y(n_131)
);


endmodule