module fake_jpeg_2649_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_61),
.Y(n_66)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_1),
.Y(n_74)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_53),
.B1(n_47),
.B2(n_40),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_73),
.B1(n_49),
.B2(n_51),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_41),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_55),
.B1(n_43),
.B2(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_65),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_81),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_55),
.B1(n_47),
.B2(n_52),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_88),
.Y(n_95)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_54),
.C(n_52),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_49),
.B(n_46),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_108)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_3),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_22),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_21),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_23),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_103),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_6),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_6),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_7),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_28),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_87),
.B1(n_76),
.B2(n_12),
.Y(n_112)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_124),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_116),
.B1(n_32),
.B2(n_33),
.Y(n_135)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_98),
.B1(n_100),
.B2(n_108),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_122),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_27),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_123),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_13),
.B(n_14),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_121),
.A2(n_20),
.B(n_24),
.Y(n_128)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_26),
.B(n_30),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_135),
.B1(n_121),
.B2(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_25),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_132),
.B(n_134),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_137),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_140),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_116),
.B(n_110),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_140),
.B(n_133),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_143),
.A2(n_129),
.B1(n_125),
.B2(n_127),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_145),
.C(n_117),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_139),
.C(n_136),
.Y(n_147)
);

OAI321xp33_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_124),
.A3(n_141),
.B1(n_135),
.B2(n_128),
.C(n_115),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_110),
.C(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_34),
.C(n_36),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_37),
.Y(n_152)
);


endmodule