module fake_jpeg_11997_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx3_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx8_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_22),
.Y(n_34)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_6),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_8),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_9),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_36),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_0),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_40),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_41),
.B1(n_46),
.B2(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_19),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_23),
.B1(n_22),
.B2(n_9),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_11),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_28),
.B1(n_27),
.B2(n_11),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_17),
.B(n_10),
.C(n_16),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_48),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_45),
.B1(n_43),
.B2(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_49),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_61),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_45),
.B(n_50),
.Y(n_62)
);

AO221x1_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_63),
.B1(n_56),
.B2(n_57),
.C(n_10),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_47),
.B(n_54),
.C(n_17),
.Y(n_63)
);

AO21x1_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_66),
.B(n_10),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_29),
.B(n_58),
.C(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_0),
.Y(n_70)
);

AOI222xp33_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_66),
.B1(n_18),
.B2(n_25),
.C1(n_1),
.C2(n_3),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_70),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g72 ( 
.A(n_71),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_27),
.C(n_1),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_0),
.Y(n_74)
);


endmodule