module fake_aes_1482_n_1457 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1457);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1457;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_533;
wire n_1010;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_659;
wire n_386;
wire n_432;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1454;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1439;
wire n_374;
wire n_718;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1219;
wire n_1120;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g328 ( .A(n_82), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_300), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_310), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_317), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_216), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_112), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_175), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_253), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_322), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_60), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_326), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_201), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_314), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_101), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_205), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_108), .Y(n_343) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_258), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_248), .Y(n_345) );
INVxp67_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_10), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_143), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_100), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_142), .Y(n_350) );
INVxp33_ASAP7_75t_SL g351 ( .A(n_98), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_55), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_41), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_213), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_254), .Y(n_355) );
CKINVDCx16_ASAP7_75t_R g356 ( .A(n_32), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_119), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_319), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_202), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_36), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_56), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_269), .Y(n_362) );
INVxp33_ASAP7_75t_SL g363 ( .A(n_20), .Y(n_363) );
CKINVDCx16_ASAP7_75t_R g364 ( .A(n_320), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_104), .Y(n_365) );
INVxp67_ASAP7_75t_L g366 ( .A(n_237), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_19), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_170), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_148), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_78), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_239), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_93), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_186), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_64), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_69), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_0), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_147), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_193), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_294), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_195), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_35), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_73), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_12), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_297), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_96), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_46), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_34), .Y(n_387) );
CKINVDCx14_ASAP7_75t_R g388 ( .A(n_64), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_70), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_144), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_63), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_164), .Y(n_392) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_215), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_296), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_257), .Y(n_395) );
CKINVDCx16_ASAP7_75t_R g396 ( .A(n_86), .Y(n_396) );
INVxp33_ASAP7_75t_L g397 ( .A(n_183), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_61), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_292), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_220), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_318), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_24), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_263), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_228), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_165), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_232), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_125), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_19), .Y(n_408) );
INVxp33_ASAP7_75t_SL g409 ( .A(n_184), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_65), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_65), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_238), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_149), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_49), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_7), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_30), .B(n_118), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_9), .Y(n_417) );
INVxp33_ASAP7_75t_SL g418 ( .A(n_100), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_18), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_264), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_51), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_282), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_265), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_226), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_59), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_153), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_187), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_83), .Y(n_428) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_261), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_10), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_72), .Y(n_431) );
INVxp67_ASAP7_75t_L g432 ( .A(n_306), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_1), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_192), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_95), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_28), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_225), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_163), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_13), .Y(n_439) );
CKINVDCx16_ASAP7_75t_R g440 ( .A(n_92), .Y(n_440) );
INVxp33_ASAP7_75t_L g441 ( .A(n_245), .Y(n_441) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_94), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_323), .B(n_235), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_2), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_229), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_101), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_167), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_321), .Y(n_448) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_35), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_92), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_252), .Y(n_451) );
NOR2xp67_ASAP7_75t_L g452 ( .A(n_161), .B(n_1), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_293), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_272), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_5), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_295), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_87), .Y(n_457) );
INVxp33_ASAP7_75t_L g458 ( .A(n_59), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_223), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_120), .B(n_87), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_139), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_97), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_0), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_103), .Y(n_464) );
INVxp67_ASAP7_75t_L g465 ( .A(n_256), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_173), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_284), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_204), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_206), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_85), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_224), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_327), .Y(n_472) );
INVxp33_ASAP7_75t_SL g473 ( .A(n_80), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_131), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_111), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_55), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_315), .Y(n_477) );
BUFx3_ASAP7_75t_L g478 ( .A(n_5), .Y(n_478) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_210), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_271), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_285), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_194), .Y(n_482) );
BUFx3_ASAP7_75t_L g483 ( .A(n_132), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_176), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_36), .Y(n_485) );
INVxp33_ASAP7_75t_SL g486 ( .A(n_324), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_50), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_298), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_20), .Y(n_489) );
INVxp33_ASAP7_75t_L g490 ( .A(n_130), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_134), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_137), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_251), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_188), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_3), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_399), .Y(n_496) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_399), .Y(n_497) );
NAND2xp33_ASAP7_75t_L g498 ( .A(n_374), .B(n_109), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_368), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_388), .Y(n_500) );
BUFx2_ASAP7_75t_L g501 ( .A(n_402), .Y(n_501) );
BUFx2_ASAP7_75t_L g502 ( .A(n_402), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_368), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_399), .Y(n_504) );
NOR2xp33_ASAP7_75t_SL g505 ( .A(n_364), .B(n_477), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_371), .Y(n_506) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_399), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_371), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_494), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_456), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_458), .B(n_2), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_458), .B(n_3), .Y(n_512) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_399), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_397), .B(n_4), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_356), .B(n_4), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_494), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_456), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_339), .B(n_6), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_329), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_385), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_403), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_456), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_397), .B(n_6), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_385), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_460), .B(n_7), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_387), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_387), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_460), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_403), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_367), .B(n_8), .Y(n_530) );
INVx4_ASAP7_75t_L g531 ( .A(n_460), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_441), .B(n_8), .Y(n_532) );
OR2x6_ASAP7_75t_L g533 ( .A(n_416), .B(n_9), .Y(n_533) );
AND2x4_ASAP7_75t_SL g534 ( .A(n_533), .B(n_329), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_501), .B(n_441), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_511), .A2(n_363), .B1(n_418), .B2(n_351), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_497), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_500), .Y(n_538) );
INVx5_ASAP7_75t_L g539 ( .A(n_522), .Y(n_539) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_497), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_522), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_501), .B(n_490), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_501), .B(n_490), .Y(n_543) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_512), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_497), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_522), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_497), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_531), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_522), .Y(n_549) );
INVx3_ASAP7_75t_L g550 ( .A(n_531), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_522), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_510), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_502), .B(n_528), .Y(n_553) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_497), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_500), .B(n_396), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_497), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_502), .B(n_431), .Y(n_557) );
NAND2xp33_ASAP7_75t_L g558 ( .A(n_528), .B(n_403), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_497), .Y(n_559) );
AO22x2_ASAP7_75t_L g560 ( .A1(n_525), .A2(n_416), .B1(n_358), .B2(n_394), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_497), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_502), .B(n_431), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_528), .B(n_334), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_507), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_528), .B(n_334), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_511), .A2(n_363), .B1(n_418), .B2(n_351), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_510), .Y(n_567) );
BUFx3_ASAP7_75t_L g568 ( .A(n_525), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_510), .Y(n_569) );
INVx4_ASAP7_75t_SL g570 ( .A(n_525), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_525), .B(n_358), .Y(n_571) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_507), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_531), .Y(n_573) );
NAND2xp33_ASAP7_75t_L g574 ( .A(n_528), .B(n_403), .Y(n_574) );
AND2x6_ASAP7_75t_L g575 ( .A(n_525), .B(n_340), .Y(n_575) );
INVx5_ASAP7_75t_L g576 ( .A(n_507), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_544), .B(n_533), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_539), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_539), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_543), .B(n_505), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_544), .B(n_533), .Y(n_581) );
BUFx3_ASAP7_75t_L g582 ( .A(n_575), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_560), .A2(n_533), .B1(n_511), .B2(n_532), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_535), .B(n_523), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_534), .A2(n_533), .B1(n_330), .B2(n_380), .Y(n_585) );
NAND2x1p5_ASAP7_75t_L g586 ( .A(n_568), .B(n_523), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_535), .B(n_523), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_560), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_539), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_552), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_570), .B(n_505), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_539), .Y(n_592) );
BUFx12f_ASAP7_75t_L g593 ( .A(n_555), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_543), .B(n_532), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_534), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_538), .B(n_515), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_552), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_570), .B(n_533), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_539), .Y(n_599) );
BUFx12f_ASAP7_75t_L g600 ( .A(n_555), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_539), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_535), .B(n_532), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_539), .Y(n_603) );
BUFx12f_ASAP7_75t_SL g604 ( .A(n_542), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_539), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_542), .B(n_499), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_567), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_548), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_570), .B(n_518), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_570), .B(n_533), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_570), .B(n_531), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_548), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_548), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_567), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_569), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g616 ( .A1(n_568), .A2(n_503), .B(n_506), .C(n_499), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_569), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_542), .B(n_503), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_538), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_534), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_553), .A2(n_512), .B(n_514), .C(n_518), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_541), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_548), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_548), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_550), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_541), .Y(n_626) );
INVx4_ASAP7_75t_L g627 ( .A(n_570), .Y(n_627) );
INVx5_ASAP7_75t_L g628 ( .A(n_575), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_546), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_546), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_551), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_550), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_551), .Y(n_633) );
INVx3_ASAP7_75t_L g634 ( .A(n_568), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_553), .B(n_506), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_568), .Y(n_636) );
NAND3xp33_ASAP7_75t_SL g637 ( .A(n_536), .B(n_566), .C(n_519), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_550), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g639 ( .A(n_550), .B(n_531), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_555), .B(n_508), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_549), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_550), .Y(n_642) );
INVx3_ASAP7_75t_L g643 ( .A(n_573), .Y(n_643) );
INVx4_ASAP7_75t_L g644 ( .A(n_575), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_557), .B(n_508), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_560), .A2(n_516), .B1(n_509), .B2(n_515), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_557), .B(n_509), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_536), .B(n_515), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_549), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_549), .Y(n_650) );
BUFx2_ASAP7_75t_L g651 ( .A(n_560), .Y(n_651) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_575), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_573), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_557), .B(n_516), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_588), .A2(n_560), .B1(n_575), .B2(n_571), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_588), .Y(n_656) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_652), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_651), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_594), .B(n_562), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_596), .B(n_566), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_598), .B(n_534), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_598), .B(n_610), .Y(n_662) );
BUFx3_ASAP7_75t_L g663 ( .A(n_652), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_596), .B(n_562), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_608), .A2(n_571), .B(n_573), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_608), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_651), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_608), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_586), .Y(n_669) );
BUFx3_ASAP7_75t_L g670 ( .A(n_652), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_586), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_619), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_648), .B(n_562), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_586), .Y(n_674) );
A2O1A1Ixp33_ASAP7_75t_L g675 ( .A1(n_621), .A2(n_565), .B(n_563), .C(n_530), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_577), .A2(n_560), .B1(n_575), .B2(n_573), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_585), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_584), .A2(n_602), .B1(n_587), .B2(n_640), .C(n_637), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_598), .B(n_575), .Y(n_679) );
AND2x4_ASAP7_75t_SL g680 ( .A(n_598), .B(n_330), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_584), .B(n_440), .Y(n_681) );
INVx3_ASAP7_75t_L g682 ( .A(n_627), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_612), .A2(n_573), .B(n_565), .Y(n_683) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_648), .A2(n_514), .B1(n_530), .B2(n_449), .C(n_442), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g685 ( .A1(n_583), .A2(n_380), .B1(n_424), .B2(n_362), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_652), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_590), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_612), .Y(n_688) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_652), .Y(n_689) );
INVx3_ASAP7_75t_L g690 ( .A(n_627), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_580), .B(n_574), .C(n_558), .Y(n_691) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_583), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_612), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_577), .A2(n_575), .B1(n_424), .B2(n_454), .Y(n_694) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_652), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_613), .A2(n_563), .B(n_558), .Y(n_696) );
NAND2x1p5_ASAP7_75t_L g697 ( .A(n_627), .B(n_478), .Y(n_697) );
INVx3_ASAP7_75t_SL g698 ( .A(n_610), .Y(n_698) );
NAND3xp33_ASAP7_75t_SL g699 ( .A(n_646), .B(n_454), .C(n_362), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_590), .Y(n_700) );
AOI21x1_ASAP7_75t_L g701 ( .A1(n_609), .A2(n_517), .B(n_537), .Y(n_701) );
NOR2xp33_ASAP7_75t_SL g702 ( .A(n_644), .B(n_466), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_587), .B(n_575), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_613), .Y(n_704) );
INVx2_ASAP7_75t_SL g705 ( .A(n_593), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_597), .Y(n_706) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_606), .B(n_466), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_597), .Y(n_708) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_610), .Y(n_709) );
BUFx2_ASAP7_75t_L g710 ( .A(n_604), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_602), .B(n_398), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_618), .B(n_337), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_645), .B(n_575), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_604), .B(n_473), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_593), .B(n_337), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_595), .A2(n_474), .B1(n_469), .B2(n_389), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_613), .Y(n_717) );
CKINVDCx11_ASAP7_75t_R g718 ( .A(n_600), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_595), .A2(n_474), .B1(n_469), .B2(n_389), .Y(n_719) );
INVx2_ASAP7_75t_SL g720 ( .A(n_600), .Y(n_720) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_610), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_625), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_582), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_647), .B(n_473), .Y(n_724) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_611), .Y(n_725) );
NAND3xp33_ASAP7_75t_L g726 ( .A(n_616), .B(n_591), .C(n_654), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_607), .Y(n_727) );
BUFx2_ASAP7_75t_L g728 ( .A(n_577), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_635), .B(n_409), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_625), .Y(n_730) );
INVx4_ASAP7_75t_L g731 ( .A(n_627), .Y(n_731) );
AOI21xp33_ASAP7_75t_L g732 ( .A1(n_620), .A2(n_574), .B(n_486), .Y(n_732) );
BUFx2_ASAP7_75t_L g733 ( .A(n_577), .Y(n_733) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_611), .Y(n_734) );
BUFx2_ASAP7_75t_L g735 ( .A(n_581), .Y(n_735) );
BUFx2_ASAP7_75t_L g736 ( .A(n_581), .Y(n_736) );
INVx3_ASAP7_75t_L g737 ( .A(n_611), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_581), .B(n_343), .Y(n_738) );
INVx4_ASAP7_75t_L g739 ( .A(n_628), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_607), .Y(n_740) );
BUFx2_ASAP7_75t_SL g741 ( .A(n_628), .Y(n_741) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_582), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_581), .A2(n_517), .B1(n_486), .B2(n_409), .Y(n_743) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_611), .Y(n_744) );
O2A1O1Ixp5_ASAP7_75t_L g745 ( .A1(n_644), .A2(n_393), .B(n_429), .C(n_344), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_614), .Y(n_746) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_582), .Y(n_747) );
INVx3_ASAP7_75t_L g748 ( .A(n_636), .Y(n_748) );
INVx4_ASAP7_75t_L g749 ( .A(n_628), .Y(n_749) );
INVx2_ASAP7_75t_SL g750 ( .A(n_628), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_644), .A2(n_517), .B1(n_478), .B2(n_370), .Y(n_751) );
BUFx2_ASAP7_75t_L g752 ( .A(n_620), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_614), .A2(n_524), .B(n_526), .C(n_520), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_615), .B(n_376), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_615), .Y(n_755) );
INVxp67_ASAP7_75t_L g756 ( .A(n_617), .Y(n_756) );
BUFx6f_ASAP7_75t_L g757 ( .A(n_628), .Y(n_757) );
BUFx4f_ASAP7_75t_L g758 ( .A(n_639), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_644), .B(n_331), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_617), .A2(n_634), .B1(n_636), .B2(n_653), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_634), .B(n_331), .Y(n_761) );
AOI221x1_ASAP7_75t_L g762 ( .A1(n_641), .A2(n_333), .B1(n_336), .B2(n_335), .C(n_332), .Y(n_762) );
INVx4_ASAP7_75t_L g763 ( .A(n_628), .Y(n_763) );
INVx2_ASAP7_75t_SL g764 ( .A(n_639), .Y(n_764) );
INVx4_ASAP7_75t_L g765 ( .A(n_636), .Y(n_765) );
INVx1_ASAP7_75t_SL g766 ( .A(n_680), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_754), .Y(n_767) );
BUFx12f_ASAP7_75t_L g768 ( .A(n_718), .Y(n_768) );
AOI222xp33_ASAP7_75t_L g769 ( .A1(n_678), .A2(n_476), .B1(n_343), .B2(n_415), .C1(n_391), .C2(n_450), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_687), .Y(n_770) );
AND2x6_ASAP7_75t_L g771 ( .A(n_661), .B(n_634), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_661), .B(n_634), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_737), .Y(n_773) );
INVx1_ASAP7_75t_SL g774 ( .A(n_680), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_699), .A2(n_643), .B1(n_636), .B2(n_391), .Y(n_775) );
A2O1A1Ixp33_ASAP7_75t_L g776 ( .A1(n_675), .A2(n_643), .B(n_622), .C(n_629), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_738), .B(n_415), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_677), .A2(n_643), .B1(n_636), .B2(n_476), .Y(n_778) );
NOR2xp67_ASAP7_75t_L g779 ( .A(n_672), .B(n_11), .Y(n_779) );
INVx4_ASAP7_75t_L g780 ( .A(n_758), .Y(n_780) );
OAI222xp33_ASAP7_75t_L g781 ( .A1(n_685), .A2(n_375), .B1(n_370), .B2(n_367), .C1(n_341), .C2(n_347), .Y(n_781) );
BUFx8_ASAP7_75t_SL g782 ( .A(n_672), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_660), .B(n_643), .Y(n_783) );
AND2x4_ASAP7_75t_L g784 ( .A(n_661), .B(n_636), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_700), .Y(n_785) );
AND2x4_ASAP7_75t_L g786 ( .A(n_669), .B(n_622), .Y(n_786) );
INVx3_ASAP7_75t_L g787 ( .A(n_758), .Y(n_787) );
BUFx2_ASAP7_75t_L g788 ( .A(n_679), .Y(n_788) );
BUFx3_ASAP7_75t_L g789 ( .A(n_718), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_706), .Y(n_790) );
NAND2x1p5_ASAP7_75t_L g791 ( .A(n_662), .B(n_626), .Y(n_791) );
OAI221xp5_ASAP7_75t_L g792 ( .A1(n_684), .A2(n_349), .B1(n_353), .B2(n_352), .C(n_328), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_708), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_677), .A2(n_632), .B1(n_638), .B2(n_625), .Y(n_794) );
INVx1_ASAP7_75t_SL g795 ( .A(n_698), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g796 ( .A1(n_675), .A2(n_629), .B(n_626), .Y(n_796) );
AND2x4_ASAP7_75t_L g797 ( .A(n_671), .B(n_630), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_727), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_740), .B(n_630), .Y(n_799) );
INVx3_ASAP7_75t_L g800 ( .A(n_731), .Y(n_800) );
AND2x4_ASAP7_75t_L g801 ( .A(n_674), .B(n_631), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_692), .A2(n_632), .B1(n_642), .B2(n_638), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_685), .A2(n_632), .B1(n_642), .B2(n_638), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_746), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_712), .B(n_664), .Y(n_805) );
AOI21xp5_ASAP7_75t_SL g806 ( .A1(n_679), .A2(n_649), .B(n_641), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_656), .A2(n_653), .B1(n_642), .B2(n_633), .Y(n_807) );
AND2x4_ASAP7_75t_L g808 ( .A(n_662), .B(n_631), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_656), .A2(n_653), .B1(n_633), .B2(n_624), .Y(n_809) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_710), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_737), .Y(n_811) );
AND2x4_ASAP7_75t_L g812 ( .A(n_662), .B(n_623), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_755), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_665), .A2(n_650), .B(n_649), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_728), .A2(n_624), .B1(n_623), .B2(n_639), .Y(n_815) );
BUFx2_ASAP7_75t_L g816 ( .A(n_679), .Y(n_816) );
INVx4_ASAP7_75t_L g817 ( .A(n_698), .Y(n_817) );
NOR2xp33_ASAP7_75t_SL g818 ( .A(n_702), .B(n_342), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_666), .Y(n_819) );
NOR2xp67_ASAP7_75t_L g820 ( .A(n_705), .B(n_11), .Y(n_820) );
O2A1O1Ixp5_ASAP7_75t_L g821 ( .A1(n_745), .A2(n_650), .B(n_479), .C(n_524), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_716), .A2(n_342), .B1(n_348), .B2(n_345), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_673), .Y(n_823) );
O2A1O1Ixp33_ASAP7_75t_SL g824 ( .A1(n_753), .A2(n_350), .B(n_354), .C(n_338), .Y(n_824) );
INVx6_ASAP7_75t_L g825 ( .A(n_715), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_681), .B(n_520), .Y(n_826) );
OR2x2_ASAP7_75t_L g827 ( .A(n_716), .B(n_526), .Y(n_827) );
OR2x2_ASAP7_75t_L g828 ( .A(n_719), .B(n_527), .Y(n_828) );
INVx1_ASAP7_75t_SL g829 ( .A(n_733), .Y(n_829) );
AND2x4_ASAP7_75t_L g830 ( .A(n_735), .B(n_578), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_736), .A2(n_579), .B1(n_589), .B2(n_578), .Y(n_831) );
OR2x6_ASAP7_75t_L g832 ( .A(n_720), .B(n_411), .Y(n_832) );
OR2x2_ASAP7_75t_L g833 ( .A(n_719), .B(n_527), .Y(n_833) );
AO31x2_ASAP7_75t_L g834 ( .A1(n_762), .A2(n_504), .A3(n_521), .B(n_496), .Y(n_834) );
OAI21x1_ASAP7_75t_L g835 ( .A1(n_701), .A2(n_422), .B(n_394), .Y(n_835) );
BUFx8_ASAP7_75t_L g836 ( .A(n_709), .Y(n_836) );
OAI211xp5_ASAP7_75t_L g837 ( .A1(n_743), .A2(n_452), .B(n_361), .C(n_365), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_658), .A2(n_605), .B1(n_579), .B2(n_589), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_725), .Y(n_839) );
INVxp67_ASAP7_75t_SL g840 ( .A(n_723), .Y(n_840) );
NAND2x1p5_ASAP7_75t_L g841 ( .A(n_709), .B(n_578), .Y(n_841) );
AND2x4_ASAP7_75t_L g842 ( .A(n_764), .B(n_579), .Y(n_842) );
INVx4_ASAP7_75t_L g843 ( .A(n_709), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_659), .B(n_589), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_725), .Y(n_845) );
AND2x4_ASAP7_75t_L g846 ( .A(n_734), .B(n_592), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_711), .B(n_360), .Y(n_847) );
NAND2x1p5_ASAP7_75t_L g848 ( .A(n_709), .B(n_592), .Y(n_848) );
INVx4_ASAP7_75t_SL g849 ( .A(n_721), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_667), .A2(n_605), .B1(n_599), .B2(n_601), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_714), .B(n_592), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_734), .Y(n_852) );
AND2x6_ASAP7_75t_L g853 ( .A(n_721), .B(n_599), .Y(n_853) );
BUFx6f_ASAP7_75t_L g854 ( .A(n_657), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_666), .Y(n_855) );
AOI222xp33_ASAP7_75t_L g856 ( .A1(n_724), .A2(n_383), .B1(n_381), .B2(n_386), .C1(n_382), .C2(n_372), .Y(n_856) );
BUFx2_ASAP7_75t_L g857 ( .A(n_723), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_744), .Y(n_858) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_721), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_668), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_714), .A2(n_605), .B1(n_601), .B2(n_603), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_744), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g863 ( .A1(n_752), .A2(n_345), .B1(n_369), .B2(n_348), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_676), .A2(n_601), .B1(n_603), .B2(n_599), .Y(n_864) );
OAI21x1_ASAP7_75t_L g865 ( .A1(n_697), .A2(n_459), .B(n_422), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_676), .A2(n_433), .B1(n_435), .B2(n_411), .Y(n_866) );
INVx2_ASAP7_75t_SL g867 ( .A(n_707), .Y(n_867) );
BUFx8_ASAP7_75t_L g868 ( .A(n_721), .Y(n_868) );
INVx8_ASAP7_75t_L g869 ( .A(n_757), .Y(n_869) );
AOI21xp5_ASAP7_75t_SL g870 ( .A1(n_657), .A2(n_379), .B(n_340), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_694), .A2(n_603), .B1(n_408), .B2(n_414), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_729), .A2(n_392), .B1(n_445), .B2(n_369), .Y(n_872) );
BUFx3_ASAP7_75t_L g873 ( .A(n_697), .Y(n_873) );
AOI22xp33_ASAP7_75t_SL g874 ( .A1(n_756), .A2(n_445), .B1(n_447), .B2(n_392), .Y(n_874) );
OR2x2_ASAP7_75t_L g875 ( .A(n_743), .B(n_410), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_703), .B(n_417), .Y(n_876) );
BUFx3_ASAP7_75t_L g877 ( .A(n_731), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_668), .Y(n_878) );
INVx3_ASAP7_75t_L g879 ( .A(n_682), .Y(n_879) );
O2A1O1Ixp33_ASAP7_75t_SL g880 ( .A1(n_753), .A2(n_355), .B(n_359), .C(n_357), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_655), .A2(n_421), .B1(n_425), .B2(n_419), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_655), .A2(n_435), .B1(n_470), .B2(n_433), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_688), .Y(n_883) );
BUFx6f_ASAP7_75t_L g884 ( .A(n_657), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_713), .B(n_428), .Y(n_885) );
NOR3xp33_ASAP7_75t_L g886 ( .A(n_726), .B(n_436), .C(n_430), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_761), .A2(n_444), .B1(n_446), .B2(n_439), .Y(n_887) );
OAI221xp5_ASAP7_75t_L g888 ( .A1(n_751), .A2(n_462), .B1(n_463), .B2(n_457), .C(n_455), .Y(n_888) );
OAI222xp33_ASAP7_75t_L g889 ( .A1(n_751), .A2(n_485), .B1(n_489), .B2(n_487), .C1(n_464), .C2(n_470), .Y(n_889) );
AOI21xp5_ASAP7_75t_L g890 ( .A1(n_696), .A2(n_498), .B(n_556), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_805), .B(n_688), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_886), .A2(n_495), .B1(n_374), .B2(n_693), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_823), .B(n_693), .Y(n_893) );
AOI221xp5_ASAP7_75t_L g894 ( .A1(n_781), .A2(n_732), .B1(n_495), .B2(n_683), .C(n_691), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_777), .B(n_704), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_792), .A2(n_759), .B1(n_374), .B2(n_760), .C(n_717), .Y(n_896) );
AOI222xp33_ASAP7_75t_L g897 ( .A1(n_767), .A2(n_374), .B1(n_759), .B2(n_346), .C1(n_366), .C2(n_432), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_769), .B(n_704), .Y(n_898) );
OAI21x1_ASAP7_75t_L g899 ( .A1(n_835), .A2(n_748), .B(n_760), .Y(n_899) );
A2O1A1Ixp33_ASAP7_75t_L g900 ( .A1(n_796), .A2(n_722), .B(n_730), .C(n_717), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_769), .B(n_722), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_783), .A2(n_374), .B1(n_730), .B2(n_765), .Y(n_902) );
INVx1_ASAP7_75t_SL g903 ( .A(n_857), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_803), .B(n_765), .Y(n_904) );
BUFx2_ASAP7_75t_L g905 ( .A(n_836), .Y(n_905) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_778), .A2(n_765), .B1(n_747), .B2(n_742), .Y(n_906) );
INVx1_ASAP7_75t_SL g907 ( .A(n_825), .Y(n_907) );
OAI211xp5_ASAP7_75t_SL g908 ( .A1(n_856), .A2(n_465), .B(n_377), .C(n_378), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_888), .A2(n_748), .B1(n_747), .B2(n_742), .Y(n_909) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_818), .A2(n_690), .B1(n_682), .B2(n_468), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_770), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_819), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_888), .A2(n_747), .B1(n_742), .B2(n_670), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_855), .Y(n_914) );
AOI222xp33_ASAP7_75t_L g915 ( .A1(n_847), .A2(n_472), .B1(n_384), .B2(n_390), .C1(n_395), .C2(n_400), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_866), .A2(n_747), .B1(n_742), .B2(n_670), .Y(n_916) );
OR2x2_ASAP7_75t_L g917 ( .A(n_766), .B(n_690), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_866), .A2(n_686), .B1(n_663), .B2(n_379), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_775), .A2(n_663), .B1(n_686), .B2(n_483), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_860), .Y(n_920) );
OAI22xp33_ASAP7_75t_L g921 ( .A1(n_822), .A2(n_468), .B1(n_480), .B2(n_447), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g922 ( .A1(n_792), .A2(n_404), .B1(n_405), .B2(n_401), .C(n_373), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_882), .A2(n_483), .B1(n_406), .B2(n_412), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_882), .A2(n_407), .B1(n_420), .B2(n_413), .Y(n_924) );
AOI222xp33_ASAP7_75t_L g925 ( .A1(n_826), .A2(n_484), .B1(n_423), .B2(n_481), .C1(n_426), .C2(n_427), .Y(n_925) );
OAI22xp33_ASAP7_75t_L g926 ( .A1(n_818), .A2(n_480), .B1(n_749), .B2(n_739), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_785), .Y(n_927) );
INVxp67_ASAP7_75t_L g928 ( .A(n_832), .Y(n_928) );
AOI21xp5_ASAP7_75t_L g929 ( .A1(n_796), .A2(n_689), .B(n_657), .Y(n_929) );
AOI22xp5_ASAP7_75t_SL g930 ( .A1(n_789), .A2(n_741), .B1(n_437), .B2(n_438), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_871), .A2(n_695), .B1(n_689), .B2(n_739), .Y(n_931) );
OR2x2_ASAP7_75t_L g932 ( .A(n_766), .B(n_12), .Y(n_932) );
AOI22xp5_ASAP7_75t_SL g933 ( .A1(n_774), .A2(n_448), .B1(n_451), .B2(n_434), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_790), .Y(n_934) );
OAI221xp5_ASAP7_75t_L g935 ( .A1(n_837), .A2(n_750), .B1(n_493), .B2(n_467), .C(n_492), .Y(n_935) );
BUFx2_ASAP7_75t_L g936 ( .A(n_836), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_774), .A2(n_695), .B1(n_689), .B2(n_749), .Y(n_937) );
OAI221xp5_ASAP7_75t_L g938 ( .A1(n_837), .A2(n_488), .B1(n_482), .B2(n_475), .C(n_453), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_878), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_875), .A2(n_471), .B1(n_459), .B2(n_461), .Y(n_940) );
INVx2_ASAP7_75t_L g941 ( .A(n_883), .Y(n_941) );
INVx3_ASAP7_75t_L g942 ( .A(n_780), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_794), .A2(n_695), .B1(n_689), .B2(n_763), .Y(n_943) );
AO21x2_ASAP7_75t_L g944 ( .A1(n_776), .A2(n_504), .B(n_496), .Y(n_944) );
AO21x2_ASAP7_75t_L g945 ( .A1(n_814), .A2(n_504), .B(n_496), .Y(n_945) );
OAI211xp5_ASAP7_75t_SL g946 ( .A1(n_856), .A2(n_498), .B(n_461), .C(n_491), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_793), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_840), .B(n_13), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_798), .B(n_695), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_804), .Y(n_950) );
OAI22xp33_ASAP7_75t_L g951 ( .A1(n_832), .A2(n_763), .B1(n_757), .B2(n_491), .Y(n_951) );
OAI21x1_ASAP7_75t_L g952 ( .A1(n_814), .A2(n_504), .B(n_496), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_791), .A2(n_757), .B1(n_443), .B2(n_403), .Y(n_953) );
AOI21xp5_ASAP7_75t_L g954 ( .A1(n_890), .A2(n_757), .B(n_556), .Y(n_954) );
AOI21xp5_ASAP7_75t_L g955 ( .A1(n_890), .A2(n_556), .B(n_545), .Y(n_955) );
AO221x2_ASAP7_75t_L g956 ( .A1(n_889), .A2(n_14), .B1(n_15), .B2(n_16), .C(n_17), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_813), .B(n_14), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_854), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_844), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_832), .B(n_15), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_881), .A2(n_521), .B1(n_513), .B2(n_507), .Y(n_961) );
AOI22xp33_ASAP7_75t_SL g962 ( .A1(n_780), .A2(n_513), .B1(n_529), .B2(n_507), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_854), .Y(n_963) );
OR2x2_ASAP7_75t_L g964 ( .A(n_827), .B(n_16), .Y(n_964) );
OAI221xp5_ASAP7_75t_L g965 ( .A1(n_867), .A2(n_887), .B1(n_833), .B2(n_828), .C(n_863), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_825), .A2(n_521), .B1(n_513), .B2(n_507), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_791), .A2(n_521), .B1(n_513), .B2(n_507), .Y(n_967) );
OAI221xp5_ASAP7_75t_L g968 ( .A1(n_874), .A2(n_507), .B1(n_513), .B2(n_529), .C(n_556), .Y(n_968) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_868), .Y(n_969) );
OAI221xp5_ASAP7_75t_L g970 ( .A1(n_851), .A2(n_513), .B1(n_529), .B2(n_564), .C(n_561), .Y(n_970) );
INVx2_ASAP7_75t_L g971 ( .A(n_854), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_808), .A2(n_529), .B1(n_513), .B2(n_537), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_799), .A2(n_529), .B1(n_21), .B2(n_17), .Y(n_973) );
CKINVDCx8_ASAP7_75t_R g974 ( .A(n_768), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_844), .Y(n_975) );
AO21x2_ASAP7_75t_L g976 ( .A1(n_824), .A2(n_545), .B(n_537), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_799), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_839), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_808), .A2(n_529), .B1(n_547), .B2(n_545), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_845), .Y(n_980) );
NOR2xp33_ASAP7_75t_L g981 ( .A(n_829), .B(n_18), .Y(n_981) );
INVx2_ASAP7_75t_SL g982 ( .A(n_868), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_884), .Y(n_983) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_786), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_884), .Y(n_985) );
OAI211xp5_ASAP7_75t_L g986 ( .A1(n_779), .A2(n_529), .B(n_559), .C(n_547), .Y(n_986) );
INVx2_ASAP7_75t_L g987 ( .A(n_884), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_876), .A2(n_547), .B1(n_561), .B2(n_559), .Y(n_988) );
OAI22xp33_ASAP7_75t_L g989 ( .A1(n_820), .A2(n_23), .B1(n_21), .B2(n_22), .Y(n_989) );
INVx2_ASAP7_75t_L g990 ( .A(n_786), .Y(n_990) );
OAI221xp5_ASAP7_75t_L g991 ( .A1(n_861), .A2(n_564), .B1(n_561), .B2(n_559), .C(n_572), .Y(n_991) );
AOI22xp5_ASAP7_75t_L g992 ( .A1(n_872), .A2(n_564), .B1(n_554), .B2(n_540), .Y(n_992) );
AOI322xp5_ASAP7_75t_L g993 ( .A1(n_810), .A2(n_22), .A3(n_23), .B1(n_24), .B2(n_25), .C1(n_26), .C2(n_27), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_885), .A2(n_554), .B1(n_572), .B2(n_540), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_885), .A2(n_554), .B1(n_572), .B2(n_540), .Y(n_995) );
BUFx6f_ASAP7_75t_L g996 ( .A(n_869), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_787), .B(n_25), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_852), .A2(n_554), .B1(n_572), .B2(n_540), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_787), .B(n_26), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_858), .A2(n_554), .B1(n_572), .B2(n_540), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_862), .A2(n_554), .B1(n_572), .B2(n_540), .Y(n_1001) );
AOI222xp33_ASAP7_75t_L g1002 ( .A1(n_889), .A2(n_27), .B1(n_28), .B2(n_29), .C1(n_30), .C2(n_31), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_797), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_797), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_788), .B(n_29), .Y(n_1005) );
OAI21x1_ASAP7_75t_L g1006 ( .A1(n_865), .A2(n_554), .B(n_540), .Y(n_1006) );
AO21x2_ASAP7_75t_L g1007 ( .A1(n_880), .A2(n_554), .B(n_540), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_801), .A2(n_572), .B1(n_33), .B2(n_31), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_807), .A2(n_34), .B1(n_32), .B2(n_33), .Y(n_1009) );
OAI21x1_ASAP7_75t_L g1010 ( .A1(n_821), .A2(n_572), .B(n_113), .Y(n_1010) );
AO31x2_ASAP7_75t_L g1011 ( .A1(n_834), .A2(n_39), .A3(n_37), .B(n_38), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g1012 ( .A(n_782), .Y(n_1012) );
BUFx4f_ASAP7_75t_SL g1013 ( .A(n_817), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_801), .A2(n_39), .B1(n_37), .B2(n_38), .Y(n_1014) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_772), .B(n_40), .Y(n_1015) );
OAI31xp33_ASAP7_75t_L g1016 ( .A1(n_908), .A2(n_829), .A3(n_795), .B(n_772), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_977), .A2(n_802), .B1(n_809), .B2(n_806), .Y(n_1017) );
OR2x2_ASAP7_75t_L g1018 ( .A(n_964), .B(n_795), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_984), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_898), .B(n_816), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_901), .A2(n_771), .B1(n_812), .B2(n_784), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_911), .Y(n_1022) );
OAI22xp33_ASAP7_75t_L g1023 ( .A1(n_965), .A2(n_817), .B1(n_873), .B2(n_800), .Y(n_1023) );
INVx2_ASAP7_75t_L g1024 ( .A(n_941), .Y(n_1024) );
AOI322xp5_ASAP7_75t_L g1025 ( .A1(n_960), .A2(n_40), .A3(n_41), .B1(n_42), .B2(n_43), .C1(n_44), .C2(n_45), .Y(n_1025) );
OAI33xp33_ASAP7_75t_L g1026 ( .A1(n_989), .A2(n_773), .A3(n_811), .B1(n_44), .B2(n_45), .B3(n_46), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_895), .B(n_812), .Y(n_1027) );
OAI211xp5_ASAP7_75t_L g1028 ( .A1(n_1002), .A2(n_870), .B(n_843), .C(n_859), .Y(n_1028) );
INVx2_ASAP7_75t_L g1029 ( .A(n_941), .Y(n_1029) );
OA21x2_ASAP7_75t_L g1030 ( .A1(n_929), .A2(n_850), .B(n_838), .Y(n_1030) );
BUFx3_ASAP7_75t_L g1031 ( .A(n_905), .Y(n_1031) );
INVx3_ASAP7_75t_L g1032 ( .A(n_996), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_891), .Y(n_1033) );
OAI33xp33_ASAP7_75t_L g1034 ( .A1(n_1009), .A2(n_42), .A3(n_43), .B1(n_47), .B2(n_48), .B3(n_49), .Y(n_1034) );
INVx3_ASAP7_75t_SL g1035 ( .A(n_1012), .Y(n_1035) );
NOR3xp33_ASAP7_75t_L g1036 ( .A(n_938), .B(n_843), .C(n_800), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_933), .B(n_842), .Y(n_1037) );
AOI221xp5_ASAP7_75t_L g1038 ( .A1(n_922), .A2(n_864), .B1(n_846), .B2(n_815), .C(n_784), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_912), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_912), .Y(n_1040) );
AOI22xp33_ASAP7_75t_SL g1041 ( .A1(n_956), .A2(n_771), .B1(n_853), .B2(n_877), .Y(n_1041) );
AND2x4_ASAP7_75t_L g1042 ( .A(n_959), .B(n_849), .Y(n_1042) );
AOI21xp5_ASAP7_75t_L g1043 ( .A1(n_975), .A2(n_869), .B(n_848), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_950), .B(n_842), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_927), .Y(n_1045) );
INVx2_ASAP7_75t_L g1046 ( .A(n_914), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_950), .B(n_834), .Y(n_1047) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_924), .A2(n_831), .B1(n_846), .B2(n_879), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g1049 ( .A1(n_981), .A2(n_771), .B1(n_830), .B2(n_853), .Y(n_1049) );
OAI221xp5_ASAP7_75t_L g1050 ( .A1(n_924), .A2(n_879), .B1(n_841), .B2(n_771), .C(n_834), .Y(n_1050) );
INVx2_ASAP7_75t_L g1051 ( .A(n_914), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_934), .B(n_830), .Y(n_1052) );
AOI222xp33_ASAP7_75t_L g1053 ( .A1(n_1013), .A2(n_849), .B1(n_853), .B2(n_50), .C1(n_51), .C2(n_52), .Y(n_1053) );
AND2x4_ASAP7_75t_L g1054 ( .A(n_990), .B(n_849), .Y(n_1054) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_947), .A2(n_841), .B1(n_48), .B2(n_52), .C(n_53), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_920), .Y(n_1056) );
OA21x2_ASAP7_75t_L g1057 ( .A1(n_952), .A2(n_853), .B(n_114), .Y(n_1057) );
INVx2_ASAP7_75t_SL g1058 ( .A(n_936), .Y(n_1058) );
NAND3xp33_ASAP7_75t_L g1059 ( .A(n_993), .B(n_576), .C(n_47), .Y(n_1059) );
NAND4xp25_ASAP7_75t_L g1060 ( .A(n_915), .B(n_53), .C(n_54), .D(n_56), .Y(n_1060) );
INVx3_ASAP7_75t_L g1061 ( .A(n_996), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_978), .B(n_54), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_980), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_956), .B(n_57), .Y(n_1064) );
OAI31xp33_ASAP7_75t_SL g1065 ( .A1(n_981), .A2(n_57), .A3(n_58), .B(n_60), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_923), .A2(n_58), .B1(n_61), .B2(n_62), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_956), .A2(n_576), .B1(n_63), .B2(n_66), .Y(n_1067) );
NOR2x1p5_ASAP7_75t_L g1068 ( .A(n_942), .B(n_62), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1015), .B(n_66), .Y(n_1069) );
AOI31xp33_ASAP7_75t_L g1070 ( .A1(n_930), .A2(n_67), .A3(n_68), .B(n_69), .Y(n_1070) );
NAND3xp33_ASAP7_75t_L g1071 ( .A(n_925), .B(n_576), .C(n_67), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_893), .Y(n_1072) );
NOR2x1_ASAP7_75t_L g1073 ( .A(n_1012), .B(n_68), .Y(n_1073) );
AOI31xp67_ASAP7_75t_L g1074 ( .A1(n_970), .A2(n_963), .A3(n_971), .B(n_958), .Y(n_1074) );
NAND5xp2_ASAP7_75t_SL g1075 ( .A(n_1014), .B(n_70), .C(n_71), .D(n_72), .E(n_73), .Y(n_1075) );
CKINVDCx9p33_ASAP7_75t_R g1076 ( .A(n_974), .Y(n_1076) );
INVx2_ASAP7_75t_SL g1077 ( .A(n_969), .Y(n_1077) );
AO21x2_ASAP7_75t_L g1078 ( .A1(n_944), .A2(n_945), .B(n_904), .Y(n_1078) );
AOI22xp5_ASAP7_75t_L g1079 ( .A1(n_928), .A2(n_71), .B1(n_74), .B2(n_75), .Y(n_1079) );
BUFx6f_ASAP7_75t_L g1080 ( .A(n_996), .Y(n_1080) );
OAI211xp5_ASAP7_75t_L g1081 ( .A1(n_1014), .A2(n_576), .B(n_75), .C(n_76), .Y(n_1081) );
OAI21xp33_ASAP7_75t_L g1082 ( .A1(n_1008), .A2(n_74), .B(n_76), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1015), .B(n_77), .Y(n_1083) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_923), .A2(n_77), .B1(n_78), .B2(n_79), .Y(n_1084) );
OAI221xp5_ASAP7_75t_L g1085 ( .A1(n_896), .A2(n_79), .B1(n_80), .B2(n_81), .C(n_82), .Y(n_1085) );
OR2x6_ASAP7_75t_L g1086 ( .A(n_982), .B(n_81), .Y(n_1086) );
AOI222xp33_ASAP7_75t_L g1087 ( .A1(n_903), .A2(n_83), .B1(n_84), .B2(n_85), .C1(n_86), .C2(n_88), .Y(n_1087) );
INVx2_ASAP7_75t_L g1088 ( .A(n_920), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_1015), .A2(n_576), .B1(n_88), .B2(n_89), .Y(n_1089) );
AOI221x1_ASAP7_75t_SL g1090 ( .A1(n_957), .A2(n_84), .B1(n_89), .B2(n_90), .C(n_91), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_939), .B(n_90), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_935), .A2(n_576), .B1(n_93), .B2(n_94), .Y(n_1092) );
INVx2_ASAP7_75t_L g1093 ( .A(n_939), .Y(n_1093) );
OA21x2_ASAP7_75t_L g1094 ( .A1(n_1010), .A2(n_899), .B(n_900), .Y(n_1094) );
OAI22xp5_ASAP7_75t_SL g1095 ( .A1(n_907), .A2(n_942), .B1(n_1008), .B2(n_932), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_948), .Y(n_1096) );
OAI222xp33_ASAP7_75t_L g1097 ( .A1(n_973), .A2(n_91), .B1(n_95), .B2(n_96), .C1(n_97), .C2(n_98), .Y(n_1097) );
AOI21xp5_ASAP7_75t_L g1098 ( .A1(n_900), .A2(n_576), .B(n_115), .Y(n_1098) );
OAI21xp33_ASAP7_75t_L g1099 ( .A1(n_940), .A2(n_99), .B(n_102), .Y(n_1099) );
OAI222xp33_ASAP7_75t_L g1100 ( .A1(n_909), .A2(n_99), .B1(n_102), .B2(n_103), .C1(n_104), .C2(n_105), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g1101 ( .A1(n_892), .A2(n_105), .B1(n_106), .B2(n_107), .C(n_108), .Y(n_1101) );
NAND3xp33_ASAP7_75t_SL g1102 ( .A(n_897), .B(n_106), .C(n_107), .Y(n_1102) );
AOI33xp33_ASAP7_75t_L g1103 ( .A1(n_940), .A2(n_110), .A3(n_116), .B1(n_117), .B2(n_121), .B3(n_122), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_997), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_990), .B(n_123), .Y(n_1105) );
AOI221xp5_ASAP7_75t_L g1106 ( .A1(n_946), .A2(n_576), .B1(n_126), .B2(n_127), .C(n_128), .Y(n_1106) );
NAND3xp33_ASAP7_75t_L g1107 ( .A(n_894), .B(n_124), .C(n_129), .Y(n_1107) );
OAI31xp33_ASAP7_75t_SL g1108 ( .A1(n_951), .A2(n_133), .A3(n_135), .B(n_136), .Y(n_1108) );
AOI22xp5_ASAP7_75t_L g1109 ( .A1(n_921), .A2(n_138), .B1(n_140), .B2(n_141), .Y(n_1109) );
OAI211xp5_ASAP7_75t_L g1110 ( .A1(n_999), .A2(n_145), .B(n_146), .C(n_150), .Y(n_1110) );
INVx2_ASAP7_75t_SL g1111 ( .A(n_996), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1005), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1011), .Y(n_1113) );
OAI21xp5_ASAP7_75t_L g1114 ( .A1(n_892), .A2(n_151), .B(n_152), .Y(n_1114) );
BUFx5_ASAP7_75t_L g1115 ( .A(n_1003), .Y(n_1115) );
NOR2x1_ASAP7_75t_SL g1116 ( .A(n_906), .B(n_154), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1011), .Y(n_1117) );
BUFx2_ASAP7_75t_L g1118 ( .A(n_1004), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_917), .B(n_155), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_902), .A2(n_156), .B1(n_157), .B2(n_158), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1011), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_902), .A2(n_159), .B1(n_160), .B2(n_162), .Y(n_1122) );
AOI21xp5_ASAP7_75t_L g1123 ( .A1(n_954), .A2(n_166), .B(n_168), .Y(n_1123) );
NAND3xp33_ASAP7_75t_L g1124 ( .A(n_966), .B(n_169), .C(n_171), .Y(n_1124) );
AOI22xp33_ASAP7_75t_SL g1125 ( .A1(n_953), .A2(n_172), .B1(n_174), .B2(n_177), .Y(n_1125) );
AOI31xp33_ASAP7_75t_L g1126 ( .A1(n_909), .A2(n_178), .A3(n_179), .B(n_180), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1011), .Y(n_1127) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_949), .Y(n_1128) );
INVx2_ASAP7_75t_L g1129 ( .A(n_945), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1027), .B(n_913), .Y(n_1130) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1024), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1063), .Y(n_1132) );
NAND2x1p5_ASAP7_75t_L g1133 ( .A(n_1031), .B(n_910), .Y(n_1133) );
OAI221xp5_ASAP7_75t_L g1134 ( .A1(n_1060), .A2(n_919), .B1(n_913), .B2(n_918), .C(n_961), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1033), .B(n_919), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1022), .Y(n_1136) );
OR2x2_ASAP7_75t_L g1137 ( .A(n_1018), .B(n_958), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1045), .Y(n_1138) );
OR2x2_ASAP7_75t_L g1139 ( .A(n_1019), .B(n_963), .Y(n_1139) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_1070), .A2(n_926), .B1(n_968), .B2(n_961), .C(n_966), .Y(n_1140) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1029), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1062), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1062), .Y(n_1143) );
OAI31xp33_ASAP7_75t_L g1144 ( .A1(n_1068), .A2(n_986), .A3(n_967), .B(n_943), .Y(n_1144) );
OAI222xp33_ASAP7_75t_L g1145 ( .A1(n_1041), .A2(n_1086), .B1(n_1064), .B2(n_1067), .C1(n_1037), .C2(n_1050), .Y(n_1145) );
BUFx2_ASAP7_75t_L g1146 ( .A(n_1080), .Y(n_1146) );
INVx3_ASAP7_75t_L g1147 ( .A(n_1080), .Y(n_1147) );
INVx2_ASAP7_75t_L g1148 ( .A(n_1039), .Y(n_1148) );
INVx8_ASAP7_75t_L g1149 ( .A(n_1086), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1072), .B(n_944), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1096), .B(n_918), .Y(n_1151) );
INVx1_ASAP7_75t_SL g1152 ( .A(n_1076), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1091), .Y(n_1153) );
BUFx2_ASAP7_75t_L g1154 ( .A(n_1080), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1069), .B(n_916), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_1126), .A2(n_916), .B1(n_994), .B2(n_995), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1091), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_1075), .A2(n_976), .B1(n_1007), .B2(n_931), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1052), .B(n_971), .Y(n_1159) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1052), .B(n_983), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1044), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1083), .B(n_983), .Y(n_1162) );
OAI221xp5_ASAP7_75t_L g1163 ( .A1(n_1065), .A2(n_995), .B1(n_994), .B2(n_992), .C(n_962), .Y(n_1163) );
AOI31xp33_ASAP7_75t_L g1164 ( .A1(n_1053), .A2(n_937), .A3(n_972), .B(n_1000), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1128), .B(n_985), .Y(n_1165) );
AOI221xp5_ASAP7_75t_L g1166 ( .A1(n_1070), .A2(n_972), .B1(n_988), .B2(n_955), .C(n_979), .Y(n_1166) );
BUFx3_ASAP7_75t_L g1167 ( .A(n_1032), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1077), .B(n_985), .Y(n_1168) );
INVx2_ASAP7_75t_L g1169 ( .A(n_1040), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1112), .B(n_987), .Y(n_1170) );
AOI22xp5_ASAP7_75t_L g1171 ( .A1(n_1053), .A2(n_976), .B1(n_1007), .B2(n_979), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1020), .B(n_987), .Y(n_1172) );
INVx4_ASAP7_75t_L g1173 ( .A(n_1042), .Y(n_1173) );
OR2x2_ASAP7_75t_L g1174 ( .A(n_1058), .B(n_998), .Y(n_1174) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_1046), .B(n_998), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1118), .Y(n_1176) );
AND2x2_ASAP7_75t_SL g1177 ( .A(n_1108), .B(n_1000), .Y(n_1177) );
NOR2xp33_ASAP7_75t_L g1178 ( .A(n_1102), .B(n_991), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1051), .B(n_1001), .Y(n_1179) );
AOI21x1_ASAP7_75t_L g1180 ( .A1(n_1113), .A2(n_1006), .B(n_1001), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1056), .B(n_988), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1088), .Y(n_1182) );
NOR3xp33_ASAP7_75t_SL g1183 ( .A(n_1023), .B(n_181), .C(n_182), .Y(n_1183) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1093), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1185 ( .A(n_1104), .B(n_185), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1086), .B(n_189), .Y(n_1186) );
AND2x2_ASAP7_75t_SL g1187 ( .A(n_1108), .B(n_190), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1115), .B(n_191), .Y(n_1188) );
NAND3xp33_ASAP7_75t_L g1189 ( .A(n_1065), .B(n_196), .C(n_197), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1047), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1047), .Y(n_1191) );
AOI33xp33_ASAP7_75t_L g1192 ( .A1(n_1055), .A2(n_198), .A3(n_199), .B1(n_200), .B2(n_203), .B3(n_207), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1087), .B(n_208), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1111), .B(n_209), .Y(n_1194) );
NAND3xp33_ASAP7_75t_L g1195 ( .A(n_1087), .B(n_211), .C(n_212), .Y(n_1195) );
AOI322xp5_ASAP7_75t_L g1196 ( .A1(n_1073), .A2(n_214), .A3(n_217), .B1(n_218), .B2(n_219), .C1(n_221), .C2(n_222), .Y(n_1196) );
NOR3xp33_ASAP7_75t_L g1197 ( .A(n_1026), .B(n_227), .C(n_230), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1090), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1032), .B(n_231), .Y(n_1199) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1061), .Y(n_1200) );
HB1xp67_ASAP7_75t_L g1201 ( .A(n_1129), .Y(n_1201) );
BUFx2_ASAP7_75t_L g1202 ( .A(n_1061), .Y(n_1202) );
INVxp67_ASAP7_75t_SL g1203 ( .A(n_1117), .Y(n_1203) );
AND2x4_ASAP7_75t_L g1204 ( .A(n_1042), .B(n_233), .Y(n_1204) );
AOI211xp5_ASAP7_75t_L g1205 ( .A1(n_1095), .A2(n_234), .B(n_236), .C(n_240), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1090), .Y(n_1206) );
INVx3_ASAP7_75t_L g1207 ( .A(n_1054), .Y(n_1207) );
NAND3xp33_ASAP7_75t_L g1208 ( .A(n_1025), .B(n_241), .C(n_242), .Y(n_1208) );
INVxp67_ASAP7_75t_L g1209 ( .A(n_1050), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1121), .Y(n_1210) );
NAND3xp33_ASAP7_75t_L g1211 ( .A(n_1055), .B(n_243), .C(n_244), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1021), .B(n_246), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1115), .B(n_247), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1127), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1105), .Y(n_1215) );
NAND3xp33_ASAP7_75t_L g1216 ( .A(n_1079), .B(n_249), .C(n_250), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1217 ( .A(n_1078), .Y(n_1217) );
OR2x2_ASAP7_75t_L g1218 ( .A(n_1066), .B(n_255), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1115), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1066), .B(n_259), .Y(n_1220) );
INVx2_ASAP7_75t_L g1221 ( .A(n_1078), .Y(n_1221) );
NAND4xp25_ASAP7_75t_L g1222 ( .A(n_1071), .B(n_260), .C(n_262), .D(n_266), .Y(n_1222) );
NOR2xp33_ASAP7_75t_L g1223 ( .A(n_1034), .B(n_267), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1115), .Y(n_1224) );
AOI221xp5_ASAP7_75t_L g1225 ( .A1(n_1084), .A2(n_268), .B1(n_270), .B2(n_273), .C(n_274), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1115), .Y(n_1226) );
AND2x4_ASAP7_75t_L g1227 ( .A(n_1054), .B(n_275), .Y(n_1227) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1084), .B(n_325), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g1229 ( .A(n_1101), .B(n_276), .Y(n_1229) );
INVxp67_ASAP7_75t_SL g1230 ( .A(n_1201), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1132), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1136), .Y(n_1232) );
NOR3xp33_ASAP7_75t_L g1233 ( .A(n_1195), .B(n_1101), .C(n_1097), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1138), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1176), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_1187), .A2(n_1082), .B1(n_1099), .B2(n_1085), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1190), .B(n_1094), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1161), .B(n_1016), .Y(n_1238) );
NAND2x1_ASAP7_75t_SL g1239 ( .A(n_1186), .B(n_1035), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1191), .B(n_1094), .Y(n_1240) );
AND2x4_ASAP7_75t_L g1241 ( .A(n_1210), .B(n_1116), .Y(n_1241) );
NAND3xp33_ASAP7_75t_L g1242 ( .A(n_1198), .B(n_1059), .C(n_1089), .Y(n_1242) );
NOR3xp33_ASAP7_75t_SL g1243 ( .A(n_1145), .B(n_1100), .C(n_1081), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1214), .B(n_1030), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1245 ( .A(n_1165), .B(n_1049), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1182), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1165), .Y(n_1247) );
OAI21xp33_ASAP7_75t_L g1248 ( .A1(n_1187), .A2(n_1126), .B(n_1103), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1209), .B(n_1030), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1209), .B(n_1119), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1201), .B(n_1017), .Y(n_1251) );
NAND5xp2_ASAP7_75t_SL g1252 ( .A(n_1177), .B(n_1085), .C(n_1028), .D(n_1092), .E(n_1110), .Y(n_1252) );
INVx3_ASAP7_75t_L g1253 ( .A(n_1219), .Y(n_1253) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1148), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1172), .B(n_1017), .Y(n_1255) );
OR2x2_ASAP7_75t_L g1256 ( .A(n_1150), .B(n_1048), .Y(n_1256) );
INVxp67_ASAP7_75t_L g1257 ( .A(n_1168), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1150), .B(n_1048), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1206), .B(n_1038), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1142), .B(n_1043), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1203), .B(n_1114), .Y(n_1261) );
AOI211xp5_ASAP7_75t_L g1262 ( .A1(n_1145), .A2(n_1036), .B(n_1114), .C(n_1106), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1170), .Y(n_1263) );
AOI221xp5_ASAP7_75t_L g1264 ( .A1(n_1143), .A2(n_1106), .B1(n_1123), .B2(n_1098), .C(n_1122), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1137), .Y(n_1265) );
OAI211xp5_ASAP7_75t_SL g1266 ( .A1(n_1152), .A2(n_1109), .B(n_1125), .C(n_1120), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1131), .Y(n_1267) );
INVx1_ASAP7_75t_SL g1268 ( .A(n_1149), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1151), .B(n_1057), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1141), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1203), .B(n_1057), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1159), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1160), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1139), .Y(n_1274) );
OA21x2_ASAP7_75t_L g1275 ( .A1(n_1221), .A2(n_1074), .B(n_1107), .Y(n_1275) );
NAND3x1_ASAP7_75t_SL g1276 ( .A(n_1144), .B(n_1124), .C(n_278), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1169), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1184), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1153), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1157), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1224), .B(n_277), .Y(n_1281) );
AOI221xp5_ASAP7_75t_L g1282 ( .A1(n_1149), .A2(n_279), .B1(n_280), .B2(n_281), .C(n_283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1174), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1215), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1135), .B(n_286), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1226), .B(n_287), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1221), .B(n_288), .Y(n_1287) );
INVx2_ASAP7_75t_L g1288 ( .A(n_1180), .Y(n_1288) );
OR2x2_ASAP7_75t_L g1289 ( .A(n_1155), .B(n_289), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1202), .Y(n_1290) );
OAI221xp5_ASAP7_75t_L g1291 ( .A1(n_1133), .A2(n_290), .B1(n_291), .B2(n_299), .C(n_301), .Y(n_1291) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1217), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1217), .B(n_302), .Y(n_1293) );
AND2x4_ASAP7_75t_L g1294 ( .A(n_1207), .B(n_303), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1162), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1200), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1130), .B(n_305), .Y(n_1297) );
INVx2_ASAP7_75t_L g1298 ( .A(n_1175), .Y(n_1298) );
NOR2xp33_ASAP7_75t_L g1299 ( .A(n_1133), .B(n_1149), .Y(n_1299) );
INVx2_ASAP7_75t_L g1300 ( .A(n_1179), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1207), .B(n_307), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1177), .B(n_308), .Y(n_1302) );
AND2x4_ASAP7_75t_L g1303 ( .A(n_1173), .B(n_309), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1173), .B(n_311), .Y(n_1304) );
NAND3xp33_ASAP7_75t_SL g1305 ( .A(n_1205), .B(n_312), .C(n_313), .Y(n_1305) );
INVx4_ASAP7_75t_L g1306 ( .A(n_1204), .Y(n_1306) );
NOR2xp33_ASAP7_75t_SL g1307 ( .A(n_1204), .B(n_316), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1249), .B(n_1171), .Y(n_1308) );
AOI21xp5_ASAP7_75t_L g1309 ( .A1(n_1248), .A2(n_1156), .B(n_1164), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1283), .B(n_1223), .Y(n_1310) );
NOR2xp33_ASAP7_75t_SL g1311 ( .A(n_1306), .B(n_1156), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1249), .B(n_1158), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1231), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1247), .B(n_1223), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1244), .B(n_1158), .Y(n_1315) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1238), .B(n_1189), .Y(n_1316) );
BUFx3_ASAP7_75t_L g1317 ( .A(n_1306), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1274), .B(n_1193), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1232), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1234), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1272), .B(n_1197), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1284), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1235), .Y(n_1323) );
INVxp67_ASAP7_75t_SL g1324 ( .A(n_1230), .Y(n_1324) );
INVxp67_ASAP7_75t_L g1325 ( .A(n_1299), .Y(n_1325) );
OAI21xp5_ASAP7_75t_SL g1326 ( .A1(n_1299), .A2(n_1222), .B(n_1196), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1244), .B(n_1197), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1328 ( .A(n_1273), .B(n_1265), .Y(n_1328) );
NAND4xp25_ASAP7_75t_L g1329 ( .A(n_1262), .B(n_1208), .C(n_1229), .D(n_1225), .Y(n_1329) );
INVxp67_ASAP7_75t_L g1330 ( .A(n_1307), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1251), .B(n_1298), .Y(n_1331) );
NAND4xp25_ASAP7_75t_L g1332 ( .A(n_1236), .B(n_1229), .C(n_1225), .D(n_1140), .Y(n_1332) );
OAI21xp5_ASAP7_75t_L g1333 ( .A1(n_1243), .A2(n_1183), .B(n_1211), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1279), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1251), .B(n_1146), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1280), .Y(n_1336) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_1259), .B(n_1185), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1246), .Y(n_1338) );
NAND4xp25_ASAP7_75t_L g1339 ( .A(n_1236), .B(n_1140), .C(n_1178), .D(n_1166), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1263), .B(n_1181), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1298), .B(n_1154), .Y(n_1341) );
NOR2xp33_ASAP7_75t_L g1342 ( .A(n_1257), .B(n_1260), .Y(n_1342) );
NOR2xp33_ASAP7_75t_L g1343 ( .A(n_1242), .B(n_1212), .Y(n_1343) );
NAND2x1p5_ASAP7_75t_L g1344 ( .A(n_1306), .B(n_1227), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1295), .Y(n_1345) );
NAND2xp67_ASAP7_75t_L g1346 ( .A(n_1302), .B(n_1220), .Y(n_1346) );
HB1xp67_ASAP7_75t_L g1347 ( .A(n_1254), .Y(n_1347) );
XOR2xp5_ASAP7_75t_L g1348 ( .A(n_1268), .B(n_1227), .Y(n_1348) );
NAND2xp5_ASAP7_75t_SL g1349 ( .A(n_1241), .B(n_1183), .Y(n_1349) );
OR2x2_ASAP7_75t_L g1350 ( .A(n_1300), .B(n_1167), .Y(n_1350) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1254), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1300), .B(n_1167), .Y(n_1352) );
OR2x2_ASAP7_75t_L g1353 ( .A(n_1245), .B(n_1147), .Y(n_1353) );
NAND3xp33_ASAP7_75t_L g1354 ( .A(n_1233), .B(n_1192), .C(n_1178), .Y(n_1354) );
INVx1_ASAP7_75t_SL g1355 ( .A(n_1239), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1237), .B(n_1147), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1357 ( .A(n_1267), .B(n_1213), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_1252), .A2(n_1134), .B1(n_1218), .B2(n_1228), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1313), .Y(n_1359) );
INVx2_ASAP7_75t_SL g1360 ( .A(n_1317), .Y(n_1360) );
NOR2xp33_ASAP7_75t_L g1361 ( .A(n_1339), .B(n_1290), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1319), .Y(n_1362) );
AOI221xp5_ASAP7_75t_L g1363 ( .A1(n_1309), .A2(n_1302), .B1(n_1250), .B2(n_1255), .C(n_1296), .Y(n_1363) );
OAI22xp33_ASAP7_75t_SL g1364 ( .A1(n_1311), .A2(n_1303), .B1(n_1258), .B2(n_1256), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1320), .Y(n_1365) );
OAI31xp33_ASAP7_75t_L g1366 ( .A1(n_1354), .A2(n_1266), .A3(n_1291), .B(n_1250), .Y(n_1366) );
OAI211xp5_ASAP7_75t_SL g1367 ( .A1(n_1333), .A2(n_1282), .B(n_1285), .C(n_1297), .Y(n_1367) );
INVxp67_ASAP7_75t_L g1368 ( .A(n_1342), .Y(n_1368) );
INVxp67_ASAP7_75t_L g1369 ( .A(n_1342), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1331), .B(n_1237), .Y(n_1370) );
AO22x2_ASAP7_75t_L g1371 ( .A1(n_1323), .A2(n_1253), .B1(n_1256), .B2(n_1258), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1331), .B(n_1240), .Y(n_1372) );
OR2x2_ASAP7_75t_L g1373 ( .A(n_1328), .B(n_1292), .Y(n_1373) );
O2A1O1Ixp33_ASAP7_75t_L g1374 ( .A1(n_1326), .A2(n_1332), .B(n_1329), .C(n_1349), .Y(n_1374) );
NAND4xp25_ASAP7_75t_L g1375 ( .A(n_1358), .B(n_1289), .C(n_1255), .D(n_1261), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1308), .B(n_1278), .Y(n_1376) );
OAI21xp5_ASAP7_75t_L g1377 ( .A1(n_1349), .A2(n_1305), .B(n_1303), .Y(n_1377) );
OAI21xp33_ASAP7_75t_L g1378 ( .A1(n_1343), .A2(n_1261), .B(n_1269), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1338), .Y(n_1379) );
NAND2xp5_ASAP7_75t_L g1380 ( .A(n_1308), .B(n_1270), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1322), .Y(n_1381) );
INVx2_ASAP7_75t_L g1382 ( .A(n_1351), .Y(n_1382) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1334), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_1345), .B(n_1277), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1315), .B(n_1240), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1315), .B(n_1292), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1335), .B(n_1271), .Y(n_1387) );
INVx1_ASAP7_75t_SL g1388 ( .A(n_1348), .Y(n_1388) );
NOR2xp33_ASAP7_75t_L g1389 ( .A(n_1343), .B(n_1241), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1336), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1312), .B(n_1253), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1392 ( .A(n_1312), .B(n_1253), .Y(n_1392) );
INVxp67_ASAP7_75t_L g1393 ( .A(n_1324), .Y(n_1393) );
AOI22xp33_ASAP7_75t_L g1394 ( .A1(n_1316), .A2(n_1241), .B1(n_1134), .B2(n_1303), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1347), .Y(n_1395) );
AOI221xp5_ASAP7_75t_L g1396 ( .A1(n_1337), .A2(n_1358), .B1(n_1316), .B2(n_1318), .C(n_1325), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1340), .B(n_1293), .Y(n_1397) );
AOI22xp33_ASAP7_75t_L g1398 ( .A1(n_1327), .A2(n_1294), .B1(n_1216), .B2(n_1293), .Y(n_1398) );
OA21x2_ASAP7_75t_L g1399 ( .A1(n_1321), .A2(n_1288), .B(n_1271), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1335), .B(n_1288), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1310), .B(n_1287), .Y(n_1401) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_1344), .A2(n_1294), .B1(n_1304), .B2(n_1301), .Y(n_1402) );
AOI22xp5_ASAP7_75t_L g1403 ( .A1(n_1337), .A2(n_1301), .B1(n_1294), .B2(n_1264), .Y(n_1403) );
XOR2x2_ASAP7_75t_L g1404 ( .A(n_1344), .B(n_1276), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1356), .B(n_1275), .Y(n_1405) );
A2O1A1Ixp33_ASAP7_75t_SL g1406 ( .A1(n_1330), .A2(n_1163), .B(n_1286), .C(n_1281), .Y(n_1406) );
AOI22xp5_ASAP7_75t_L g1407 ( .A1(n_1355), .A2(n_1286), .B1(n_1281), .B2(n_1166), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1356), .B(n_1341), .Y(n_1408) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1352), .Y(n_1409) );
OAI21xp5_ASAP7_75t_SL g1410 ( .A1(n_1327), .A2(n_1163), .B(n_1213), .Y(n_1410) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1341), .Y(n_1411) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1350), .Y(n_1412) );
AOI211xp5_ASAP7_75t_L g1413 ( .A1(n_1374), .A2(n_1364), .B(n_1366), .C(n_1396), .Y(n_1413) );
BUFx2_ASAP7_75t_L g1414 ( .A(n_1360), .Y(n_1414) );
INVx2_ASAP7_75t_L g1415 ( .A(n_1382), .Y(n_1415) );
NOR3xp33_ASAP7_75t_L g1416 ( .A(n_1361), .B(n_1276), .C(n_1367), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1373), .Y(n_1417) );
NAND3xp33_ASAP7_75t_L g1418 ( .A(n_1361), .B(n_1377), .C(n_1394), .Y(n_1418) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_1375), .A2(n_1368), .B1(n_1369), .B2(n_1363), .Y(n_1419) );
OAI22xp5_ASAP7_75t_L g1420 ( .A1(n_1360), .A2(n_1389), .B1(n_1407), .B2(n_1393), .Y(n_1420) );
AOI221xp5_ASAP7_75t_L g1421 ( .A1(n_1371), .A2(n_1378), .B1(n_1410), .B2(n_1389), .C(n_1409), .Y(n_1421) );
HB1xp67_ASAP7_75t_L g1422 ( .A(n_1399), .Y(n_1422) );
NAND2xp5_ASAP7_75t_L g1423 ( .A(n_1371), .B(n_1399), .Y(n_1423) );
AOI222xp33_ASAP7_75t_L g1424 ( .A1(n_1371), .A2(n_1388), .B1(n_1405), .B2(n_1406), .C1(n_1392), .C2(n_1391), .Y(n_1424) );
XNOR2x1_ASAP7_75t_L g1425 ( .A(n_1404), .B(n_1403), .Y(n_1425) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1381), .Y(n_1426) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1383), .Y(n_1427) );
OAI211xp5_ASAP7_75t_L g1428 ( .A1(n_1413), .A2(n_1424), .B(n_1421), .C(n_1416), .Y(n_1428) );
OA22x2_ASAP7_75t_L g1429 ( .A1(n_1420), .A2(n_1402), .B1(n_1405), .B2(n_1362), .Y(n_1429) );
NAND4xp75_ASAP7_75t_L g1430 ( .A(n_1423), .B(n_1399), .C(n_1404), .D(n_1314), .Y(n_1430) );
AOI21xp33_ASAP7_75t_SL g1431 ( .A1(n_1425), .A2(n_1398), .B(n_1406), .Y(n_1431) );
O2A1O1Ixp33_ASAP7_75t_L g1432 ( .A1(n_1418), .A2(n_1359), .B(n_1365), .C(n_1379), .Y(n_1432) );
OAI211xp5_ASAP7_75t_SL g1433 ( .A1(n_1416), .A2(n_1376), .B(n_1380), .C(n_1390), .Y(n_1433) );
OAI22xp5_ASAP7_75t_L g1434 ( .A1(n_1419), .A2(n_1317), .B1(n_1412), .B2(n_1385), .Y(n_1434) );
NAND5xp2_ASAP7_75t_L g1435 ( .A(n_1419), .B(n_1401), .C(n_1346), .D(n_1397), .E(n_1400), .Y(n_1435) );
AOI211xp5_ASAP7_75t_L g1436 ( .A1(n_1422), .A2(n_1353), .B(n_1386), .C(n_1400), .Y(n_1436) );
NAND3xp33_ASAP7_75t_L g1437 ( .A(n_1428), .B(n_1414), .C(n_1426), .Y(n_1437) );
CKINVDCx20_ASAP7_75t_R g1438 ( .A(n_1434), .Y(n_1438) );
AOI221xp5_ASAP7_75t_L g1439 ( .A1(n_1431), .A2(n_1427), .B1(n_1417), .B2(n_1395), .C(n_1384), .Y(n_1439) );
OAI211xp5_ASAP7_75t_SL g1440 ( .A1(n_1432), .A2(n_1192), .B(n_1412), .C(n_1415), .Y(n_1440) );
XNOR2xp5_ASAP7_75t_L g1441 ( .A(n_1430), .B(n_1387), .Y(n_1441) );
HB1xp67_ASAP7_75t_L g1442 ( .A(n_1429), .Y(n_1442) );
OAI221xp5_ASAP7_75t_L g1443 ( .A1(n_1442), .A2(n_1429), .B1(n_1433), .B2(n_1436), .C(n_1435), .Y(n_1443) );
XNOR2xp5_ASAP7_75t_SL g1444 ( .A(n_1441), .B(n_1411), .Y(n_1444) );
INVxp33_ASAP7_75t_SL g1445 ( .A(n_1437), .Y(n_1445) );
OAI211xp5_ASAP7_75t_SL g1446 ( .A1(n_1439), .A2(n_1188), .B(n_1194), .C(n_1357), .Y(n_1446) );
OAI21xp5_ASAP7_75t_L g1447 ( .A1(n_1438), .A2(n_1408), .B(n_1387), .Y(n_1447) );
INVx3_ASAP7_75t_SL g1448 ( .A(n_1445), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1447), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1444), .Y(n_1450) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1443), .Y(n_1451) );
OAI22x1_ASAP7_75t_L g1452 ( .A1(n_1448), .A2(n_1451), .B1(n_1450), .B2(n_1449), .Y(n_1452) );
INVx4_ASAP7_75t_L g1453 ( .A(n_1448), .Y(n_1453) );
BUFx3_ASAP7_75t_L g1454 ( .A(n_1453), .Y(n_1454) );
AOI222xp33_ASAP7_75t_L g1455 ( .A1(n_1452), .A2(n_1446), .B1(n_1440), .B2(n_1372), .C1(n_1370), .C2(n_1199), .Y(n_1455) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1454), .Y(n_1456) );
AOI21xp5_ASAP7_75t_L g1457 ( .A1(n_1456), .A2(n_1455), .B(n_1188), .Y(n_1457) );
endmodule