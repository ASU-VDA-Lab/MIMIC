module fake_jpeg_14508_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_49),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_28),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_51),
.A2(n_59),
.B(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_28),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_23),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_34),
.B1(n_36),
.B2(n_23),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_34),
.B1(n_20),
.B2(n_29),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_63),
.A2(n_50),
.B1(n_42),
.B2(n_43),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_26),
.B1(n_21),
.B2(n_34),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_38),
.B1(n_47),
.B2(n_45),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_66),
.B(n_36),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_39),
.B(n_28),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_41),
.C(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_70),
.B(n_84),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_77),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_18),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_73),
.B(n_76),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_41),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_74),
.Y(n_142)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_27),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_24),
.B1(n_33),
.B2(n_29),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_113),
.B1(n_114),
.B2(n_49),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_83),
.Y(n_116)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_33),
.B(n_20),
.C(n_24),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_55),
.B(n_27),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_20),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_R g115 ( 
.A(n_91),
.B(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_19),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_98),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_65),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_96),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_24),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_33),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_99),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_59),
.B(n_31),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_102),
.B(n_106),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_29),
.B(n_30),
.C(n_35),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_109),
.B1(n_48),
.B2(n_50),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_60),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_31),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_19),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_111),
.B(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_18),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_57),
.A2(n_38),
.B1(n_47),
.B2(n_45),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_57),
.A2(n_45),
.B1(n_44),
.B2(n_47),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_103),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_44),
.B1(n_26),
.B2(n_21),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_124),
.B1(n_133),
.B2(n_137),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_21),
.B1(n_26),
.B2(n_44),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_26),
.B1(n_21),
.B2(n_41),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_34),
.B1(n_23),
.B2(n_36),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_147),
.A2(n_149),
.B1(n_154),
.B2(n_86),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_130),
.B1(n_129),
.B2(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_76),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_77),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_152),
.B(n_157),
.Y(n_194)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_100),
.B1(n_70),
.B2(n_72),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_87),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_126),
.Y(n_158)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_159),
.B(n_161),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_74),
.C(n_81),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_173),
.C(n_86),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_97),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_74),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_125),
.B(n_80),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_164),
.B(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_98),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_91),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_171),
.Y(n_207)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_123),
.B(n_78),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_133),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_96),
.C(n_85),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_94),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_125),
.B1(n_115),
.B2(n_141),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_176),
.A2(n_182),
.B1(n_184),
.B2(n_189),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_115),
.B(n_120),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_191),
.B(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_128),
.B1(n_135),
.B2(n_136),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_183),
.B(n_198),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_135),
.B1(n_136),
.B2(n_117),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_137),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_204),
.C(n_158),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_163),
.A2(n_102),
.B1(n_119),
.B2(n_109),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_121),
.B(n_122),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_203),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_154),
.A2(n_139),
.B1(n_132),
.B2(n_131),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_196),
.A2(n_197),
.B(n_173),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_148),
.A2(n_139),
.B1(n_89),
.B2(n_104),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_205),
.B1(n_206),
.B2(n_50),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_132),
.B(n_82),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_150),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_92),
.C(n_144),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_147),
.A2(n_107),
.B1(n_71),
.B2(n_90),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_147),
.A2(n_71),
.B1(n_75),
.B2(n_105),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_207),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_223),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_155),
.Y(n_211)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_146),
.Y(n_215)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_166),
.Y(n_216)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_200),
.B(n_170),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_226),
.C(n_188),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_158),
.B1(n_167),
.B2(n_156),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_219),
.A2(n_224),
.B1(n_229),
.B2(n_236),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_180),
.A2(n_153),
.B(n_151),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_235),
.B(n_190),
.Y(n_254)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_171),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_144),
.B1(n_30),
.B2(n_35),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_181),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_95),
.C(n_48),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_185),
.A2(n_36),
.B1(n_99),
.B2(n_35),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_11),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_233),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_10),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_175),
.B(n_99),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_177),
.B(n_10),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_190),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_43),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_192),
.B1(n_30),
.B2(n_99),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_228),
.A2(n_187),
.B1(n_183),
.B2(n_199),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_219),
.B1(n_209),
.B2(n_211),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_248),
.C(n_256),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_188),
.C(n_199),
.Y(n_248)
);

OA21x2_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_206),
.B(n_189),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_210),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_255),
.B(n_229),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_175),
.C(n_205),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_192),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_261),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_43),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_217),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_268),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_266),
.A2(n_267),
.B1(n_270),
.B2(n_281),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_238),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_223),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_222),
.B1(n_208),
.B2(n_235),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_214),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_240),
.A2(n_222),
.B1(n_231),
.B2(n_220),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_277),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_235),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_241),
.Y(n_287)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_280),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_247),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_282),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_252),
.B(n_237),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_253),
.A2(n_236),
.B1(n_221),
.B2(n_213),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_255),
.B(n_212),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_242),
.C(n_248),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_286),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_256),
.C(n_261),
.Y(n_286)
);

XNOR2x1_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_281),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_254),
.C(n_245),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_297),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

AO221x1_ASAP7_75t_L g295 ( 
.A1(n_264),
.A2(n_262),
.B1(n_259),
.B2(n_251),
.C(n_246),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_291),
.B(n_296),
.Y(n_302)
);

OAI322xp33_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_266),
.A3(n_269),
.B1(n_272),
.B2(n_246),
.C1(n_270),
.C2(n_273),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_251),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_299),
.B(n_301),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_250),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_306),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_274),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_304),
.Y(n_323)
);

AO22x1_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_250),
.B1(n_224),
.B2(n_233),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_309),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_289),
.A2(n_257),
.B1(n_42),
.B2(n_9),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_42),
.B1(n_8),
.B2(n_9),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_310),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_298),
.A2(n_36),
.B1(n_7),
.B2(n_9),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_6),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_288),
.A2(n_6),
.B1(n_16),
.B2(n_15),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_314),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_285),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_314)
);

AOI211xp5_ASAP7_75t_L g319 ( 
.A1(n_308),
.A2(n_292),
.B(n_293),
.C(n_294),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_313),
.B1(n_309),
.B2(n_314),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_286),
.B(n_287),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_4),
.B(n_12),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_285),
.B1(n_5),
.B2(n_7),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_322),
.A2(n_325),
.B1(n_12),
.B2(n_1),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_17),
.C(n_5),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_324),
.B(n_0),
.Y(n_333)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_303),
.B(n_5),
.CI(n_15),
.CON(n_325),
.SN(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_310),
.C(n_305),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_327),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_328),
.A2(n_333),
.B(n_322),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_17),
.C(n_7),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_330),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_12),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_332),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_17),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_325),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_326),
.A2(n_317),
.B(n_321),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_329),
.B(n_318),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_335),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_339),
.A2(n_340),
.B(n_341),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_337),
.B(n_334),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_332),
.C(n_331),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_345),
.B(n_0),
.Y(n_346)
);


endmodule