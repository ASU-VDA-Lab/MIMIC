module fake_jpeg_28661_n_316 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_12),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_46),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_12),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_25),
.B(n_8),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_62),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_8),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_75),
.Y(n_88)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_63),
.Y(n_77)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_25),
.B(n_30),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_30),
.B(n_31),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_69),
.Y(n_96)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_40),
.Y(n_84)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_31),
.B(n_1),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g112 ( 
.A(n_72),
.B(n_73),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_18),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_34),
.B(n_21),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_34),
.B1(n_39),
.B2(n_38),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_81),
.A2(n_105),
.B1(n_106),
.B2(n_121),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_84),
.B(n_108),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_26),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_91),
.B(n_92),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_26),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_42),
.A2(n_40),
.B1(n_35),
.B2(n_38),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_93),
.A2(n_104),
.B1(n_109),
.B2(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_102),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_39),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_47),
.A2(n_40),
.B1(n_16),
.B2(n_37),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_51),
.A2(n_16),
.B1(n_37),
.B2(n_36),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_56),
.B1(n_33),
.B2(n_36),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_33),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_115),
.Y(n_146)
);

NAND2x1_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_40),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_49),
.A2(n_32),
.B1(n_21),
.B2(n_18),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_59),
.B1(n_54),
.B2(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_32),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_21),
.B1(n_18),
.B2(n_3),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_116),
.A2(n_117),
.B1(n_0),
.B2(n_9),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_61),
.A2(n_18),
.B1(n_21),
.B2(n_0),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_69),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_62),
.B(n_5),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_124),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_62),
.B(n_5),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_127),
.B(n_132),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_11),
.B1(n_10),
.B2(n_0),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_152),
.B1(n_163),
.B2(n_83),
.Y(n_168)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_0),
.B1(n_10),
.B2(n_112),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_138),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_88),
.A2(n_93),
.B(n_109),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_139),
.A2(n_149),
.B(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_96),
.B(n_90),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_142),
.B(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_77),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_99),
.Y(n_145)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_99),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_153),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_88),
.B(n_86),
.C(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_86),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_150),
.B(n_132),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_80),
.B(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_154),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_110),
.B1(n_118),
.B2(n_95),
.Y(n_152)
);

BUFx8_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_100),
.B(n_113),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_94),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_120),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_100),
.A2(n_113),
.B1(n_119),
.B2(n_79),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_164),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_123),
.A2(n_94),
.B1(n_111),
.B2(n_114),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_89),
.A2(n_111),
.B(n_114),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_128),
.Y(n_167)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_183),
.B1(n_195),
.B2(n_127),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_103),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_178),
.Y(n_201)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_103),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_135),
.B(n_147),
.Y(n_210)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_120),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_162),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_184),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_134),
.B1(n_149),
.B2(n_139),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_126),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_159),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_190),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_157),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_199),
.Y(n_209)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_151),
.B1(n_164),
.B2(n_152),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_132),
.B(n_154),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_188),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_153),
.B(n_138),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_224),
.Y(n_243)
);

NAND2x1_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_132),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_202),
.A2(n_223),
.B(n_225),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_172),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_203),
.B(n_212),
.Y(n_248)
);

OAI22x1_ASAP7_75t_SL g204 ( 
.A1(n_171),
.A2(n_130),
.B1(n_154),
.B2(n_158),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_204),
.A2(n_223),
.B1(n_202),
.B2(n_217),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_208),
.C(n_206),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_160),
.B1(n_143),
.B2(n_133),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_211),
.A2(n_217),
.B1(n_218),
.B2(n_223),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_153),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_178),
.C(n_197),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_228),
.C(n_220),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_173),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_222),
.Y(n_231)
);

OAI32xp33_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_166),
.A3(n_177),
.B1(n_167),
.B2(n_191),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_186),
.B1(n_197),
.B2(n_174),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_196),
.B1(n_175),
.B2(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_194),
.Y(n_222)
);

OR2x6_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_179),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_169),
.B(n_193),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_167),
.A2(n_181),
.B(n_191),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_169),
.B(n_170),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_219),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_170),
.C(n_182),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_187),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_198),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_234),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_223),
.B(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_236),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_198),
.B1(n_177),
.B2(n_181),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_223),
.B(n_201),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_207),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_238),
.B(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_245),
.B1(n_249),
.B2(n_225),
.Y(n_254)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_218),
.B(n_208),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_200),
.A2(n_209),
.B1(n_202),
.B2(n_211),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_221),
.C(n_214),
.Y(n_256)
);

XOR2x2_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_213),
.Y(n_252)
);

OAI322xp33_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_255),
.A3(n_249),
.B1(n_242),
.B2(n_266),
.C1(n_254),
.C2(n_264),
.Y(n_271)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_264),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_267),
.C(n_247),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_231),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_263),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_244),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_248),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_232),
.B(n_236),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_214),
.C(n_206),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_262),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_269),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_256),
.C(n_267),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_233),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_257),
.A2(n_247),
.B(n_243),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_265),
.B(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_243),
.B(n_241),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_265),
.B1(n_255),
.B2(n_230),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_284),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_252),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_283),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_277),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_233),
.C(n_237),
.Y(n_288)
);

NAND4xp25_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_289),
.C(n_269),
.D(n_274),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_SL g289 ( 
.A(n_273),
.B(n_237),
.C(n_239),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_293),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_288),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_289),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_269),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_287),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_268),
.C(n_270),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_297),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_268),
.C(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_287),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_280),
.C(n_290),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_302),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_306),
.B(n_296),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_304),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_307),
.B(n_310),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_305),
.C(n_298),
.Y(n_311)
);

AOI321xp33_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_307),
.A3(n_309),
.B1(n_292),
.B2(n_301),
.C(n_303),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_312),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_292),
.Y(n_316)
);


endmodule