module fake_jpeg_13347_n_428 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_428);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_428;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_46),
.B(n_48),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_16),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_47),
.Y(n_133)
);

BUFx12f_ASAP7_75t_SL g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_50),
.B(n_51),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

CKINVDCx9p33_ASAP7_75t_R g57 ( 
.A(n_23),
.Y(n_57)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_15),
.B(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_58),
.B(n_67),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g144 ( 
.A(n_59),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_15),
.B(n_10),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_71),
.Y(n_97)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_31),
.B(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_76),
.B(n_78),
.Y(n_142)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

BUFx16f_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_29),
.B(n_1),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_91),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_40),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_22),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_45),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_27),
.B1(n_29),
.B2(n_43),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_106),
.A2(n_121),
.B1(n_61),
.B2(n_53),
.Y(n_173)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_57),
.A2(n_29),
.B1(n_42),
.B2(n_43),
.Y(n_121)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_20),
.B1(n_34),
.B2(n_41),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_27),
.B1(n_43),
.B2(n_42),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_48),
.B(n_28),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_84),
.Y(n_152)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_52),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_91),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_140),
.B(n_37),
.Y(n_186)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g146 ( 
.A(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_146),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_46),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_153),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_148),
.A2(n_150),
.B1(n_65),
.B2(n_73),
.Y(n_196)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_106),
.A2(n_77),
.B1(n_81),
.B2(n_87),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_152),
.B(n_144),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_50),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_105),
.A2(n_56),
.B1(n_59),
.B2(n_47),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_156),
.Y(n_217)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_142),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_162),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_97),
.B(n_36),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_163),
.B(n_178),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_133),
.A2(n_59),
.B1(n_47),
.B2(n_25),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_85),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_169),
.Y(n_225)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_80),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_120),
.A2(n_35),
.B1(n_19),
.B2(n_25),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_173),
.A2(n_179),
.B1(n_103),
.B2(n_54),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_122),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_174),
.B(n_184),
.Y(n_228)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_107),
.Y(n_177)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_117),
.B(n_36),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_121),
.A2(n_41),
.B1(n_34),
.B2(n_20),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_28),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_180),
.B(n_187),
.Y(n_205)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

CKINVDCx12_ASAP7_75t_R g183 ( 
.A(n_110),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_183),
.Y(n_230)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_188),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_111),
.B(n_22),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_138),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_132),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_131),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_207),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_196),
.A2(n_116),
.B1(n_100),
.B2(n_156),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_35),
.Y(n_207)
);

NOR2x1_ASAP7_75t_R g210 ( 
.A(n_166),
.B(n_103),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

NAND2xp33_ASAP7_75t_SL g211 ( 
.A(n_169),
.B(n_166),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_211),
.B(n_175),
.C(n_165),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_224),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_154),
.B(n_169),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_95),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_159),
.B(n_144),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_218),
.B(n_223),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_220),
.A2(n_221),
.B1(n_226),
.B2(n_191),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_157),
.A2(n_93),
.B1(n_141),
.B2(n_55),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_167),
.B(n_151),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_151),
.B(n_181),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_149),
.A2(n_93),
.B1(n_60),
.B2(n_132),
.Y(n_226)
);

AND2x6_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_8),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_257),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_228),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_234),
.B(n_238),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_160),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_235),
.B(n_241),
.C(n_214),
.Y(n_284)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_228),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_171),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_240),
.B(n_243),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_176),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_184),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_244),
.A2(n_256),
.B1(n_217),
.B2(n_208),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_185),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_245),
.B(n_247),
.Y(n_288)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_95),
.B(n_177),
.C(n_92),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_246),
.A2(n_261),
.B(n_175),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_193),
.B(n_174),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_255),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_250),
.A2(n_260),
.B1(n_208),
.B2(n_217),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_204),
.B(n_99),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_251),
.B(n_253),
.Y(n_296)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_201),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_254),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_188),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_196),
.A2(n_100),
.B1(n_116),
.B2(n_182),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

AND2x6_ASAP7_75t_L g258 ( 
.A(n_195),
.B(n_7),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_264),
.Y(n_281)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_198),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_259),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_220),
.A2(n_83),
.B1(n_34),
.B2(n_41),
.Y(n_260)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_216),
.A2(n_26),
.B(n_172),
.C(n_94),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_213),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_265),
.A2(n_219),
.B(n_213),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_194),
.B1(n_197),
.B2(n_225),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_269),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_231),
.A2(n_197),
.B1(n_221),
.B2(n_226),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_271),
.A2(n_272),
.B1(n_276),
.B2(n_279),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_231),
.A2(n_211),
.B1(n_225),
.B2(n_203),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_225),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_273),
.B(n_278),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_232),
.A2(n_218),
.B(n_210),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_275),
.A2(n_258),
.B(n_259),
.Y(n_312)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_229),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_244),
.A2(n_229),
.B1(n_214),
.B2(n_198),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_239),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_284),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_285),
.B(n_265),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_254),
.Y(n_286)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_236),
.B(n_199),
.C(n_227),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_SL g301 ( 
.A(n_287),
.B(n_232),
.C(n_257),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_260),
.A2(n_227),
.B1(n_219),
.B2(n_206),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_292),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_26),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_246),
.B(n_254),
.Y(n_306)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_299),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_254),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_300),
.B(n_317),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_301),
.A2(n_306),
.B(n_275),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_271),
.A2(n_249),
.B1(n_233),
.B2(n_261),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_304),
.A2(n_322),
.B1(n_323),
.B2(n_289),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_242),
.Y(n_305)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_283),
.Y(n_307)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_307),
.Y(n_339)
);

AND2x6_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_270),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_308),
.A2(n_312),
.B(n_281),
.Y(n_324)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_252),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_319),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_296),
.B(n_237),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_314),
.Y(n_328)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_291),
.Y(n_317)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_267),
.Y(n_318)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_318),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_282),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_288),
.B(n_264),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_320),
.B(n_321),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_286),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_272),
.A2(n_256),
.B1(n_263),
.B2(n_262),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_279),
.A2(n_158),
.B1(n_145),
.B2(n_165),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_324),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_325),
.A2(n_44),
.B(n_21),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_301),
.A2(n_295),
.B(n_285),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_326),
.A2(n_330),
.B(n_345),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_311),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_341),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_312),
.A2(n_268),
.B(n_267),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_273),
.C(n_284),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_347),
.C(n_298),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_309),
.A2(n_287),
.B(n_266),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_334),
.B(n_322),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_303),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_315),
.B(n_278),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_343),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_277),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_344),
.A2(n_346),
.B1(n_310),
.B2(n_316),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_305),
.A2(n_294),
.B(n_290),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_302),
.A2(n_294),
.B1(n_290),
.B2(n_293),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_293),
.C(n_110),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_347),
.B(n_302),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_319),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_351),
.B(n_353),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_341),
.A2(n_304),
.B1(n_297),
.B2(n_303),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_352),
.B(n_361),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_297),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_354),
.A2(n_367),
.B(n_44),
.Y(n_382)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_333),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_357),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_307),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_345),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_337),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_362),
.C(n_325),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_364),
.B1(n_340),
.B2(n_339),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_318),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_338),
.C(n_326),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_328),
.A2(n_323),
.B1(n_308),
.B2(n_316),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_98),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_366),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_331),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_368),
.A2(n_382),
.B(n_21),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_363),
.A2(n_337),
.B1(n_330),
.B2(n_324),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_369),
.A2(n_350),
.B1(n_365),
.B2(n_356),
.Y(n_383)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_371),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g386 ( 
.A(n_372),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_346),
.C(n_344),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_376),
.C(n_378),
.Y(n_393)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_379),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_340),
.C(n_339),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_335),
.C(n_336),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_363),
.A2(n_335),
.B1(n_336),
.B2(n_20),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_383),
.A2(n_393),
.B1(n_389),
.B2(n_385),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_370),
.B(n_348),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_388),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_366),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_387),
.B(n_172),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_353),
.Y(n_388)
);

A2O1A1Ixp33_ASAP7_75t_L g389 ( 
.A1(n_380),
.A2(n_362),
.B(n_350),
.C(n_360),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_389),
.A2(n_392),
.B(n_113),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_127),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_381),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g394 ( 
.A(n_368),
.B(n_8),
.CI(n_45),
.CON(n_394),
.SN(n_394)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_1),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_377),
.B1(n_374),
.B2(n_380),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_395),
.A2(n_402),
.B1(n_403),
.B2(n_394),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_393),
.B(n_375),
.C(n_370),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_404),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_398),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_127),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_399),
.B(n_390),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_401),
.A2(n_388),
.B1(n_394),
.B2(n_74),
.Y(n_409)
);

BUFx12f_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_405),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_406),
.B(n_408),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_404),
.B(n_386),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_409),
.A2(n_407),
.B1(n_410),
.B2(n_398),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_94),
.C(n_84),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_410),
.B(n_412),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_404),
.A2(n_64),
.B(n_70),
.Y(n_412)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_414),
.Y(n_418)
);

A2O1A1Ixp33_ASAP7_75t_L g416 ( 
.A1(n_409),
.A2(n_397),
.B(n_400),
.C(n_3),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_416),
.B(n_411),
.Y(n_419)
);

AOI21x1_ASAP7_75t_L g422 ( 
.A1(n_419),
.A2(n_416),
.B(n_2),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_413),
.A2(n_411),
.B(n_64),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_420),
.A2(n_415),
.B(n_417),
.Y(n_421)
);

AOI322xp5_ASAP7_75t_L g423 ( 
.A1(n_421),
.A2(n_422),
.A3(n_418),
.B1(n_37),
.B2(n_3),
.C1(n_4),
.C2(n_1),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_423),
.B(n_1),
.Y(n_424)
);

AO21x1_ASAP7_75t_L g425 ( 
.A1(n_424),
.A2(n_2),
.B(n_3),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_425),
.Y(n_426)
);

AOI221xp5_ASAP7_75t_L g427 ( 
.A1(n_426),
.A2(n_63),
.B1(n_79),
.B2(n_6),
.C(n_2),
.Y(n_427)
);

OAI311xp33_ASAP7_75t_L g428 ( 
.A1(n_427),
.A2(n_2),
.A3(n_3),
.B1(n_6),
.C1(n_254),
.Y(n_428)
);


endmodule