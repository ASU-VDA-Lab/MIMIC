module fake_jpeg_27802_n_339 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_13),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_8),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_43),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_42),
.B(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_49),
.Y(n_102)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_62),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_22),
.C(n_19),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_45),
.C(n_33),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_30),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_74),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_72),
.B(n_76),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_31),
.B1(n_22),
.B2(n_19),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_95),
.B1(n_101),
.B2(n_104),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_22),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_53),
.Y(n_77)
);

NAND2x1_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_30),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_78),
.A2(n_105),
.B(n_107),
.Y(n_132)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_29),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_90),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_21),
.B(n_14),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_0),
.B(n_1),
.Y(n_112)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_99),
.Y(n_127)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_92),
.B(n_93),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_18),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_18),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_94),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_31),
.B1(n_30),
.B2(n_26),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_57),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_56),
.A2(n_31),
.B1(n_34),
.B2(n_26),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_86),
.B1(n_84),
.B2(n_79),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_48),
.A2(n_25),
.B1(n_17),
.B2(n_33),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g105 ( 
.A(n_51),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_55),
.B(n_15),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_87),
.C(n_72),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_111),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_45),
.C(n_41),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_116),
.B(n_120),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_68),
.B1(n_126),
.B2(n_82),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_73),
.B(n_15),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_25),
.B(n_32),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_33),
.C(n_32),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_131),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_33),
.C(n_32),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_80),
.B1(n_90),
.B2(n_92),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_127),
.B1(n_115),
.B2(n_131),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_106),
.Y(n_142)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_151),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_78),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_147),
.B(n_150),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_161),
.B1(n_139),
.B2(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_102),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_156),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_71),
.Y(n_153)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_83),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_122),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_1),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_111),
.CI(n_5),
.CON(n_180),
.SN(n_180)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_71),
.Y(n_158)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_109),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_127),
.B(n_102),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_165),
.Y(n_181)
);

AND2x4_ASAP7_75t_SL g163 ( 
.A(n_120),
.B(n_91),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_163),
.A2(n_166),
.B(n_167),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_116),
.B(n_103),
.Y(n_166)
);

INVx2_ASAP7_75t_R g167 ( 
.A(n_132),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_112),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_169),
.A2(n_170),
.B(n_182),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_129),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_171),
.A2(n_184),
.B1(n_188),
.B2(n_29),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_159),
.B(n_127),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_159),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_191),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_132),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_135),
.B(n_124),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_166),
.B1(n_140),
.B2(n_162),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_133),
.B1(n_121),
.B2(n_136),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_125),
.B1(n_146),
.B2(n_88),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_151),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_135),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_139),
.B(n_124),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_197),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_141),
.A2(n_121),
.B(n_136),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_150),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_202),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_194),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

CKINVDCx12_ASAP7_75t_R g204 ( 
.A(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_204),
.B(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_182),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_147),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_208),
.A2(n_213),
.B(n_181),
.Y(n_250)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_195),
.C(n_184),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_216),
.C(n_229),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_170),
.A2(n_157),
.B(n_144),
.Y(n_213)
);

NOR2x1_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_89),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_225),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_221),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_81),
.C(n_32),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_178),
.B1(n_175),
.B2(n_179),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_173),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_81),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_230),
.Y(n_254)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_227),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_169),
.A2(n_24),
.B1(n_23),
.B2(n_17),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_24),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_171),
.A2(n_24),
.B1(n_23),
.B2(n_6),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_182),
.A2(n_24),
.B1(n_23),
.B2(n_7),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_226),
.A2(n_177),
.B1(n_185),
.B2(n_192),
.Y(n_239)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_187),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_39),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_203),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_237),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_238),
.A2(n_243),
.B1(n_247),
.B2(n_206),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_239),
.A2(n_228),
.B1(n_206),
.B2(n_218),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_203),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_240),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_207),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_244),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_200),
.B1(n_180),
.B2(n_176),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_176),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_212),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_249),
.B(n_224),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_211),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_205),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_255),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_257),
.B(n_259),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_252),
.B(n_201),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_181),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_265),
.Y(n_276)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_267),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_208),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_220),
.C(n_186),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_233),
.C(n_254),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_273),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_179),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_180),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_231),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_243),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_277),
.B(n_282),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_248),
.C(n_224),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_251),
.C(n_239),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_285),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_247),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_233),
.C(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_245),
.C(n_246),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_2),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_291),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_231),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_244),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_2),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_272),
.B1(n_271),
.B2(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_270),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_300),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_293),
.A2(n_274),
.B1(n_256),
.B2(n_255),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_306),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_292),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_248),
.B1(n_261),
.B2(n_262),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_305),
.C(n_284),
.Y(n_317)
);

BUFx12_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

XOR2x1_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_291),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_309),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_276),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_313),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_277),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_283),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_283),
.B(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_316),
.A2(n_302),
.B1(n_298),
.B2(n_307),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_323),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_325),
.C(n_315),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_304),
.B(n_282),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_322),
.A2(n_324),
.B(n_314),
.Y(n_330)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_23),
.B1(n_5),
.B2(n_7),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_321),
.B(n_314),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_324),
.C(n_322),
.Y(n_328)
);

AOI322xp5_ASAP7_75t_L g332 ( 
.A1(n_328),
.A2(n_330),
.A3(n_2),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_331),
.C(n_329),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_8),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_9),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_9),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_10),
.Y(n_339)
);


endmodule