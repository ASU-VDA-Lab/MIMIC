module real_jpeg_11924_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_341, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_341;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_4),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_79),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_79),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_4),
.A2(n_67),
.B1(n_68),
.B2(n_79),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_6),
.A2(n_67),
.B1(n_68),
.B2(n_83),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_83),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_83),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_7),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_41),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_8),
.A2(n_41),
.B1(n_67),
.B2(n_68),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_41),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_8),
.A2(n_41),
.B1(n_56),
.B2(n_57),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_9),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_94),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_94),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_9),
.A2(n_56),
.B1(n_57),
.B2(n_94),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_10),
.A2(n_67),
.B1(n_68),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_10),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_176),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_176),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_176),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_12),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_66),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_66),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_12),
.A2(n_56),
.B1(n_57),
.B2(n_66),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_13),
.A2(n_67),
.B1(n_68),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_13),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_13),
.B(n_57),
.C(n_71),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_13),
.B(n_92),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_13),
.A2(n_127),
.B(n_180),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_13),
.A2(n_25),
.B(n_91),
.C(n_207),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_164),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_13),
.B(n_22),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_13),
.B(n_32),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_14),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_136),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_14),
.A2(n_67),
.B1(n_68),
.B2(n_136),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_136),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_15),
.A2(n_37),
.B1(n_56),
.B2(n_57),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_15),
.A2(n_37),
.B1(n_67),
.B2(n_68),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_149)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_42),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_29),
.B(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_22),
.A2(n_29),
.B1(n_36),
.B2(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_22),
.A2(n_29),
.B1(n_40),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_23),
.A2(n_78),
.B(n_80),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_23),
.A2(n_30),
.B1(n_78),
.B2(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_23),
.B(n_82),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_23),
.A2(n_30),
.B1(n_103),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_23),
.A2(n_80),
.B(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_23),
.A2(n_30),
.B1(n_135),
.B2(n_278),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_23)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g264 ( 
.A(n_24),
.B(n_26),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_25),
.A2(n_26),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

AOI32xp33_ASAP7_75t_L g263 ( 
.A1(n_25),
.A2(n_28),
.A3(n_33),
.B1(n_251),
.B2(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_29),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_30),
.A2(n_135),
.B(n_137),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_30),
.A2(n_33),
.B(n_164),
.C(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_38),
.B(n_339),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_39),
.B(n_336),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_335),
.B(n_337),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_323),
.B(n_334),
.Y(n_45)
);

AO21x1_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_152),
.B(n_320),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_139),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_114),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_49),
.B(n_114),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_84),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_50),
.B(n_85),
.C(n_100),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_54),
.B(n_77),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_51),
.A2(n_52),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_63),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_53),
.A2(n_54),
.B1(n_77),
.B2(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_60),
.B(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_55),
.A2(n_60),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_55),
.B(n_181),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_55),
.A2(n_60),
.B1(n_126),
.B2(n_268),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_57),
.B1(n_71),
.B2(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_56),
.B(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_60),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_60),
.B(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_62),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B1(n_74),
.B2(n_76),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_65),
.A2(n_69),
.B1(n_76),
.B2(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_68),
.B1(n_90),
.B2(n_91),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_67),
.B(n_168),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_68),
.A2(n_90),
.B(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_76),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_69),
.B(n_166),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_69),
.A2(n_76),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_69),
.A2(n_76),
.B1(n_131),
.B2(n_257),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_75),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_73),
.A2(n_175),
.B(n_177),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_73),
.B(n_164),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_73),
.A2(n_177),
.B(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_76),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_100),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_86),
.B(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_97),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_87),
.A2(n_93),
.B1(n_95),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_87),
.A2(n_95),
.B1(n_108),
.B2(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_87),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_87),
.A2(n_95),
.B1(n_227),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_87),
.A2(n_213),
.B(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_92),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_88),
.B(n_214),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_88),
.A2(n_92),
.B(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_92),
.B(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_95),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_95),
.A2(n_133),
.B(n_228),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_98),
.A2(n_163),
.B(n_165),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_98),
.A2(n_165),
.B(n_239),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_104),
.B2(n_113),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_102),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_SL g150 ( 
.A(n_102),
.B(n_105),
.C(n_110),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_102),
.B(n_143),
.C(n_150),
.Y(n_333)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_110),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_110),
.B(n_144),
.C(n_148),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.C(n_121),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_120),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_121),
.B(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_132),
.C(n_134),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_122),
.A2(n_123),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_124),
.A2(n_129),
.B1(n_130),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_124),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_127),
.A2(n_179),
.B(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_127),
.A2(n_128),
.B1(n_209),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_127),
.A2(n_128),
.B1(n_234),
.B2(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_128),
.A2(n_186),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_128),
.B(n_164),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_128),
.A2(n_194),
.B(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_132),
.B(n_134),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_138),
.B(n_249),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_139),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_151),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_140),
.B(n_151),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_145),
.Y(n_329)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_149),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_314),
.B(n_319),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_302),
.B(n_313),
.Y(n_153)
);

OAI321xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_270),
.A3(n_295),
.B1(n_300),
.B2(n_301),
.C(n_341),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_243),
.B(n_269),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_221),
.B(n_242),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_202),
.B(n_220),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_182),
.B(n_201),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_169),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_160),
.B(n_169),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_162),
.B1(n_167),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_178),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_174),
.C(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_190),
.B(n_200),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_184),
.B(n_188),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_195),
.B(n_199),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_192),
.B(n_193),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_203),
.B(n_204),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_215),
.C(n_219),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_208),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_215),
.B1(n_218),
.B2(n_219),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_222),
.B(n_223),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_235),
.B2(n_236),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_238),
.C(n_240),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_230),
.C(n_233),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_244),
.B(n_245),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_259),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_246),
.B(n_260),
.C(n_261),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_252),
.B2(n_258),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_253),
.C(n_255),
.Y(n_284)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_285),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_281),
.C(n_284),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_272),
.A2(n_273),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_279),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_279),
.C(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_277),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_281),
.B(n_284),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_283),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_294),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_289),
.C(n_294),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_293),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_292),
.C(n_293),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_312),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_312),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_307),
.C(n_308),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_333),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_333),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_332),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_328),
.B1(n_330),
.B2(n_331),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_330),
.C(n_332),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_336),
.Y(n_339)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);


endmodule