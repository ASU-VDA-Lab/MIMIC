module fake_netlist_1_57_n_20 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_20);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
OR2x2_ASAP7_75t_L g11 ( .A(n_4), .B(n_7), .Y(n_11) );
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_9), .B(n_0), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_5), .B(n_6), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_3), .B(n_10), .Y(n_15) );
OAI211xp5_ASAP7_75t_SL g16 ( .A1(n_12), .A2(n_2), .B(n_8), .C(n_13), .Y(n_16) );
INVx2_ASAP7_75t_SL g17 ( .A(n_16), .Y(n_17) );
NOR2xp33_ASAP7_75t_SL g18 ( .A(n_17), .B(n_14), .Y(n_18) );
NAND3xp33_ASAP7_75t_L g19 ( .A(n_18), .B(n_11), .C(n_15), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
endmodule