module fake_jpeg_26713_n_312 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_SL g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_36),
.Y(n_41)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_28),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_40),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_37),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_24),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_55),
.Y(n_60)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_39),
.B1(n_34),
.B2(n_17),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_67),
.B1(n_63),
.B2(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_72),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_30),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_34),
.B1(n_17),
.B2(n_32),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_68),
.B1(n_52),
.B2(n_33),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_17),
.B1(n_32),
.B2(n_40),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_17),
.B1(n_29),
.B2(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_24),
.B1(n_16),
.B2(n_20),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_70),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_71),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_49),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_42),
.B1(n_56),
.B2(n_54),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_89),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_88),
.A2(n_95),
.B(n_33),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_54),
.B1(n_42),
.B2(n_16),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_92),
.B1(n_99),
.B2(n_103),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_16),
.B1(n_22),
.B2(n_52),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_41),
.B(n_47),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_60),
.B(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_108),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_20),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_70),
.B(n_27),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_29),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_58),
.B1(n_80),
.B2(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_45),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_110),
.B(n_124),
.Y(n_150)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_106),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_82),
.C(n_73),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_121),
.C(n_115),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_15),
.B(n_26),
.C(n_25),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_19),
.B(n_15),
.Y(n_149)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_100),
.B1(n_101),
.B2(n_107),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_105),
.Y(n_139)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_30),
.B1(n_77),
.B2(n_69),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_101),
.B1(n_100),
.B2(n_86),
.Y(n_138)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_102),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_62),
.B1(n_30),
.B2(n_37),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_126),
.A2(n_87),
.B1(n_86),
.B2(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_83),
.B(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_131),
.Y(n_136)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_29),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_79),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_134),
.Y(n_174)
);

OAI22x1_ASAP7_75t_L g135 ( 
.A1(n_128),
.A2(n_93),
.B1(n_95),
.B2(n_88),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_135),
.A2(n_158),
.B(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_157),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_154),
.B1(n_147),
.B2(n_157),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_142),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_101),
.B1(n_98),
.B2(n_104),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_107),
.B1(n_28),
.B2(n_21),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_106),
.B1(n_90),
.B2(n_30),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_152),
.B1(n_119),
.B2(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_129),
.B(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_156),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_21),
.B1(n_15),
.B2(n_106),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_21),
.B1(n_37),
.B2(n_15),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_112),
.A2(n_71),
.B1(n_26),
.B2(n_19),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_25),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_123),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_57),
.B1(n_15),
.B2(n_26),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_119),
.B1(n_122),
.B2(n_118),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_187),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_164),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_117),
.B(n_116),
.C(n_131),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_188),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_172),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_117),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_113),
.B(n_114),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_133),
.C(n_151),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_176),
.B1(n_186),
.B2(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_113),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_179),
.B(n_182),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_180),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_25),
.Y(n_181)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_19),
.Y(n_182)
);

AO22x1_ASAP7_75t_SL g183 ( 
.A1(n_139),
.A2(n_57),
.B1(n_71),
.B2(n_2),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_159),
.B(n_147),
.Y(n_184)
);

NOR4xp25_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_177),
.C(n_178),
.D(n_164),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_146),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_142),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_0),
.Y(n_187)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_0),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_0),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_165),
.B(n_189),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_167),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_202),
.B1(n_161),
.B2(n_171),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_138),
.B1(n_155),
.B2(n_146),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_208),
.B1(n_176),
.B2(n_175),
.Y(n_226)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_1),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_13),
.C(n_12),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_215),
.C(n_183),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_166),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_3),
.Y(n_211)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_213),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_12),
.C(n_11),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_217),
.A2(n_201),
.B(n_214),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_197),
.B(n_186),
.CI(n_168),
.CON(n_220),
.SN(n_220)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_168),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_225),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_190),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_226),
.A2(n_235),
.B1(n_196),
.B2(n_195),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_230),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_209),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_232),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_190),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_192),
.A2(n_162),
.B1(n_174),
.B2(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_209),
.B(n_162),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_233),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_185),
.C(n_170),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_227),
.C(n_232),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_188),
.B1(n_170),
.B2(n_5),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_228),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_239),
.B1(n_208),
.B2(n_236),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_191),
.C(n_222),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_230),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_219),
.Y(n_255)
);

AOI21xp33_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_214),
.B(n_192),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_252),
.B(n_223),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_224),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_249),
.B(n_234),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_201),
.B(n_206),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_250),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_220),
.A2(n_206),
.B(n_212),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_258),
.C(n_265),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_242),
.B1(n_248),
.B2(n_226),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_254),
.B(n_255),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_245),
.B(n_220),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_256),
.A2(n_262),
.B1(n_253),
.B2(n_245),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_263),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_212),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

BUFx12_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_210),
.B1(n_191),
.B2(n_205),
.Y(n_266)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_249),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_251),
.B(n_238),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_272),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_263),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_277),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_241),
.B1(n_211),
.B2(n_204),
.Y(n_282)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_205),
.B1(n_250),
.B2(n_252),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_258),
.B1(n_260),
.B2(n_235),
.Y(n_280)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_288),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_241),
.C(n_203),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_285),
.C(n_287),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_271),
.B(n_10),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_289),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_3),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_4),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_270),
.B(n_272),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_294),
.B(n_7),
.Y(n_304)
);

AOI321xp33_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_268),
.A3(n_267),
.B1(n_276),
.B2(n_278),
.C(n_279),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_5),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_298),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_290),
.B(n_280),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_295),
.B(n_290),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_300),
.A2(n_301),
.B(n_303),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_288),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_6),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_304),
.A2(n_296),
.B(n_299),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_291),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_305),
.B(n_302),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_7),
.B1(n_8),
.B2(n_295),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_7),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_8),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_8),
.Y(n_312)
);


endmodule