module fake_jpeg_29386_n_378 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_378);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_378;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_14),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_0),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_73),
.Y(n_107)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_54),
.Y(n_89)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_56),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_59),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_32),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_65),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_76),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_34),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_27),
.Y(n_100)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_34),
.B1(n_41),
.B2(n_38),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_83),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_34),
.B1(n_38),
.B2(n_21),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_31),
.B1(n_24),
.B2(n_28),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_28),
.B1(n_31),
.B2(n_20),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_46),
.B1(n_45),
.B2(n_48),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_90),
.A2(n_103),
.B1(n_110),
.B2(n_114),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_20),
.B1(n_42),
.B2(n_39),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_100),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_34),
.B1(n_21),
.B2(n_39),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_94),
.A2(n_95),
.B1(n_118),
.B2(n_120),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_34),
.B1(n_21),
.B2(n_30),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_30),
.B1(n_42),
.B2(n_23),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_102),
.B(n_105),
.C(n_22),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_61),
.A2(n_36),
.B1(n_35),
.B2(n_43),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_51),
.A2(n_36),
.B1(n_35),
.B2(n_43),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_37),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_119),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_60),
.A2(n_37),
.B1(n_27),
.B2(n_21),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_63),
.A2(n_27),
.B1(n_21),
.B2(n_22),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_75),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_78),
.B1(n_3),
.B2(n_4),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_67),
.A2(n_27),
.B1(n_7),
.B2(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_0),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_67),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_55),
.A2(n_22),
.B1(n_9),
.B2(n_8),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_124),
.B1(n_70),
.B2(n_50),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_67),
.A2(n_9),
.B1(n_8),
.B2(n_7),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_78),
.B1(n_77),
.B2(n_71),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_126),
.A2(n_92),
.B1(n_93),
.B2(n_104),
.Y(n_176)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_128),
.B(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_59),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_131),
.B(n_145),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_109),
.Y(n_132)
);

OR2x2_ASAP7_75t_SL g133 ( 
.A(n_91),
.B(n_68),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_162),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_136),
.A2(n_143),
.B1(n_101),
.B2(n_97),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_68),
.B(n_70),
.C(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_138),
.B(n_141),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_70),
.Y(n_139)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_100),
.A3(n_90),
.B1(n_114),
.B2(n_110),
.Y(n_171)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_49),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_56),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_96),
.B(n_58),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_147),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_96),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_106),
.B(n_58),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_58),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_80),
.B(n_76),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_153),
.Y(n_180)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_80),
.B(n_22),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

BUFx4f_ASAP7_75t_SL g205 ( 
.A(n_157),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

BUFx24_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_159),
.A2(n_164),
.B1(n_97),
.B2(n_81),
.Y(n_185)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_163),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_1),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_167),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_116),
.B(n_52),
.Y(n_163)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_87),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_22),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_121),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_148),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_112),
.C(n_111),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_181),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_189),
.B1(n_136),
.B2(n_191),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_155),
.B1(n_133),
.B2(n_150),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_193),
.B1(n_202),
.B2(n_165),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_130),
.B(n_117),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_112),
.C(n_111),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_204),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_161),
.B(n_125),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_104),
.B1(n_99),
.B2(n_93),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_189),
.A2(n_135),
.B1(n_166),
.B2(n_149),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_92),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_191),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_129),
.B(n_81),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_197),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_99),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_125),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_206),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_200),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_134),
.A2(n_108),
.B1(n_3),
.B2(n_4),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_139),
.B(n_138),
.C(n_134),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_1),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_208),
.A2(n_220),
.B1(n_222),
.B2(n_225),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_209),
.A2(n_213),
.B1(n_214),
.B2(n_216),
.Y(n_270)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_215),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_204),
.A2(n_127),
.B1(n_159),
.B2(n_158),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_137),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_217),
.Y(n_242)
);

NAND2x1_ASAP7_75t_SL g219 ( 
.A(n_201),
.B(n_152),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_219),
.A2(n_192),
.B(n_205),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_169),
.A2(n_154),
.B1(n_160),
.B2(n_164),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_198),
.A2(n_108),
.B1(n_157),
.B2(n_146),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_171),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_223)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_205),
.B(n_190),
.C(n_192),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_169),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_186),
.A2(n_5),
.B1(n_172),
.B2(n_181),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_238),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_229),
.B(n_230),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_5),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_231),
.B(n_232),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_182),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_196),
.Y(n_235)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_199),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_237),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_174),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_195),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_173),
.Y(n_241)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_224),
.A2(n_172),
.B(n_197),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_245),
.A2(n_264),
.B(n_234),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_184),
.C(n_175),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_250),
.C(n_257),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_175),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_249),
.B(n_223),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_177),
.C(n_187),
.Y(n_250)
);

INVx11_ASAP7_75t_SL g253 ( 
.A(n_235),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_208),
.A2(n_176),
.B1(n_206),
.B2(n_177),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_256),
.A2(n_267),
.B1(n_214),
.B2(n_221),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_188),
.C(n_173),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_188),
.C(n_203),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_228),
.C(n_216),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_219),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_263),
.A2(n_266),
.B(n_231),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_228),
.A2(n_205),
.B(n_203),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_219),
.A2(n_207),
.B(n_190),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_239),
.A2(n_190),
.B1(n_207),
.B2(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_269),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_272),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_244),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_275),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_233),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_276),
.B(n_284),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_290),
.C(n_292),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_270),
.A2(n_223),
.B1(n_210),
.B2(n_218),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_278),
.A2(n_281),
.B1(n_287),
.B2(n_263),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_283),
.B(n_265),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_234),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_223),
.B1(n_218),
.B2(n_211),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_227),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_291),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_243),
.B(n_229),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_285),
.A2(n_246),
.B1(n_262),
.B2(n_255),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_236),
.Y(n_286)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_252),
.A2(n_245),
.B1(n_257),
.B2(n_247),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_267),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_288),
.Y(n_301)
);

NOR3xp33_ASAP7_75t_SL g289 ( 
.A(n_247),
.B(n_223),
.C(n_215),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_289),
.B(n_266),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_260),
.C(n_250),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_241),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_252),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_293),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_258),
.Y(n_294)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_296),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_298),
.A2(n_251),
.B1(n_294),
.B2(n_226),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_261),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_268),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_288),
.A3(n_278),
.B1(n_283),
.B2(n_281),
.C1(n_287),
.C2(n_282),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_292),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_285),
.B1(n_277),
.B2(n_280),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_274),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_255),
.C(n_261),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_314),
.C(n_259),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_265),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_286),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_313),
.A2(n_274),
.B(n_259),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_268),
.C(n_269),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_300),
.A2(n_272),
.B(n_279),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_315),
.B(n_320),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_306),
.Y(n_316)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_306),
.Y(n_317)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_317),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_291),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_318),
.B(n_331),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_319),
.A2(n_298),
.B1(n_303),
.B2(n_297),
.Y(n_340)
);

BUFx12_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_321),
.Y(n_341)
);

INVx13_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_273),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_326),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_327),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_313),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_330),
.C(n_305),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_258),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_342),
.C(n_344),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_340),
.B(n_343),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_310),
.C(n_314),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_312),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_334),
.A2(n_307),
.B1(n_301),
.B2(n_331),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_347),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_299),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_339),
.A2(n_323),
.B1(n_304),
.B2(n_295),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_348),
.A2(n_354),
.B(n_352),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_335),
.A2(n_301),
.B1(n_303),
.B2(n_295),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_350),
.B(n_345),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_327),
.Y(n_351)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_351),
.Y(n_363)
);

AO21x1_ASAP7_75t_L g352 ( 
.A1(n_343),
.A2(n_315),
.B(n_328),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_352),
.B(n_319),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_321),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_353),
.A2(n_332),
.B1(n_316),
.B2(n_317),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_332),
.A2(n_321),
.B(n_322),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_347),
.B(n_336),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_355),
.A2(n_354),
.B(n_344),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_357),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_360),
.C(n_349),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_349),
.B(n_318),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_361),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_346),
.A2(n_342),
.B(n_338),
.Y(n_362)
);

MAJx2_ASAP7_75t_L g365 ( 
.A(n_362),
.B(n_346),
.C(n_351),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_365),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_353),
.C(n_338),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_366),
.B(n_369),
.Y(n_373)
);

AO21x1_ASAP7_75t_L g372 ( 
.A1(n_367),
.A2(n_363),
.B(n_358),
.Y(n_372)
);

BUFx24_ASAP7_75t_SL g371 ( 
.A(n_368),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_371),
.A2(n_372),
.B(n_370),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_373),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_374),
.A2(n_350),
.B(n_325),
.Y(n_376)
);

O2A1O1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_376),
.A2(n_363),
.B(n_375),
.C(n_360),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_377),
.A2(n_251),
.B(n_311),
.Y(n_378)
);


endmodule