module real_aes_2813_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_836, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_837, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_836;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_837;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_335;
wire n_177;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g179 ( .A(n_0), .B(n_153), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_1), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_2), .B(n_114), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_3), .Y(n_832) );
INVx1_ASAP7_75t_L g144 ( .A(n_4), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_5), .B(n_137), .Y(n_206) );
NAND2xp33_ASAP7_75t_SL g249 ( .A(n_6), .B(n_143), .Y(n_249) );
INVx1_ASAP7_75t_L g241 ( .A(n_7), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_8), .B(n_211), .Y(n_499) );
INVx1_ASAP7_75t_L g480 ( .A(n_9), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_10), .Y(n_114) );
AND2x2_ASAP7_75t_L g204 ( .A(n_11), .B(n_161), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_12), .Y(n_563) );
INVx2_ASAP7_75t_L g159 ( .A(n_13), .Y(n_159) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_14), .Y(n_115) );
INVx1_ASAP7_75t_L g507 ( .A(n_15), .Y(n_507) );
AOI221x1_ASAP7_75t_L g244 ( .A1(n_16), .A2(n_146), .B1(n_245), .B2(n_247), .C(n_248), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_17), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g111 ( .A(n_18), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_19), .Y(n_799) );
INVx1_ASAP7_75t_L g505 ( .A(n_20), .Y(n_505) );
INVx1_ASAP7_75t_SL g517 ( .A(n_21), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_22), .B(n_138), .Y(n_495) );
AOI221xp5_ASAP7_75t_SL g168 ( .A1(n_23), .A2(n_44), .B1(n_137), .B2(n_146), .C(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_24), .A2(n_146), .B(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_25), .B(n_153), .Y(n_209) );
AOI33xp33_ASAP7_75t_L g472 ( .A1(n_26), .A2(n_56), .A3(n_192), .B1(n_199), .B2(n_473), .B3(n_474), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_27), .A2(n_42), .B1(n_824), .B2(n_825), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_27), .Y(n_825) );
INVx1_ASAP7_75t_L g557 ( .A(n_28), .Y(n_557) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_29), .A2(n_119), .B1(n_120), .B2(n_126), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_29), .Y(n_126) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_30), .A2(n_93), .B(n_159), .Y(n_158) );
OR2x2_ASAP7_75t_L g162 ( .A(n_30), .B(n_93), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_31), .B(n_155), .Y(n_154) );
INVxp67_ASAP7_75t_L g243 ( .A(n_32), .Y(n_243) );
AND2x2_ASAP7_75t_L g230 ( .A(n_33), .B(n_167), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_34), .B(n_190), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_35), .A2(n_146), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_36), .B(n_660), .Y(n_659) );
CKINVDCx16_ASAP7_75t_R g783 ( .A(n_36), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_37), .B(n_155), .Y(n_170) );
AND2x2_ASAP7_75t_L g143 ( .A(n_38), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g147 ( .A(n_38), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g198 ( .A(n_38), .Y(n_198) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_39), .B(n_113), .C(n_115), .Y(n_112) );
OR2x6_ASAP7_75t_L g787 ( .A(n_39), .B(n_788), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_40), .A2(n_73), .B1(n_820), .B2(n_821), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_40), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_41), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_42), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_43), .B(n_190), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_45), .A2(n_121), .B1(n_122), .B2(n_123), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_45), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_46), .A2(n_175), .B1(n_211), .B2(n_489), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_47), .A2(n_85), .B1(n_146), .B2(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_48), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_49), .B(n_138), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_50), .B(n_153), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_51), .B(n_157), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_52), .B(n_138), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_53), .Y(n_492) );
AND2x2_ASAP7_75t_L g182 ( .A(n_54), .B(n_167), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_55), .B(n_167), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_57), .B(n_138), .Y(n_463) );
INVx1_ASAP7_75t_L g140 ( .A(n_58), .Y(n_140) );
INVx1_ASAP7_75t_L g150 ( .A(n_58), .Y(n_150) );
AND2x2_ASAP7_75t_L g464 ( .A(n_59), .B(n_167), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_60), .A2(n_78), .B1(n_190), .B2(n_196), .C(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_61), .B(n_190), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_62), .B(n_137), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_63), .B(n_175), .Y(n_565) );
AOI21xp5_ASAP7_75t_SL g525 ( .A1(n_64), .A2(n_196), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g221 ( .A(n_65), .B(n_167), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_66), .B(n_155), .Y(n_180) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_67), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_68), .B(n_153), .Y(n_218) );
INVx1_ASAP7_75t_L g502 ( .A(n_69), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_70), .A2(n_146), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g461 ( .A(n_71), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_72), .B(n_155), .Y(n_210) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_73), .B(n_157), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_73), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_74), .A2(n_196), .B(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_75), .A2(n_97), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_75), .Y(n_124) );
INVx1_ASAP7_75t_L g142 ( .A(n_76), .Y(n_142) );
INVx1_ASAP7_75t_L g148 ( .A(n_76), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_77), .B(n_190), .Y(n_475) );
AND2x2_ASAP7_75t_L g519 ( .A(n_79), .B(n_247), .Y(n_519) );
INVx1_ASAP7_75t_L g503 ( .A(n_80), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_81), .A2(n_196), .B(n_516), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_82), .A2(n_187), .B(n_196), .C(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_83), .A2(n_88), .B1(n_137), .B2(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_84), .B(n_137), .Y(n_219) );
INVx1_ASAP7_75t_L g110 ( .A(n_86), .Y(n_110) );
AND2x2_ASAP7_75t_SL g523 ( .A(n_87), .B(n_247), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_89), .A2(n_196), .B1(n_470), .B2(n_471), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_90), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_91), .B(n_153), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_92), .A2(n_146), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g527 ( .A(n_94), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_95), .B(n_155), .Y(n_217) );
AND2x2_ASAP7_75t_L g476 ( .A(n_96), .B(n_247), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_97), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_98), .A2(n_555), .B(n_556), .C(n_558), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_99), .B(n_137), .Y(n_181) );
INVxp67_ASAP7_75t_L g246 ( .A(n_100), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_101), .B(n_155), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_102), .A2(n_146), .B(n_151), .Y(n_145) );
BUFx2_ASAP7_75t_L g810 ( .A(n_103), .Y(n_810) );
BUFx2_ASAP7_75t_SL g830 ( .A(n_103), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_104), .B(n_138), .Y(n_528) );
AOI21xp33_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_116), .B(n_831), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_107), .Y(n_834) );
INVx3_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_112), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_110), .B(n_111), .Y(n_788) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_115), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_115), .B(n_446), .Y(n_445) );
OR2x6_ASAP7_75t_SL g793 ( .A(n_115), .B(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_115), .B(n_794), .Y(n_804) );
OR2x2_ASAP7_75t_L g808 ( .A(n_115), .B(n_787), .Y(n_808) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_811), .Y(n_116) );
A2O1A1Ixp33_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_127), .B(n_785), .C(n_789), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g785 ( .A1(n_118), .A2(n_786), .B(n_787), .Y(n_785) );
INVxp67_ASAP7_75t_SL g796 ( .A(n_118), .Y(n_796) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_443), .B(n_445), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx3_ASAP7_75t_SL g795 ( .A(n_129), .Y(n_795) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_335), .Y(n_129) );
NOR3xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_263), .C(n_313), .Y(n_130) );
OAI211xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_183), .B(n_231), .C(n_252), .Y(n_131) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_163), .Y(n_132) );
AND2x2_ASAP7_75t_L g262 ( .A(n_133), .B(n_164), .Y(n_262) );
INVx1_ASAP7_75t_L g393 ( .A(n_133), .Y(n_393) );
NOR2x1p5_ASAP7_75t_L g425 ( .A(n_133), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g236 ( .A(n_134), .B(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g284 ( .A(n_134), .Y(n_284) );
OR2x2_ASAP7_75t_L g288 ( .A(n_134), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_134), .B(n_166), .Y(n_300) );
OR2x2_ASAP7_75t_L g322 ( .A(n_134), .B(n_166), .Y(n_322) );
AND2x4_ASAP7_75t_L g328 ( .A(n_134), .B(n_292), .Y(n_328) );
OR2x2_ASAP7_75t_L g345 ( .A(n_134), .B(n_238), .Y(n_345) );
INVx1_ASAP7_75t_L g380 ( .A(n_134), .Y(n_380) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_134), .Y(n_402) );
OR2x2_ASAP7_75t_L g416 ( .A(n_134), .B(n_349), .Y(n_416) );
AND2x4_ASAP7_75t_SL g420 ( .A(n_134), .B(n_238), .Y(n_420) );
OR2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_160), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_145), .B(n_157), .Y(n_135) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_143), .Y(n_137) );
INVx1_ASAP7_75t_L g250 ( .A(n_138), .Y(n_250) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
AND2x6_ASAP7_75t_L g153 ( .A(n_139), .B(n_148), .Y(n_153) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g155 ( .A(n_141), .B(n_150), .Y(n_155) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx5_ASAP7_75t_L g156 ( .A(n_143), .Y(n_156) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_143), .Y(n_558) );
AND2x2_ASAP7_75t_L g149 ( .A(n_144), .B(n_150), .Y(n_149) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_144), .Y(n_193) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
BUFx3_ASAP7_75t_L g194 ( .A(n_147), .Y(n_194) );
INVx2_ASAP7_75t_L g200 ( .A(n_148), .Y(n_200) );
AND2x4_ASAP7_75t_L g196 ( .A(n_149), .B(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g192 ( .A(n_150), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_154), .B(n_156), .Y(n_151) );
INVxp67_ASAP7_75t_L g506 ( .A(n_153), .Y(n_506) );
INVxp67_ASAP7_75t_L g508 ( .A(n_155), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_156), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_156), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_156), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_156), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_156), .A2(n_227), .B(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_156), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
INVx1_ASAP7_75t_L g470 ( .A(n_156), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_156), .A2(n_462), .B(n_480), .C(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_156), .A2(n_495), .B(n_496), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_156), .B(n_211), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_156), .A2(n_462), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_156), .A2(n_462), .B(n_527), .C(n_528), .Y(n_526) );
INVx2_ASAP7_75t_SL g187 ( .A(n_157), .Y(n_187) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_157), .A2(n_478), .B(n_482), .Y(n_477) );
BUFx4f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx3_ASAP7_75t_L g175 ( .A(n_158), .Y(n_175) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_159), .B(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g211 ( .A(n_159), .B(n_162), .Y(n_211) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_161), .Y(n_167) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g372 ( .A(n_164), .B(n_328), .Y(n_372) );
AND2x2_ASAP7_75t_L g419 ( .A(n_164), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_173), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g235 ( .A(n_166), .Y(n_235) );
AND2x2_ASAP7_75t_L g282 ( .A(n_166), .B(n_173), .Y(n_282) );
INVx2_ASAP7_75t_L g289 ( .A(n_166), .Y(n_289) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_166), .Y(n_410) );
BUFx3_ASAP7_75t_L g426 ( .A(n_166), .Y(n_426) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_172), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_167), .Y(n_220) );
INVx2_ASAP7_75t_L g251 ( .A(n_173), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_173), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g349 ( .A(n_173), .B(n_289), .Y(n_349) );
INVx1_ASAP7_75t_L g367 ( .A(n_173), .Y(n_367) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_173), .Y(n_383) );
INVx1_ASAP7_75t_L g405 ( .A(n_173), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_173), .B(n_284), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_173), .B(n_238), .Y(n_442) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AOI21x1_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_182), .Y(n_174) );
INVx4_ASAP7_75t_L g247 ( .A(n_175), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_175), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_181), .Y(n_176) );
INVx1_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_202), .Y(n_184) );
AND2x4_ASAP7_75t_L g256 ( .A(n_185), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g267 ( .A(n_185), .Y(n_267) );
AND2x2_ASAP7_75t_L g272 ( .A(n_185), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g307 ( .A(n_185), .B(n_212), .Y(n_307) );
AND2x2_ASAP7_75t_L g317 ( .A(n_185), .B(n_213), .Y(n_317) );
OR2x2_ASAP7_75t_L g397 ( .A(n_185), .B(n_312), .Y(n_397) );
OAI322xp33_ASAP7_75t_L g427 ( .A1(n_185), .A2(n_340), .A3(n_379), .B1(n_412), .B2(n_428), .C1(n_429), .C2(n_430), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_185), .B(n_410), .Y(n_428) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g261 ( .A(n_186), .Y(n_261) );
AOI21x1_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_201), .Y(n_186) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_187), .A2(n_468), .B(n_476), .Y(n_467) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_187), .A2(n_468), .B(n_476), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_195), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_190), .A2(n_196), .B1(n_240), .B2(n_242), .Y(n_239) );
INVx1_ASAP7_75t_L g566 ( .A(n_190), .Y(n_566) );
AND2x4_ASAP7_75t_L g190 ( .A(n_191), .B(n_194), .Y(n_190) );
INVx1_ASAP7_75t_L g490 ( .A(n_191), .Y(n_490) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
OR2x6_ASAP7_75t_L g462 ( .A(n_192), .B(n_200), .Y(n_462) );
INVxp33_ASAP7_75t_L g473 ( .A(n_192), .Y(n_473) );
INVx1_ASAP7_75t_L g491 ( .A(n_194), .Y(n_491) );
INVxp67_ASAP7_75t_L g564 ( .A(n_196), .Y(n_564) );
NOR2x1p5_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVx1_ASAP7_75t_L g474 ( .A(n_199), .Y(n_474) );
INVx3_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_202), .A2(n_374), .B1(n_378), .B2(n_381), .Y(n_373) );
AOI211xp5_ASAP7_75t_L g433 ( .A1(n_202), .A2(n_434), .B(n_435), .C(n_438), .Y(n_433) );
AND2x4_ASAP7_75t_SL g202 ( .A(n_203), .B(n_212), .Y(n_202) );
AND2x4_ASAP7_75t_L g255 ( .A(n_203), .B(n_223), .Y(n_255) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_203), .Y(n_259) );
INVx5_ASAP7_75t_L g271 ( .A(n_203), .Y(n_271) );
INVx2_ASAP7_75t_L g280 ( .A(n_203), .Y(n_280) );
AND2x2_ASAP7_75t_L g303 ( .A(n_203), .B(n_213), .Y(n_303) );
AND2x2_ASAP7_75t_L g332 ( .A(n_203), .B(n_222), .Y(n_332) );
OR2x2_ASAP7_75t_L g341 ( .A(n_203), .B(n_261), .Y(n_341) );
OR2x2_ASAP7_75t_L g356 ( .A(n_203), .B(n_270), .Y(n_356) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_211), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_211), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_211), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_211), .B(n_246), .Y(n_245) );
NOR3xp33_ASAP7_75t_L g248 ( .A(n_211), .B(n_249), .C(n_250), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_211), .A2(n_525), .B(n_529), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_212), .B(n_232), .Y(n_231) );
INVx3_ASAP7_75t_SL g340 ( .A(n_212), .Y(n_340) );
AND2x2_ASAP7_75t_L g363 ( .A(n_212), .B(n_271), .Y(n_363) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_222), .Y(n_212) );
INVx2_ASAP7_75t_L g257 ( .A(n_213), .Y(n_257) );
AND2x2_ASAP7_75t_L g260 ( .A(n_213), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g274 ( .A(n_213), .B(n_223), .Y(n_274) );
INVx1_ASAP7_75t_L g278 ( .A(n_213), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_213), .B(n_223), .Y(n_312) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_213), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_213), .B(n_271), .Y(n_387) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_220), .B(n_221), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_219), .Y(n_214) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_220), .A2(n_224), .B(n_230), .Y(n_223) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_220), .A2(n_224), .B(n_230), .Y(n_270) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_220), .A2(n_513), .B(n_519), .Y(n_512) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_223), .Y(n_293) );
AND2x2_ASAP7_75t_L g377 ( .A(n_223), .B(n_261), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_229), .Y(n_224) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_236), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_233), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OR2x6_ASAP7_75t_SL g441 ( .A(n_234), .B(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_235), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_235), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g389 ( .A(n_235), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_236), .A2(n_298), .B1(n_301), .B2(n_308), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_237), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g333 ( .A(n_237), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_237), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_SL g388 ( .A(n_237), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_251), .Y(n_237) );
AND2x2_ASAP7_75t_L g283 ( .A(n_238), .B(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g292 ( .A(n_238), .Y(n_292) );
OAI22xp33_ASAP7_75t_L g350 ( .A1(n_238), .A2(n_299), .B1(n_351), .B2(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g358 ( .A(n_238), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_238), .B(n_352), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_238), .B(n_282), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_238), .B(n_289), .Y(n_431) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_244), .Y(n_238) );
INVx3_ASAP7_75t_L g456 ( .A(n_247), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_247), .A2(n_456), .B1(n_554), .B2(n_559), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_250), .A2(n_462), .B1(n_502), .B2(n_503), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_250), .B(n_557), .Y(n_556) );
OAI21xp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_258), .B(n_262), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
NAND4xp25_ASAP7_75t_SL g301 ( .A(n_254), .B(n_302), .C(n_304), .D(n_306), .Y(n_301) );
INVx2_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_255), .B(n_362), .Y(n_391) );
AND2x2_ASAP7_75t_L g418 ( .A(n_255), .B(n_256), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_255), .B(n_278), .Y(n_429) );
INVx1_ASAP7_75t_L g294 ( .A(n_256), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_256), .A2(n_319), .B1(n_330), .B2(n_333), .Y(n_329) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_256), .B(n_269), .C(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_256), .B(n_271), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_256), .B(n_279), .Y(n_422) );
AND2x2_ASAP7_75t_L g354 ( .A(n_257), .B(n_261), .Y(n_354) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_257), .Y(n_415) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g310 ( .A(n_259), .Y(n_310) );
INVx1_ASAP7_75t_L g400 ( .A(n_260), .Y(n_400) );
AND2x2_ASAP7_75t_L g407 ( .A(n_260), .B(n_271), .Y(n_407) );
BUFx2_ASAP7_75t_L g362 ( .A(n_261), .Y(n_362) );
NAND3xp33_ASAP7_75t_SL g263 ( .A(n_264), .B(n_285), .C(n_297), .Y(n_263) );
OAI31xp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_272), .A3(n_275), .B(n_281), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_265), .A2(n_319), .B1(n_323), .B2(n_324), .Y(n_318) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
OR2x2_ASAP7_75t_L g304 ( .A(n_267), .B(n_305), .Y(n_304) );
NOR2x1_ASAP7_75t_L g330 ( .A(n_267), .B(n_331), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_268), .A2(n_370), .B(n_400), .C(n_401), .Y(n_399) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_269), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_270), .B(n_278), .Y(n_305) );
AND2x2_ASAP7_75t_L g323 ( .A(n_270), .B(n_303), .Y(n_323) );
AND2x2_ASAP7_75t_L g440 ( .A(n_273), .B(n_362), .Y(n_440) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g296 ( .A(n_274), .B(n_280), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_279), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_279), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g371 ( .A(n_279), .B(n_354), .Y(n_371) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_280), .B(n_354), .Y(n_360) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g352 ( .A(n_282), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_283), .B(n_383), .Y(n_382) );
AOI32xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_293), .A3(n_294), .B1(n_295), .B2(n_836), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_286), .A2(n_371), .B1(n_407), .B2(n_408), .C(n_411), .Y(n_406) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_289), .Y(n_334) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g299 ( .A(n_291), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g404 ( .A(n_292), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_293), .B(n_315), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_295), .A2(n_338), .B1(n_342), .B2(n_346), .C(n_350), .Y(n_337) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI211xp5_ASAP7_75t_L g313 ( .A1(n_300), .A2(n_314), .B(n_318), .C(n_329), .Y(n_313) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI322xp33_ASAP7_75t_L g411 ( .A1(n_306), .A2(n_316), .A3(n_365), .B1(n_412), .B2(n_413), .C1(n_414), .C2(n_416), .Y(n_411) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AOI21xp33_ASAP7_75t_L g438 ( .A1(n_309), .A2(n_439), .B(n_441), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g395 ( .A1(n_315), .A2(n_396), .B(n_398), .C(n_399), .Y(n_395) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g437 ( .A(n_322), .B(n_403), .Y(n_437) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVxp67_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_328), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g412 ( .A(n_328), .Y(n_412) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI31xp33_ASAP7_75t_L g368 ( .A1(n_332), .A2(n_369), .A3(n_371), .B(n_372), .Y(n_368) );
NOR2x1_ASAP7_75t_L g335 ( .A(n_336), .B(n_394), .Y(n_335) );
NAND5xp2_ASAP7_75t_L g336 ( .A(n_337), .B(n_357), .C(n_368), .D(n_373), .E(n_384), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AOI21xp33_ASAP7_75t_L g435 ( .A1(n_340), .A2(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g408 ( .A(n_344), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B(n_361), .C(n_364), .Y(n_357) );
INVxp33_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
OR2x2_ASAP7_75t_L g386 ( .A(n_362), .B(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_365), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g436 ( .A(n_377), .Y(n_436) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .B(n_390), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI21xp33_ASAP7_75t_L g390 ( .A1(n_386), .A2(n_391), .B(n_392), .Y(n_390) );
NAND4xp25_ASAP7_75t_L g394 ( .A(n_395), .B(n_406), .C(n_417), .D(n_433), .Y(n_394) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_404), .B(n_425), .Y(n_424) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g434 ( .A(n_416), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_421), .B2(n_423), .C(n_427), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g786 ( .A(n_445), .Y(n_786) );
INVx2_ASAP7_75t_L g817 ( .A(n_446), .Y(n_817) );
OR2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_780), .Y(n_446) );
NOR4xp25_ASAP7_75t_L g447 ( .A(n_448), .B(n_659), .C(n_683), .D(n_749), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_448), .A2(n_683), .B1(n_783), .B2(n_837), .Y(n_784) );
NAND3x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_611), .C(n_645), .Y(n_448) );
NOR3x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_570), .C(n_590), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_545), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_483), .B1(n_534), .B2(n_542), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_465), .Y(n_452) );
AND2x2_ASAP7_75t_L g709 ( .A(n_453), .B(n_639), .Y(n_709) );
INVx1_ASAP7_75t_L g716 ( .A(n_453), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_453), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_453), .B(n_579), .Y(n_768) );
OR2x2_ASAP7_75t_L g778 ( .A(n_453), .B(n_779), .Y(n_778) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2x1p5_ASAP7_75t_L g599 ( .A(n_454), .B(n_536), .Y(n_599) );
AND2x4_ASAP7_75t_L g627 ( .A(n_454), .B(n_541), .Y(n_627) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g575 ( .A(n_455), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_455), .B(n_467), .Y(n_665) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_455), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_455), .B(n_552), .Y(n_702) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B(n_464), .Y(n_455) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_456), .A2(n_457), .B(n_464), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx2_ASAP7_75t_L g497 ( .A(n_462), .Y(n_497) );
INVxp67_ASAP7_75t_L g555 ( .A(n_462), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_465), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g773 ( .A(n_465), .B(n_610), .Y(n_773) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g763 ( .A(n_466), .B(n_702), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_477), .Y(n_466) );
INVx2_ASAP7_75t_L g541 ( .A(n_467), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_469), .B(n_475), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g537 ( .A(n_477), .Y(n_537) );
INVx2_ASAP7_75t_L g551 ( .A(n_477), .Y(n_551) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_477), .Y(n_576) );
INVx1_ASAP7_75t_L g589 ( .A(n_477), .Y(n_589) );
INVxp67_ASAP7_75t_L g608 ( .A(n_477), .Y(n_608) );
AND2x4_ASAP7_75t_L g639 ( .A(n_477), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_520), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_510), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g681 ( .A(n_486), .B(n_668), .Y(n_681) );
AND2x2_ASAP7_75t_L g705 ( .A(n_486), .B(n_521), .Y(n_705) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_498), .Y(n_486) );
INVx2_ASAP7_75t_L g533 ( .A(n_487), .Y(n_533) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_487), .Y(n_548) );
INVx1_ASAP7_75t_L g605 ( .A(n_487), .Y(n_605) );
AND2x4_ASAP7_75t_L g614 ( .A(n_487), .B(n_532), .Y(n_614) );
AND2x2_ASAP7_75t_L g670 ( .A(n_487), .B(n_522), .Y(n_670) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_493), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .C(n_492), .Y(n_489) );
INVx3_ASAP7_75t_L g532 ( .A(n_498), .Y(n_532) );
AND2x2_ASAP7_75t_L g544 ( .A(n_498), .B(n_512), .Y(n_544) );
INVx2_ASAP7_75t_L g583 ( .A(n_498), .Y(n_583) );
NOR2x1_ASAP7_75t_SL g596 ( .A(n_498), .B(n_522), .Y(n_596) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_504), .B(n_509), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B1(n_507), .B2(n_508), .Y(n_504) );
INVx1_ASAP7_75t_L g698 ( .A(n_510), .Y(n_698) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g621 ( .A(n_511), .Y(n_621) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_512), .Y(n_579) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_512), .Y(n_595) );
AND2x2_ASAP7_75t_L g603 ( .A(n_512), .B(n_532), .Y(n_603) );
INVx1_ASAP7_75t_L g643 ( .A(n_512), .Y(n_643) );
INVx1_ASAP7_75t_L g668 ( .A(n_512), .Y(n_668) );
OR2x2_ASAP7_75t_L g729 ( .A(n_512), .B(n_522), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
OA211x2_ASAP7_75t_L g750 ( .A1(n_520), .A2(n_751), .B(n_753), .C(n_760), .Y(n_750) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
AND2x2_ASAP7_75t_L g671 ( .A(n_521), .B(n_544), .Y(n_671) );
AND2x2_ASAP7_75t_SL g689 ( .A(n_521), .B(n_531), .Y(n_689) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g543 ( .A(n_522), .Y(n_543) );
INVx2_ASAP7_75t_L g585 ( .A(n_522), .Y(n_585) );
AND2x4_ASAP7_75t_L g648 ( .A(n_522), .B(n_605), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_522), .B(n_644), .Y(n_699) );
AND2x2_ASAP7_75t_L g742 ( .A(n_522), .B(n_583), .Y(n_742) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_531), .B(n_643), .Y(n_736) );
AND2x2_ASAP7_75t_L g756 ( .A(n_531), .B(n_579), .Y(n_756) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g644 ( .A(n_532), .Y(n_644) );
INVx1_ASAP7_75t_L g618 ( .A(n_533), .Y(n_618) );
NOR2xp67_ASAP7_75t_SL g534 ( .A(n_535), .B(n_538), .Y(n_534) );
INVx1_ASAP7_75t_L g712 ( .A(n_535), .Y(n_712) );
NOR2xp67_ASAP7_75t_L g759 ( .A(n_535), .B(n_713), .Y(n_759) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g732 ( .A(n_537), .B(n_574), .Y(n_732) );
OAI211xp5_ASAP7_75t_L g720 ( .A1(n_538), .A2(n_721), .B(n_724), .C(n_733), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g764 ( .A1(n_538), .A2(n_758), .B(n_765), .C(n_769), .Y(n_764) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g649 ( .A(n_539), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g568 ( .A(n_540), .Y(n_568) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_540), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g624 ( .A(n_540), .B(n_574), .Y(n_624) );
NOR2xp67_ASAP7_75t_L g734 ( .A(n_540), .B(n_574), .Y(n_734) );
AND2x2_ASAP7_75t_L g607 ( .A(n_541), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g658 ( .A(n_541), .Y(n_658) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
AND2x4_ASAP7_75t_SL g547 ( .A(n_543), .B(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g604 ( .A(n_543), .B(n_605), .Y(n_604) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_543), .B(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g652 ( .A(n_543), .B(n_653), .Y(n_652) );
NOR2xp67_ASAP7_75t_SL g735 ( .A(n_543), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_SL g546 ( .A(n_544), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_SL g775 ( .A(n_544), .B(n_617), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_549), .Y(n_545) );
INVx2_ASAP7_75t_SL g743 ( .A(n_549), .Y(n_743) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_567), .Y(n_549) );
INVx3_ASAP7_75t_L g666 ( .A(n_550), .Y(n_666) );
AND2x2_ASAP7_75t_L g687 ( .A(n_550), .B(n_678), .Y(n_687) );
AND2x2_ASAP7_75t_L g745 ( .A(n_550), .B(n_627), .Y(n_745) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx2_ASAP7_75t_L g574 ( .A(n_552), .Y(n_574) );
INVx1_ASAP7_75t_L g610 ( .A(n_552), .Y(n_610) );
INVx1_ASAP7_75t_L g630 ( .A(n_552), .Y(n_630) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_560), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .B1(n_565), .B2(n_566), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVxp67_ASAP7_75t_L g713 ( .A(n_567), .Y(n_713) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g573 ( .A(n_569), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g640 ( .A(n_569), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_577), .B1(n_580), .B2(n_586), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
AND2x2_ASAP7_75t_L g587 ( .A(n_573), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g598 ( .A(n_573), .Y(n_598) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g647 ( .A(n_578), .B(n_648), .Y(n_647) );
BUFx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVxp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g667 ( .A(n_582), .B(n_668), .Y(n_667) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g675 ( .A(n_583), .Y(n_675) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g723 ( .A(n_585), .B(n_614), .Y(n_723) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_587), .A2(n_681), .B(n_682), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_597), .B(n_600), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g646 ( .A(n_596), .B(n_620), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_597), .A2(n_704), .B1(n_706), .B2(n_708), .Y(n_703) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_606), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_SL g653 ( .A(n_603), .Y(n_653) );
AND2x2_ASAP7_75t_L g682 ( .A(n_604), .B(n_620), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_604), .B(n_642), .Y(n_714) );
AND2x2_ASAP7_75t_L g718 ( .A(n_604), .B(n_675), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g662 ( .A1(n_606), .A2(n_663), .B(n_667), .Y(n_662) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
AND2x2_ASAP7_75t_L g623 ( .A(n_607), .B(n_624), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g700 ( .A(n_607), .B(n_701), .Y(n_700) );
BUFx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g692 ( .A(n_610), .Y(n_692) );
NOR2x1_ASAP7_75t_L g611 ( .A(n_612), .B(n_635), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_622), .B1(n_625), .B2(n_631), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx4_ASAP7_75t_L g634 ( .A(n_614), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_614), .B(n_620), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_614), .B(n_767), .Y(n_766) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_617), .A2(n_641), .B(n_705), .Y(n_704) );
AND2x4_ASAP7_75t_L g740 ( .A(n_617), .B(n_642), .Y(n_740) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g722 ( .A(n_619), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g758 ( .A(n_620), .B(n_742), .Y(n_758) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g638 ( .A(n_624), .B(n_639), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g657 ( .A(n_624), .B(n_658), .Y(n_657) );
OAI22xp5_ASAP7_75t_SL g635 ( .A1(n_625), .A2(n_636), .B1(n_637), .B2(n_641), .Y(n_635) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g752 ( .A(n_629), .B(n_639), .Y(n_752) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g650 ( .A(n_630), .Y(n_650) );
AND2x2_ASAP7_75t_L g676 ( .A(n_630), .B(n_639), .Y(n_676) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_632), .B(n_773), .Y(n_772) );
BUFx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_633), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g727 ( .A(n_634), .Y(n_727) );
INVx1_ASAP7_75t_L g739 ( .A(n_636), .Y(n_739) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_638), .A2(n_682), .B1(n_761), .B2(n_762), .Y(n_760) );
AND2x2_ASAP7_75t_L g677 ( .A(n_639), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g748 ( .A(n_639), .B(n_701), .Y(n_748) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI211xp5_ASAP7_75t_SL g651 ( .A1(n_642), .A2(n_652), .B(n_654), .C(n_655), .Y(n_651) );
AND2x2_ASAP7_75t_SL g761 ( .A(n_642), .B(n_648), .Y(n_761) );
AND2x4_ASAP7_75t_SL g642 ( .A(n_643), .B(n_644), .Y(n_642) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_643), .Y(n_695) );
O2A1O1Ixp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B(n_649), .C(n_651), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_646), .A2(n_674), .B1(n_676), .B2(n_677), .Y(n_673) );
INVx2_ASAP7_75t_L g654 ( .A(n_648), .Y(n_654) );
AND2x2_ASAP7_75t_L g674 ( .A(n_648), .B(n_675), .Y(n_674) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_648), .Y(n_741) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVxp67_ASAP7_75t_L g782 ( .A(n_660), .Y(n_782) );
NOR2x1_ASAP7_75t_SL g660 ( .A(n_661), .B(n_672), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_669), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_663), .A2(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g693 ( .A(n_665), .Y(n_693) );
INVx1_ASAP7_75t_L g769 ( .A(n_666), .Y(n_769) );
AND2x2_ASAP7_75t_L g707 ( .A(n_670), .B(n_695), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_671), .B(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_673), .B(n_680), .Y(n_672) );
AND2x2_ASAP7_75t_L g774 ( .A(n_676), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2x1_ASAP7_75t_L g683 ( .A(n_684), .B(n_719), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_703), .C(n_710), .Y(n_684) );
OAI222xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B1(n_690), .B2(n_694), .C1(n_696), .C2(n_700), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2x1_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx2_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g746 ( .A(n_705), .Y(n_746) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_714), .B1(n_715), .B2(n_717), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NOR2xp67_ASAP7_75t_SL g719 ( .A(n_720), .B(n_737), .Y(n_719) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_730), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_727), .B(n_748), .Y(n_747) );
INVx2_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g779 ( .A(n_732), .Y(n_779) );
NAND2xp33_ASAP7_75t_SL g733 ( .A(n_734), .B(n_735), .Y(n_733) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_743), .B1(n_744), .B2(n_746), .C(n_747), .Y(n_737) );
NOR4xp25_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .C(n_741), .D(n_742), .Y(n_738) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g781 ( .A1(n_749), .A2(n_782), .B(n_783), .Y(n_781) );
NAND4xp75_ASAP7_75t_L g749 ( .A(n_750), .B(n_764), .C(n_770), .D(n_776), .Y(n_749) );
INVx3_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g753 ( .A(n_754), .B(n_759), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NOR2x1_ASAP7_75t_L g770 ( .A(n_771), .B(n_774), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_784), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_787), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_796), .B(n_797), .Y(n_789) );
INVxp33_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND2x1_ASAP7_75t_SL g791 ( .A(n_792), .B(n_795), .Y(n_791) );
CKINVDCx11_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
OR3x1_ASAP7_75t_L g797 ( .A(n_798), .B(n_805), .C(n_809), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_798), .A2(n_813), .B(n_816), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
BUFx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
BUFx3_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
BUFx2_ASAP7_75t_R g815 ( .A(n_804), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
BUFx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_827), .Y(n_811) );
INVx1_ASAP7_75t_SL g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
XNOR2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_822), .B1(n_823), .B2(n_826), .Y(n_818) );
INVx1_ASAP7_75t_L g826 ( .A(n_819), .Y(n_826) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
CKINVDCx11_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
CKINVDCx8_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
endmodule