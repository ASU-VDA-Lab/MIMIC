module fake_jpeg_3271_n_593 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_593);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_593;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_80),
.Y(n_132)
);

BUFx6f_ASAP7_75t_SL g63 ( 
.A(n_57),
.Y(n_63)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_66),
.B(n_71),
.Y(n_135)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_18),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_72),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_20),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_75),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_78),
.Y(n_188)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_26),
.A2(n_0),
.B(n_1),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_83),
.A2(n_47),
.B(n_45),
.Y(n_127)
);

BUFx2_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g129 ( 
.A(n_84),
.B(n_121),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_89),
.Y(n_189)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_94),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_91),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_36),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_21),
.B(n_17),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_100),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_28),
.B(n_2),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_37),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_106),
.Y(n_149)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_37),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_109),
.B(n_117),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_112),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_116),
.Y(n_194)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_42),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_21),
.B(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_120),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_47),
.B(n_3),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_23),
.B(n_16),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_122),
.B(n_41),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_123),
.B(n_19),
.Y(n_192)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_46),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_39),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_127),
.A2(n_22),
.B(n_7),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_84),
.B(n_46),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_137),
.B(n_148),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_86),
.A2(n_59),
.B1(n_53),
.B2(n_40),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_138),
.A2(n_146),
.B1(n_162),
.B2(n_165),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_73),
.A2(n_59),
.B1(n_53),
.B2(n_58),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_142),
.A2(n_157),
.B1(n_174),
.B2(n_178),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_88),
.A2(n_58),
.B1(n_59),
.B2(n_43),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_144),
.A2(n_198),
.B1(n_110),
.B2(n_101),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_87),
.A2(n_58),
.B1(n_45),
.B2(n_43),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_64),
.B(n_50),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_68),
.B(n_55),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_153),
.B(n_154),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_67),
.B(n_50),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_76),
.A2(n_55),
.B1(n_52),
.B2(n_49),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_SL g160 ( 
.A(n_74),
.Y(n_160)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_160),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_97),
.A2(n_45),
.B1(n_43),
.B2(n_34),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_85),
.A2(n_103),
.B1(n_95),
.B2(n_72),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_78),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_173),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_70),
.A2(n_34),
.B1(n_33),
.B2(n_19),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_92),
.A2(n_41),
.B1(n_33),
.B2(n_34),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_79),
.A2(n_19),
.B1(n_33),
.B2(n_48),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_190),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_81),
.B(n_52),
.C(n_49),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_61),
.C(n_30),
.Y(n_211)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_75),
.B(n_48),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_91),
.B(n_44),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_200),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_192),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_93),
.A2(n_44),
.B1(n_39),
.B2(n_27),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_115),
.B(n_27),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_SL g203 ( 
.A1(n_123),
.A2(n_23),
.B(n_30),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_203),
.A2(n_25),
.B(n_9),
.Y(n_258)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_204),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_143),
.B(n_121),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_206),
.B(n_213),
.Y(n_278)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_140),
.Y(n_210)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_210),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_211),
.B(n_216),
.Y(n_284)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_212),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_150),
.B(n_116),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_145),
.Y(n_214)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_214),
.Y(n_290)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_215),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_102),
.Y(n_216)
);

BUFx12_ASAP7_75t_L g217 ( 
.A(n_156),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_217),
.Y(n_311)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_218),
.Y(n_331)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_135),
.B(n_105),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_220),
.B(n_227),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_129),
.B(n_114),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_221),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_142),
.A2(n_113),
.B1(n_112),
.B2(n_111),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_222),
.A2(n_275),
.B1(n_133),
.B2(n_179),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_132),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_223),
.B(n_228),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_224),
.A2(n_138),
.B1(n_146),
.B2(n_162),
.Y(n_285)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_126),
.Y(n_225)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_152),
.B(n_3),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_226),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_141),
.B(n_3),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_158),
.B(n_189),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_139),
.B(n_4),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_230),
.B(n_238),
.Y(n_315)
);

O2A1O1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_165),
.A2(n_30),
.B(n_22),
.C(n_7),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_231),
.A2(n_130),
.B(n_177),
.Y(n_309)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_232),
.Y(n_282)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_128),
.Y(n_233)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_30),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_252),
.C(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_170),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_235),
.Y(n_304)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_236),
.Y(n_312)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_180),
.Y(n_237)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_164),
.B(n_5),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_171),
.B(n_5),
.Y(n_239)
);

AOI21xp33_ASAP7_75t_L g322 ( 
.A1(n_239),
.A2(n_240),
.B(n_247),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_171),
.B(n_5),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_193),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_242),
.B(n_249),
.Y(n_325)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_147),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_245),
.Y(n_314)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_147),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_246),
.Y(n_324)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_176),
.Y(n_248)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_125),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_250),
.Y(n_318)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_251),
.Y(n_319)
);

AND2x2_ASAP7_75t_SL g252 ( 
.A(n_170),
.B(n_22),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_126),
.Y(n_253)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_133),
.Y(n_254)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_254),
.Y(n_328)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_155),
.Y(n_255)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_255),
.Y(n_335)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_155),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_256),
.B(n_257),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_136),
.B(n_6),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_258),
.A2(n_131),
.B(n_196),
.Y(n_305)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_163),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_259),
.B(n_260),
.Y(n_329)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_163),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_125),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_261),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_159),
.B(n_25),
.C(n_12),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_263),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g264 ( 
.A(n_176),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_264),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_170),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_265),
.A2(n_131),
.B1(n_187),
.B2(n_134),
.Y(n_299)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_161),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_266),
.Y(n_333)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_270),
.Y(n_288)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_161),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_188),
.B(n_7),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_273),
.Y(n_293)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_151),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_178),
.A2(n_25),
.B1(n_13),
.B2(n_14),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_234),
.B(n_187),
.C(n_151),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_281),
.B(n_292),
.C(n_298),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_285),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_229),
.A2(n_183),
.B1(n_174),
.B2(n_201),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_SL g292 ( 
.A(n_208),
.B(n_186),
.C(n_130),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_229),
.A2(n_201),
.B1(n_199),
.B2(n_197),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_224),
.A2(n_199),
.B1(n_197),
.B2(n_179),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_207),
.B(n_205),
.C(n_211),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_299),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_144),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_313),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_303),
.A2(n_326),
.B1(n_332),
.B2(n_248),
.Y(n_363)
);

OAI21xp33_ASAP7_75t_SL g337 ( 
.A1(n_305),
.A2(n_309),
.B(n_268),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_271),
.A2(n_169),
.B1(n_167),
.B2(n_196),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_310),
.A2(n_330),
.B1(n_225),
.B2(n_253),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_226),
.B(n_195),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_275),
.A2(n_169),
.B1(n_167),
.B2(n_134),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_316),
.A2(n_330),
.B1(n_309),
.B2(n_299),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g326 ( 
.A1(n_205),
.A2(n_177),
.B1(n_195),
.B2(n_25),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_222),
.A2(n_195),
.B1(n_13),
.B2(n_14),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_221),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_274),
.A2(n_12),
.B(n_15),
.C(n_16),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_334),
.B(n_269),
.Y(n_339)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_280),
.Y(n_336)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_336),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_337),
.B(n_361),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_310),
.A2(n_268),
.B1(n_252),
.B2(n_270),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_338),
.A2(n_344),
.B1(n_357),
.B2(n_363),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_339),
.A2(n_359),
.B(n_365),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_340),
.Y(n_386)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_288),
.Y(n_341)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_341),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_209),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_343),
.B(n_346),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_323),
.B(n_245),
.Y(n_346)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_280),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_348),
.Y(n_397)
);

MAJx2_ASAP7_75t_L g349 ( 
.A(n_298),
.B(n_252),
.C(n_268),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_360),
.Y(n_396)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_350),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_315),
.B(n_262),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_351),
.B(n_364),
.Y(n_418)
);

O2A1O1Ixp33_ASAP7_75t_L g352 ( 
.A1(n_302),
.A2(n_231),
.B(n_250),
.C(n_256),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_352),
.A2(n_324),
.B(n_314),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g353 ( 
.A(n_276),
.B(n_204),
.C(n_219),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_358),
.Y(n_387)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_354),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_293),
.B(n_232),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_355),
.B(n_362),
.Y(n_399)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_356),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_303),
.A2(n_266),
.B1(n_241),
.B2(n_237),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_325),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_291),
.A2(n_235),
.B1(n_265),
.B2(n_246),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_284),
.B(n_210),
.Y(n_360)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_329),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_289),
.B(n_215),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_267),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_366),
.B(n_370),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_278),
.B(n_243),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_372),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_278),
.A2(n_254),
.B1(n_243),
.B2(n_264),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_368),
.A2(n_304),
.B1(n_333),
.B2(n_328),
.Y(n_391)
);

AND2x2_ASAP7_75t_SL g369 ( 
.A(n_277),
.B(n_264),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_369),
.B(n_379),
.Y(n_421)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_297),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_305),
.A2(n_217),
.B(n_244),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_371),
.A2(n_378),
.B(n_312),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_293),
.B(n_12),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_321),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_380),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_311),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_374),
.B(n_375),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_312),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_301),
.B(n_15),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_376),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_322),
.A2(n_217),
.B(n_244),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_277),
.B(n_281),
.Y(n_379)
);

AO21x2_ASAP7_75t_L g380 ( 
.A1(n_294),
.A2(n_295),
.B(n_332),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_301),
.B(n_287),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_381),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g382 ( 
.A(n_334),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_382),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_345),
.A2(n_289),
.B1(n_296),
.B2(n_283),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_384),
.B(n_394),
.Y(n_425)
);

XOR2x2_ASAP7_75t_SL g388 ( 
.A(n_342),
.B(n_292),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_349),
.Y(n_423)
);

AOI322xp5_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_296),
.A3(n_313),
.B1(n_283),
.B2(n_311),
.C1(n_287),
.C2(n_333),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_389),
.A2(n_378),
.B(n_351),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_390),
.A2(n_419),
.B(n_420),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_391),
.A2(n_380),
.B1(n_344),
.B2(n_375),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_319),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_398),
.C(n_405),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_345),
.A2(n_328),
.B1(n_317),
.B2(n_319),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_335),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_380),
.A2(n_317),
.B1(n_335),
.B2(n_300),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_357),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_365),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_403),
.B(n_411),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_347),
.B(n_308),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_368),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_SL g412 ( 
.A(n_347),
.B(n_304),
.C(n_306),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_414),
.C(n_369),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_369),
.B(n_282),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_377),
.A2(n_306),
.B1(n_314),
.B2(n_324),
.Y(n_419)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_406),
.Y(n_422)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_422),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_423),
.B(n_396),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_426),
.B(n_398),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_446),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_358),
.C(n_341),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_428),
.B(n_455),
.C(n_424),
.Y(n_459)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_406),
.Y(n_429)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_429),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_410),
.A2(n_380),
.B1(n_350),
.B2(n_363),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_431),
.B1(n_437),
.B2(n_445),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_410),
.A2(n_380),
.B1(n_359),
.B2(n_367),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_415),
.Y(n_432)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_432),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_417),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_438),
.Y(n_465)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_415),
.Y(n_435)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_436),
.Y(n_471)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_399),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_413),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_439),
.B(n_440),
.Y(n_468)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_413),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_395),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_442),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_397),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_397),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_444),
.Y(n_464)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_395),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_416),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_447),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_400),
.B(n_355),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_449),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_420),
.A2(n_371),
.B(n_377),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_450),
.A2(n_409),
.B(n_390),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_364),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_451),
.Y(n_457)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_386),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_452),
.A2(n_453),
.B1(n_386),
.B2(n_354),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_408),
.B(n_372),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_392),
.A2(n_338),
.B1(n_352),
.B2(n_339),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_454),
.A2(n_392),
.B1(n_411),
.B2(n_394),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_421),
.B(n_365),
.C(n_356),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_459),
.B(n_481),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_460),
.B(n_450),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_424),
.B(n_393),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_472),
.C(n_474),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_426),
.B(n_405),
.C(n_412),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_428),
.B(n_396),
.C(n_414),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_480),
.C(n_483),
.Y(n_510)
);

AOI22x1_ASAP7_75t_L g476 ( 
.A1(n_431),
.A2(n_392),
.B1(n_402),
.B2(n_384),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_476),
.A2(n_477),
.B1(n_479),
.B2(n_385),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_478),
.A2(n_447),
.B(n_444),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_430),
.A2(n_385),
.B1(n_408),
.B2(n_418),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_423),
.B(n_388),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_409),
.Y(n_481)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_482),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_427),
.B(n_404),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_448),
.B(n_404),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_484),
.B(n_453),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_434),
.A2(n_419),
.B(n_387),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_485),
.B(n_448),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_464),
.B(n_442),
.Y(n_486)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_486),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_465),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_487),
.B(n_503),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_488),
.A2(n_500),
.B(n_505),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_461),
.A2(n_437),
.B1(n_425),
.B2(n_436),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_489),
.A2(n_494),
.B1(n_479),
.B2(n_477),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_491),
.B(n_495),
.Y(n_530)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_458),
.Y(n_493)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_493),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_461),
.A2(n_425),
.B1(n_438),
.B2(n_454),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_484),
.Y(n_496)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_496),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_480),
.B(n_434),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_498),
.B(n_499),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_459),
.B(n_449),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_501),
.A2(n_457),
.B1(n_471),
.B2(n_476),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_460),
.B(n_451),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_502),
.B(n_508),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_470),
.B(n_433),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_458),
.Y(n_504)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_504),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_478),
.A2(n_441),
.B(n_446),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_464),
.B(n_443),
.Y(n_506)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_506),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_473),
.B(n_422),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_507),
.B(n_511),
.Y(n_532)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_462),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_462),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_452),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_471),
.B(n_429),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_514),
.A2(n_529),
.B1(n_489),
.B2(n_494),
.Y(n_537)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_518),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_519),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_486),
.A2(n_485),
.B(n_463),
.Y(n_520)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_520),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_490),
.B(n_472),
.C(n_469),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_521),
.B(n_523),
.C(n_524),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_490),
.B(n_474),
.C(n_475),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_499),
.B(n_481),
.C(n_483),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_500),
.A2(n_476),
.B(n_468),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_525),
.A2(n_391),
.B(n_467),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_492),
.A2(n_445),
.B1(n_466),
.B2(n_456),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_497),
.B(n_440),
.C(n_439),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_531),
.B(n_506),
.C(n_510),
.Y(n_539)
);

AOI21xp33_ASAP7_75t_L g533 ( 
.A1(n_513),
.A2(n_505),
.B(n_507),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_533),
.A2(n_549),
.B(n_520),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_537),
.A2(n_544),
.B1(n_525),
.B2(n_519),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_531),
.B(n_497),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_538),
.B(n_540),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_539),
.B(n_521),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_523),
.B(n_524),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_527),
.B(n_383),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_541),
.B(n_545),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_512),
.B(n_511),
.Y(n_542)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_542),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_516),
.A2(n_488),
.B1(n_491),
.B2(n_510),
.Y(n_544)
);

FAx1_ASAP7_75t_SL g545 ( 
.A(n_530),
.B(n_498),
.CI(n_495),
.CON(n_545),
.SN(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_532),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_546),
.B(n_547),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_515),
.B(n_401),
.Y(n_547)
);

AOI21x1_ASAP7_75t_L g563 ( 
.A1(n_548),
.A2(n_522),
.B(n_532),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_515),
.A2(n_435),
.B(n_432),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_550),
.B(n_551),
.Y(n_571)
);

FAx1_ASAP7_75t_SL g552 ( 
.A(n_544),
.B(n_530),
.CI(n_502),
.CON(n_552),
.SN(n_552)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_552),
.B(n_560),
.Y(n_565)
);

AO21x1_ASAP7_75t_L g574 ( 
.A1(n_553),
.A2(n_562),
.B(n_545),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_543),
.A2(n_528),
.B(n_522),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_554),
.A2(n_563),
.B(n_548),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_543),
.A2(n_526),
.B(n_517),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_556),
.A2(n_542),
.B(n_535),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_539),
.B(n_540),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_559),
.B(n_534),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_538),
.B(n_514),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_537),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_558),
.B(n_534),
.Y(n_564)
);

OAI21x1_ASAP7_75t_SL g581 ( 
.A1(n_564),
.A2(n_566),
.B(n_568),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_567),
.B(n_569),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_555),
.A2(n_549),
.B(n_526),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_558),
.B(n_536),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_570),
.A2(n_574),
.B(n_373),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_SL g572 ( 
.A1(n_562),
.A2(n_536),
.B1(n_528),
.B2(n_529),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_572),
.A2(n_551),
.B1(n_557),
.B2(n_554),
.Y(n_575)
);

MAJx2_ASAP7_75t_L g573 ( 
.A(n_560),
.B(n_545),
.C(n_348),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_573),
.B(n_552),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_575),
.A2(n_340),
.B1(n_318),
.B2(n_308),
.Y(n_585)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_576),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_565),
.A2(n_561),
.B(n_336),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_577),
.A2(n_579),
.B(n_580),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_571),
.B(n_370),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_578),
.B(n_565),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_582),
.B(n_583),
.C(n_585),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_581),
.A2(n_362),
.B(n_318),
.Y(n_583)
);

NOR2xp67_ASAP7_75t_L g587 ( 
.A(n_584),
.B(n_586),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_587),
.A2(n_588),
.B1(n_279),
.B2(n_320),
.Y(n_590)
);

OAI311xp33_ASAP7_75t_L g588 ( 
.A1(n_582),
.A2(n_576),
.A3(n_282),
.B1(n_300),
.C1(n_320),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_590),
.A2(n_589),
.B(n_279),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_290),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_592),
.A2(n_290),
.B(n_331),
.Y(n_593)
);


endmodule