module fake_jpeg_31114_n_537 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_537);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_537;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_53),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_90),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_56),
.Y(n_151)
);

NAND2x1_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_37),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_57),
.B(n_63),
.Y(n_155)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_61),
.Y(n_156)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_17),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_66),
.Y(n_158)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_72),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_73),
.A2(n_46),
.B1(n_38),
.B2(n_45),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_81),
.Y(n_113)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_87),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_27),
.B(n_17),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_27),
.B(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_101),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_22),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_106),
.B(n_23),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_108),
.B(n_109),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_71),
.Y(n_116)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_63),
.B(n_50),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_129),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_57),
.B(n_19),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_82),
.B(n_19),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_157),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_91),
.A2(n_48),
.B1(n_34),
.B2(n_32),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_148),
.A2(n_68),
.B1(n_76),
.B2(n_67),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_71),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_149),
.B(n_152),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_84),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_48),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_83),
.B(n_23),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_162),
.A2(n_31),
.B1(n_35),
.B2(n_44),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_56),
.B(n_46),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_166),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_73),
.B(n_45),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_72),
.B(n_38),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_41),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_35),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_169),
.B(n_204),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_161),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_170),
.B(n_199),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_124),
.B(n_42),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_171),
.B(n_178),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g272 ( 
.A(n_172),
.Y(n_272)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_117),
.B(n_84),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_175),
.B(n_211),
.C(n_128),
.Y(n_258)
);

BUFx16f_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_176),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_177),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_42),
.Y(n_178)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_181),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_184),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_145),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_185),
.Y(n_238)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_186),
.Y(n_257)
);

CKINVDCx12_ASAP7_75t_R g187 ( 
.A(n_126),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_189),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_131),
.A2(n_105),
.B1(n_104),
.B2(n_98),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_190),
.A2(n_210),
.B1(n_128),
.B2(n_138),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_118),
.B(n_34),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_192),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_48),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_126),
.B(n_48),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_198),
.Y(n_242)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_197),
.Y(n_261)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_134),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_120),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_120),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_200),
.B(n_203),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_201),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_202),
.A2(n_158),
.B1(n_156),
.B2(n_119),
.Y(n_260)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_125),
.B(n_31),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_206),
.B(n_209),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_115),
.B(n_53),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_208),
.B(n_222),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_148),
.A2(n_99),
.B1(n_102),
.B2(n_78),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_96),
.C(n_59),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_114),
.B(n_43),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_216),
.Y(n_249)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_226),
.B1(n_141),
.B2(n_140),
.Y(n_239)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_139),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_218),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_114),
.B(n_43),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_217),
.A2(n_44),
.B1(n_95),
.B2(n_94),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_116),
.Y(n_218)
);

BUFx12_ASAP7_75t_L g219 ( 
.A(n_135),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_219),
.Y(n_229)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_220),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_140),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_221),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_115),
.B(n_60),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_223),
.B(n_224),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_114),
.B(n_48),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_123),
.B(n_66),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_225),
.B(n_227),
.Y(n_268)
);

CKINVDCx12_ASAP7_75t_R g226 ( 
.A(n_140),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_123),
.B(n_61),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_167),
.B1(n_165),
.B2(n_138),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_231),
.A2(n_233),
.B1(n_253),
.B2(n_260),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_245),
.A2(n_247),
.B1(n_252),
.B2(n_262),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_207),
.A2(n_133),
.B1(n_147),
.B2(n_77),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_199),
.A2(n_56),
.B(n_64),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_250),
.A2(n_208),
.B(n_225),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_169),
.A2(n_79),
.B1(n_88),
.B2(n_159),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_210),
.A2(n_165),
.B1(n_54),
.B2(n_146),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g255 ( 
.A1(n_204),
.A2(n_64),
.B(n_146),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_258),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_180),
.A2(n_158),
.B1(n_156),
.B2(n_119),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_194),
.A2(n_136),
.B1(n_141),
.B2(n_69),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_264),
.A2(n_233),
.B1(n_253),
.B2(n_272),
.Y(n_314)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_175),
.B(n_145),
.Y(n_266)
);

OR2x4_ASAP7_75t_L g309 ( 
.A(n_266),
.B(n_176),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_199),
.B(n_179),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_269),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_211),
.B(n_151),
.C(n_122),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_237),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_275),
.B(n_278),
.Y(n_328)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_277),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_183),
.Y(n_278)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_234),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_279),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_240),
.B(n_249),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_281),
.B(n_282),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_184),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_256),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_283),
.B(n_285),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_173),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_286),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_205),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_256),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_208),
.Y(n_289)
);

FAx1_ASAP7_75t_SL g318 ( 
.A(n_289),
.B(n_292),
.CI(n_267),
.CON(n_318),
.SN(n_318)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_296),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_268),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_260),
.A2(n_181),
.B1(n_188),
.B2(n_201),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_293),
.A2(n_304),
.B(n_313),
.Y(n_347)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_222),
.B1(n_227),
.B2(n_225),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_295),
.A2(n_306),
.B1(n_271),
.B2(n_238),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_241),
.B(n_175),
.Y(n_296)
);

INVx4_ASAP7_75t_SL g298 ( 
.A(n_244),
.Y(n_298)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_299),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_300),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_186),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_310),
.Y(n_325)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_229),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_302),
.Y(n_349)
);

OAI32xp33_ASAP7_75t_L g303 ( 
.A1(n_247),
.A2(n_220),
.A3(n_80),
.B1(n_222),
.B2(n_189),
.Y(n_303)
);

OAI32xp33_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_262),
.A3(n_309),
.B1(n_313),
.B2(n_266),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_255),
.A2(n_170),
.B(n_227),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_305),
.A2(n_265),
.B(n_251),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_268),
.A2(n_172),
.B1(n_193),
.B2(n_136),
.Y(n_306)
);

INVx13_ASAP7_75t_L g307 ( 
.A(n_234),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_307),
.Y(n_322)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_243),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_308),
.Y(n_342)
);

NAND2xp33_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_274),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_197),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_230),
.B(n_203),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_315),
.Y(n_327)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_229),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_312),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g313 ( 
.A(n_255),
.B(n_70),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_297),
.B1(n_280),
.B2(n_245),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_242),
.B(n_206),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_316),
.A2(n_336),
.B1(n_244),
.B2(n_263),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_330),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_287),
.A2(n_250),
.B(n_265),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_319),
.A2(n_259),
.B(n_185),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_324),
.A2(n_343),
.B1(n_306),
.B2(n_291),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_326),
.A2(n_319),
.B(n_304),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_274),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_305),
.A2(n_176),
.B(n_265),
.C(n_272),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_SL g379 ( 
.A(n_332),
.B(n_333),
.C(n_298),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_287),
.A2(n_274),
.B1(n_271),
.B2(n_235),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_288),
.B(n_228),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_301),
.C(n_289),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_310),
.B(n_236),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_345),
.Y(n_376)
);

AO22x1_ASAP7_75t_L g341 ( 
.A1(n_303),
.A2(n_280),
.B1(n_289),
.B2(n_295),
.Y(n_341)
);

O2A1O1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_341),
.A2(n_346),
.B(n_263),
.C(n_257),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_280),
.A2(n_272),
.B1(n_232),
.B2(n_236),
.Y(n_343)
);

XNOR2x1_ASAP7_75t_SL g344 ( 
.A(n_292),
.B(n_228),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_352),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_288),
.B(n_238),
.Y(n_345)
);

AO21x2_ASAP7_75t_L g346 ( 
.A1(n_275),
.A2(n_238),
.B(n_232),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g352 ( 
.A(n_292),
.B(n_248),
.C(n_219),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_328),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_353),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_286),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_355),
.B(n_357),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_356),
.B(n_366),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_329),
.B(n_312),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_321),
.Y(n_358)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_359),
.Y(n_388)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_331),
.Y(n_360)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_327),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_365),
.Y(n_397)
);

AND2x6_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_290),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_339),
.Y(n_367)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_367),
.Y(n_396)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_350),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_369),
.A2(n_324),
.B1(n_316),
.B2(n_332),
.Y(n_391)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

OAI32xp33_ASAP7_75t_L g371 ( 
.A1(n_341),
.A2(n_291),
.A3(n_302),
.B1(n_257),
.B2(n_259),
.Y(n_371)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_371),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g372 ( 
.A(n_327),
.B(n_15),
.C(n_12),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_373),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_340),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_326),
.A2(n_248),
.B(n_300),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_374),
.A2(n_379),
.B(n_378),
.Y(n_393)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_351),
.Y(n_375)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_375),
.Y(n_413)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_350),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_380),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_381),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_317),
.B(n_277),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_317),
.B(n_299),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_385),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_383),
.A2(n_386),
.B1(n_334),
.B2(n_332),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_384),
.A2(n_374),
.B(n_346),
.Y(n_405)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_343),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_336),
.A2(n_213),
.B1(n_195),
.B2(n_174),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_353),
.B(n_320),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_390),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_391),
.A2(n_403),
.B1(n_386),
.B2(n_356),
.Y(n_422)
);

OAI21xp33_ASAP7_75t_L g392 ( 
.A1(n_379),
.A2(n_320),
.B(n_344),
.Y(n_392)
);

HAxp5_ASAP7_75t_SL g428 ( 
.A(n_392),
.B(n_354),
.CON(n_428),
.SN(n_428)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_393),
.A2(n_410),
.B(n_346),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_367),
.B(n_325),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_404),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_401),
.A2(n_337),
.B1(n_368),
.B2(n_377),
.Y(n_441)
);

OAI32xp33_ASAP7_75t_L g402 ( 
.A1(n_385),
.A2(n_325),
.A3(n_330),
.B1(n_345),
.B2(n_346),
.Y(n_402)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_402),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_381),
.A2(n_323),
.B1(n_322),
.B2(n_332),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_382),
.B(n_376),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_405),
.A2(n_346),
.B(n_371),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_361),
.A2(n_332),
.B(n_347),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_348),
.Y(n_415)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_415),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_354),
.B(n_362),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_416),
.B(n_337),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_361),
.A2(n_347),
.B1(n_352),
.B2(n_349),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_410),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_393),
.A2(n_383),
.B(n_384),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g460 ( 
.A(n_418),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_421),
.B(n_443),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_422),
.A2(n_428),
.B1(n_440),
.B2(n_444),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_366),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_423),
.B(n_439),
.Y(n_451)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_416),
.Y(n_425)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_425),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_342),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_431),
.Y(n_459)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_387),
.Y(n_427)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_401),
.A2(n_369),
.B1(n_365),
.B2(n_363),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_434),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_338),
.C(n_363),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_435),
.C(n_438),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_360),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_437),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_318),
.C(n_375),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_397),
.A2(n_359),
.B1(n_358),
.B2(n_370),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_436),
.A2(n_408),
.B1(n_396),
.B2(n_405),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_395),
.B(n_409),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_318),
.C(n_323),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_307),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_441),
.A2(n_413),
.B1(n_407),
.B2(n_388),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_442),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_390),
.B(n_17),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_414),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_450),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_391),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_448),
.B(n_428),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_424),
.A2(n_396),
.B1(n_389),
.B2(n_394),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_398),
.C(n_406),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_455),
.C(n_464),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_430),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_454),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_406),
.C(n_404),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_389),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_394),
.C(n_388),
.Y(n_457)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_457),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_400),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_461),
.B(n_439),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_429),
.B(n_440),
.C(n_441),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_440),
.B(n_400),
.C(n_413),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_466),
.B(n_420),
.C(n_418),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_465),
.A2(n_434),
.B(n_421),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_467),
.A2(n_475),
.B(n_477),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_468),
.B(n_473),
.Y(n_489)
);

AO21x1_ASAP7_75t_L g469 ( 
.A1(n_460),
.A2(n_420),
.B(n_419),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_472),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_465),
.A2(n_419),
.B(n_430),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_447),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_478),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_427),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_445),
.Y(n_484)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_463),
.A2(n_444),
.B1(n_407),
.B2(n_387),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_479),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_130),
.Y(n_496)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_462),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_482),
.B(n_483),
.Y(n_486)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_459),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_484),
.B(n_496),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_479),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_485),
.B(n_13),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_474),
.A2(n_452),
.B(n_466),
.Y(n_487)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_487),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_480),
.A2(n_449),
.B1(n_461),
.B2(n_448),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_491),
.A2(n_471),
.B1(n_473),
.B2(n_469),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_453),
.C(n_455),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_494),
.C(n_495),
.Y(n_505)
);

OAI321xp33_ASAP7_75t_L g493 ( 
.A1(n_467),
.A2(n_456),
.A3(n_464),
.B1(n_451),
.B2(n_411),
.C(n_452),
.Y(n_493)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_493),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_470),
.B(n_451),
.C(n_177),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_472),
.B(n_279),
.C(n_122),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_497),
.A2(n_130),
.B(n_143),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_468),
.B(n_219),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_498),
.B(n_475),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_502),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_488),
.A2(n_481),
.B(n_206),
.Y(n_504)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_504),
.Y(n_515)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_506),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_486),
.B(n_14),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_507),
.B(n_508),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_494),
.C(n_496),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_499),
.B(n_12),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_510),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_490),
.A2(n_16),
.B(n_215),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_511),
.A2(n_490),
.B(n_495),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_514),
.B(n_518),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_512),
.A2(n_484),
.B1(n_489),
.B2(n_32),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_503),
.A2(n_489),
.B1(n_32),
.B2(n_143),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_521),
.C(n_511),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_505),
.A2(n_103),
.B1(n_80),
.B2(n_65),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_525),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_515),
.A2(n_510),
.B1(n_505),
.B2(n_508),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_523),
.A2(n_527),
.B1(n_519),
.B2(n_516),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_500),
.C(n_41),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_514),
.A2(n_500),
.B(n_215),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_526),
.A2(n_516),
.B(n_513),
.Y(n_529)
);

AOI322xp5_ASAP7_75t_L g527 ( 
.A1(n_513),
.A2(n_0),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_529),
.C(n_524),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_532),
.B(n_5),
.Y(n_533)
);

AOI322xp5_ASAP7_75t_L g532 ( 
.A1(n_530),
.A2(n_527),
.A3(n_41),
.B1(n_6),
.B2(n_7),
.C1(n_4),
.C2(n_10),
.Y(n_532)
);

AOI322xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C1(n_11),
.C2(n_412),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_7),
.B(n_8),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_535),
.B(n_8),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_536),
.B(n_10),
.Y(n_537)
);


endmodule