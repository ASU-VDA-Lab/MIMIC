module fake_jpeg_2219_n_201 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_201);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_59),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g88 ( 
.A(n_76),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_82),
.Y(n_84)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_92),
.C(n_1),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_65),
.B1(n_51),
.B2(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_78),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_65),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_78),
.C(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_93),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_52),
.B1(n_53),
.B2(n_68),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_53),
.B1(n_68),
.B2(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_66),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_109),
.B1(n_114),
.B2(n_105),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_100),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_76),
.C(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_68),
.B1(n_53),
.B2(n_76),
.Y(n_102)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_102),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_107),
.Y(n_122)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_88),
.Y(n_123)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_114),
.Y(n_117)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_77),
.B1(n_64),
.B2(n_60),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_73),
.B1(n_64),
.B2(n_70),
.Y(n_132)
);

NOR2xp67_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_85),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_58),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_119),
.B(n_7),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_136),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_87),
.C(n_77),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_131),
.C(n_40),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_2),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_73),
.C(n_71),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_113),
.B1(n_70),
.B2(n_6),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_2),
.Y(n_136)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_112),
.B(n_71),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_33),
.B(n_30),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_3),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_141),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_137),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_3),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_145),
.Y(n_171)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_151),
.B1(n_154),
.B2(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_46),
.C(n_41),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_150),
.C(n_127),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_149),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_4),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_5),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_39),
.B1(n_38),
.B2(n_36),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_5),
.B(n_6),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_157),
.B(n_14),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_116),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_160),
.C(n_8),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_156),
.B(n_159),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

AOI322xp5_ASAP7_75t_SL g180 ( 
.A1(n_164),
.A2(n_165),
.A3(n_168),
.B1(n_173),
.B2(n_176),
.C1(n_152),
.C2(n_154),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_158),
.A2(n_120),
.B(n_128),
.C(n_126),
.D(n_29),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_126),
.B(n_9),
.C(n_10),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_175),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_27),
.B(n_26),
.C(n_25),
.D(n_23),
.Y(n_168)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_138),
.C(n_151),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_157),
.C(n_153),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_SL g173 ( 
.A(n_146),
.B(n_10),
.C(n_11),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_12),
.B(n_13),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_162),
.Y(n_189)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_178),
.A2(n_175),
.B1(n_162),
.B2(n_169),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_SL g186 ( 
.A(n_180),
.B(n_167),
.C(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_189),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_161),
.B(n_165),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_188),
.B(n_190),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_22),
.B(n_17),
.C(n_18),
.D(n_19),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_179),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_195),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_185),
.B1(n_178),
.B2(n_177),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_186),
.Y(n_196)
);

AOI221xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_192),
.B1(n_194),
.B2(n_18),
.C(n_19),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_197),
.B(n_17),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_21),
.B(n_15),
.Y(n_200)
);

AOI221xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_15),
.B1(n_20),
.B2(n_21),
.C(n_179),
.Y(n_201)
);


endmodule