module fake_netlist_6_2448_n_28 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_8, n_28);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_8;

output n_28;

wire n_16;
wire n_10;
wire n_21;
wire n_24;
wire n_18;
wire n_15;
wire n_27;
wire n_14;
wire n_22;
wire n_26;
wire n_13;
wire n_11;
wire n_17;
wire n_23;
wire n_12;
wire n_20;
wire n_19;
wire n_25;

AND2x2_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_4),
.Y(n_10)
);

AOI22xp33_ASAP7_75t_L g11 ( 
.A1(n_9),
.A2(n_2),
.B1(n_3),
.B2(n_8),
.Y(n_11)
);

OR2x2_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_4),
.Y(n_12)
);

OAI21xp33_ASAP7_75t_L g13 ( 
.A1(n_5),
.A2(n_6),
.B(n_2),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_6),
.Y(n_17)
);

AO31x2_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_0),
.A3(n_13),
.B(n_10),
.Y(n_18)
);

AO21x2_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_13),
.B(n_12),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

NAND4xp25_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_17),
.C(n_16),
.D(n_12),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_16),
.B(n_15),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_19),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_19),
.B1(n_10),
.B2(n_21),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_19),
.B1(n_11),
.B2(n_12),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_18),
.B1(n_25),
.B2(n_17),
.Y(n_28)
);


endmodule