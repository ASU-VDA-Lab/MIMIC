module fake_jpeg_17517_n_85 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_85);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_85;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx14_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_2),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_12),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_24),
.Y(n_32)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_18),
.B1(n_22),
.B2(n_16),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_39),
.B1(n_27),
.B2(n_1),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_19),
.C(n_8),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_15),
.B1(n_21),
.B2(n_20),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_40),
.B1(n_31),
.B2(n_25),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_16),
.B1(n_13),
.B2(n_9),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_21),
.B(n_19),
.C(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_47),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_50),
.B1(n_42),
.B2(n_21),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_31),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_53),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_28),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_27),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_37),
.C(n_32),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_56),
.C(n_28),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_28),
.C(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_53),
.B1(n_50),
.B2(n_44),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_40),
.B(n_49),
.Y(n_65)
);

AOI221xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_59),
.B1(n_55),
.B2(n_45),
.C(n_28),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_54),
.C(n_55),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_70),
.B(n_71),
.Y(n_75)
);

OAI322xp33_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_65),
.A3(n_68),
.B1(n_64),
.B2(n_28),
.C1(n_45),
.C2(n_10),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_73),
.A2(n_72),
.B(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_0),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_10),
.C(n_5),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_78),
.B(n_0),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_5),
.B1(n_1),
.B2(n_2),
.Y(n_80)
);

AO21x1_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_81),
.B(n_4),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g84 ( 
.A(n_83),
.B(n_4),
.CI(n_77),
.CON(n_84),
.SN(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_82),
.Y(n_85)
);


endmodule