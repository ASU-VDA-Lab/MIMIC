module fake_netlist_1_10515_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
CKINVDCx5p33_ASAP7_75t_R g3 ( .A(n_2), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
CKINVDCx11_ASAP7_75t_R g5 ( .A(n_4), .Y(n_5) );
BUFx3_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
OAI21x1_ASAP7_75t_L g7 ( .A1(n_6), .A2(n_3), .B(n_0), .Y(n_7) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
AOI22xp33_ASAP7_75t_L g10 ( .A1(n_7), .A2(n_5), .B1(n_0), .B2(n_1), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
OAI21xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_10), .B(n_1), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
endmodule