module fake_jpeg_10181_n_169 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

AOI21xp33_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_5),
.B(n_8),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_22),
.A2(n_11),
.B1(n_12),
.B2(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_20),
.B1(n_12),
.B2(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_37),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_9),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_12),
.B1(n_23),
.B2(n_20),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_20),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_21),
.B1(n_17),
.B2(n_11),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_21),
.B1(n_11),
.B2(n_16),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_21),
.B(n_36),
.C(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_58),
.B(n_60),
.Y(n_77)
);

BUFx24_ASAP7_75t_SL g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_60),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_65),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_67),
.B1(n_44),
.B2(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_39),
.B1(n_36),
.B2(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_55),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_28),
.B(n_29),
.Y(n_90)
);

AO22x1_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_45),
.B1(n_51),
.B2(n_54),
.Y(n_71)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_16),
.B1(n_19),
.B2(n_35),
.Y(n_92)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_75),
.B1(n_76),
.B2(n_47),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_45),
.B1(n_36),
.B2(n_34),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_64),
.B1(n_31),
.B2(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_80),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_45),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_64),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_50),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_24),
.C(n_26),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_86),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_88),
.Y(n_101)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_28),
.CI(n_38),
.CON(n_88),
.SN(n_88)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_7),
.B(n_6),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_92),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_70),
.Y(n_104)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_95),
.Y(n_99)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_96),
.B(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_108),
.C(n_88),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_81),
.B1(n_76),
.B2(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_66),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_79),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_74),
.B1(n_66),
.B2(n_55),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_95),
.B1(n_87),
.B2(n_83),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_118),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_122),
.B1(n_100),
.B2(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_121),
.C(n_38),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_88),
.B1(n_86),
.B2(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_86),
.B(n_48),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_103),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_104),
.C(n_98),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_56),
.B1(n_48),
.B2(n_16),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_131),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_103),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_114),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_113),
.B1(n_116),
.B2(n_120),
.Y(n_135)
);

NOR4xp25_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_48),
.C(n_6),
.D(n_5),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_56),
.C(n_24),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_133),
.C(n_35),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_38),
.C(n_35),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_128),
.B(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_141),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_138),
.C(n_19),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_118),
.B(n_122),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_16),
.C(n_1),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_127),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_139),
.A2(n_125),
.B1(n_133),
.B2(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_140),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_149),
.C(n_16),
.Y(n_155)
);

NOR4xp25_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_5),
.C(n_6),
.D(n_2),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_147),
.B(n_150),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_35),
.C(n_29),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_153),
.B(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_0),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_148),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_155),
.A2(n_150),
.B(n_1),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_157),
.A2(n_156),
.B1(n_2),
.B2(n_3),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_0),
.B(n_1),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_1),
.B(n_2),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_161),
.B(n_162),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_159),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_160),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_3),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_165),
.B1(n_4),
.B2(n_14),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_4),
.C(n_14),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_168),
.B(n_4),
.Y(n_169)
);


endmodule