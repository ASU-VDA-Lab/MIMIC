module real_aes_564_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g530 ( .A(n_0), .B(n_147), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_1), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_2), .B(n_129), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_3), .B(n_145), .Y(n_164) );
INVx1_ASAP7_75t_L g136 ( .A(n_4), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_5), .B(n_129), .Y(n_461) );
NAND2xp33_ASAP7_75t_SL g515 ( .A(n_6), .B(n_135), .Y(n_515) );
INVx1_ASAP7_75t_L g508 ( .A(n_7), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_8), .Y(n_106) );
AND2x2_ASAP7_75t_L g459 ( .A(n_9), .B(n_150), .Y(n_459) );
AND2x2_ASAP7_75t_L g166 ( .A(n_10), .B(n_154), .Y(n_166) );
AND2x2_ASAP7_75t_L g175 ( .A(n_11), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g151 ( .A(n_12), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_13), .B(n_145), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_14), .Y(n_110) );
AOI221x1_ASAP7_75t_L g511 ( .A1(n_15), .A2(n_138), .B1(n_176), .B2(n_512), .C(n_514), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_16), .B(n_129), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_17), .B(n_129), .Y(n_209) );
INVx1_ASAP7_75t_L g114 ( .A(n_18), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_19), .A2(n_86), .B1(n_129), .B2(n_239), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_20), .A2(n_138), .B(n_463), .Y(n_462) );
AOI221xp5_ASAP7_75t_SL g520 ( .A1(n_21), .A2(n_34), .B1(n_129), .B2(n_138), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_22), .B(n_147), .Y(n_464) );
OR2x2_ASAP7_75t_L g152 ( .A(n_23), .B(n_85), .Y(n_152) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_23), .A2(n_85), .B(n_151), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_24), .B(n_145), .Y(n_502) );
INVxp67_ASAP7_75t_L g510 ( .A(n_25), .Y(n_510) );
AND2x2_ASAP7_75t_L g483 ( .A(n_26), .B(n_149), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_27), .A2(n_138), .B(n_529), .Y(n_528) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_28), .A2(n_176), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_29), .B(n_145), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_30), .A2(n_138), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_31), .B(n_145), .Y(n_193) );
AND2x2_ASAP7_75t_L g135 ( .A(n_32), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g139 ( .A(n_32), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g247 ( .A(n_32), .Y(n_247) );
OR2x6_ASAP7_75t_L g112 ( .A(n_33), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_35), .B(n_129), .Y(n_165) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_36), .A2(n_78), .B1(n_138), .B2(n_245), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_37), .B(n_145), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_38), .B(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_39), .B(n_147), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_40), .A2(n_138), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_41), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g533 ( .A(n_42), .B(n_149), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_43), .B(n_149), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_44), .B(n_129), .Y(n_181) );
INVx1_ASAP7_75t_L g132 ( .A(n_45), .Y(n_132) );
INVx1_ASAP7_75t_L g142 ( .A(n_45), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_46), .B(n_145), .Y(n_173) );
AND2x2_ASAP7_75t_L g200 ( .A(n_47), .B(n_149), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_48), .B(n_129), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_49), .B(n_147), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_50), .B(n_147), .Y(n_192) );
AND2x2_ASAP7_75t_L g474 ( .A(n_51), .B(n_149), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_52), .B(n_129), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_53), .B(n_145), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_54), .B(n_129), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_55), .A2(n_138), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_56), .B(n_147), .Y(n_472) );
AND2x2_ASAP7_75t_SL g503 ( .A(n_57), .B(n_150), .Y(n_503) );
AND2x2_ASAP7_75t_L g215 ( .A(n_58), .B(n_150), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_59), .A2(n_138), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_60), .B(n_145), .Y(n_465) );
AND2x2_ASAP7_75t_SL g493 ( .A(n_61), .B(n_154), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_62), .B(n_147), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_63), .B(n_147), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_64), .A2(n_89), .B1(n_138), .B2(n_245), .Y(n_244) );
AOI221x1_ASAP7_75t_L g117 ( .A1(n_65), .A2(n_118), .B1(n_727), .B2(n_728), .C(n_730), .Y(n_117) );
CKINVDCx14_ASAP7_75t_R g727 ( .A(n_65), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_66), .B(n_145), .Y(n_212) );
INVx1_ASAP7_75t_L g134 ( .A(n_67), .Y(n_134) );
INVx1_ASAP7_75t_L g140 ( .A(n_67), .Y(n_140) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_68), .A2(n_99), .B1(n_116), .B2(n_733), .C1(n_737), .C2(n_748), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_68), .A2(n_729), .B1(n_743), .B2(n_744), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_68), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_69), .B(n_147), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_70), .A2(n_138), .B(n_204), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_71), .A2(n_138), .B(n_143), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_72), .A2(n_138), .B(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g195 ( .A(n_73), .B(n_150), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_74), .B(n_149), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_75), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_76), .B(n_129), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_77), .A2(n_80), .B1(n_129), .B2(n_239), .Y(n_491) );
INVx1_ASAP7_75t_L g115 ( .A(n_79), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_81), .B(n_147), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_82), .B(n_147), .Y(n_523) );
AND2x2_ASAP7_75t_L g153 ( .A(n_83), .B(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_84), .A2(n_138), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_87), .B(n_145), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_88), .A2(n_138), .B(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_90), .B(n_145), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_91), .Y(n_739) );
BUFx2_ASAP7_75t_L g214 ( .A(n_92), .Y(n_214) );
INVxp67_ASAP7_75t_L g513 ( .A(n_93), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_94), .B(n_145), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_95), .A2(n_138), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_96), .B(n_129), .Y(n_532) );
BUFx2_ASAP7_75t_L g107 ( .A(n_97), .Y(n_107) );
BUFx2_ASAP7_75t_SL g752 ( .A(n_97), .Y(n_752) );
INVx1_ASAP7_75t_SL g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_108), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_SL g736 ( .A(n_105), .B(n_107), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_105), .A2(n_750), .B(n_753), .Y(n_749) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g740 ( .A(n_109), .Y(n_740) );
BUFx3_ASAP7_75t_L g747 ( .A(n_109), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x6_ASAP7_75t_SL g448 ( .A(n_110), .B(n_111), .Y(n_448) );
AND2x6_ASAP7_75t_SL g450 ( .A(n_110), .B(n_112), .Y(n_450) );
OR2x2_ASAP7_75t_L g732 ( .A(n_110), .B(n_112), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVxp33_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21x1_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_446), .B(n_449), .Y(n_118) );
AO22x2_ASAP7_75t_L g728 ( .A1(n_119), .A2(n_447), .B1(n_450), .B2(n_729), .Y(n_728) );
INVx4_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_354), .Y(n_120) );
NOR3xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_277), .C(n_312), .Y(n_121) );
OAI211xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_177), .B(n_229), .C(n_267), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_156), .Y(n_124) );
AND2x2_ASAP7_75t_L g260 ( .A(n_125), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_125), .B(n_266), .Y(n_300) );
AND2x2_ASAP7_75t_L g325 ( .A(n_125), .B(n_280), .Y(n_325) );
INVx4_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx2_ASAP7_75t_L g232 ( .A(n_126), .Y(n_232) );
OR2x2_ASAP7_75t_L g263 ( .A(n_126), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g271 ( .A(n_126), .B(n_167), .Y(n_271) );
AND2x2_ASAP7_75t_L g279 ( .A(n_126), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g306 ( .A(n_126), .B(n_307), .Y(n_306) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_126), .B(n_309), .Y(n_317) );
AND2x4_ASAP7_75t_L g334 ( .A(n_126), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g372 ( .A(n_126), .Y(n_372) );
AND2x4_ASAP7_75t_SL g377 ( .A(n_126), .B(n_157), .Y(n_377) );
OR2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_153), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_137), .B(n_149), .Y(n_127) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_135), .Y(n_129) );
INVx1_ASAP7_75t_L g516 ( .A(n_130), .Y(n_516) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
AND2x6_ASAP7_75t_L g147 ( .A(n_131), .B(n_140), .Y(n_147) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g145 ( .A(n_133), .B(n_142), .Y(n_145) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx5_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
AND2x2_ASAP7_75t_L g141 ( .A(n_136), .B(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_136), .Y(n_242) );
AND2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
BUFx3_ASAP7_75t_L g243 ( .A(n_139), .Y(n_243) );
INVx2_ASAP7_75t_L g249 ( .A(n_140), .Y(n_249) );
AND2x4_ASAP7_75t_L g245 ( .A(n_141), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g241 ( .A(n_142), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_146), .B(n_148), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_147), .B(n_214), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_148), .A2(n_163), .B(n_164), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_148), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_148), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_148), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_148), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_148), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_148), .A2(n_464), .B(n_465), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_148), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_148), .A2(n_480), .B(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_148), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_148), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_148), .A2(n_530), .B(n_531), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_149), .Y(n_159) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_149), .A2(n_238), .B(n_244), .Y(n_237) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_149), .A2(n_520), .B(n_524), .Y(n_519) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x4_ASAP7_75t_L g186 ( .A(n_151), .B(n_152), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_154), .A2(n_209), .B(n_210), .Y(n_208) );
INVx2_ASAP7_75t_SL g489 ( .A(n_154), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_154), .A2(n_498), .B(n_499), .Y(n_497) );
BUFx4f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g168 ( .A(n_155), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_156), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_156), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_167), .Y(n_156) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_157), .Y(n_272) );
INVx2_ASAP7_75t_L g308 ( .A(n_157), .Y(n_308) );
INVx1_ASAP7_75t_L g335 ( .A(n_157), .Y(n_335) );
AND2x2_ASAP7_75t_L g434 ( .A(n_157), .B(n_344), .Y(n_434) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_158), .Y(n_266) );
AND2x2_ASAP7_75t_L g280 ( .A(n_158), .B(n_167), .Y(n_280) );
AOI21x1_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_166), .Y(n_158) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_159), .A2(n_468), .B(n_474), .Y(n_467) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_159), .A2(n_477), .B(n_483), .Y(n_476) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_159), .A2(n_477), .B(n_483), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_165), .Y(n_160) );
INVx2_ASAP7_75t_L g309 ( .A(n_167), .Y(n_309) );
INVx2_ASAP7_75t_L g344 ( .A(n_167), .Y(n_344) );
OR2x2_ASAP7_75t_L g429 ( .A(n_167), .B(n_261), .Y(n_429) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_175), .Y(n_167) );
INVx4_ASAP7_75t_L g176 ( .A(n_168), .Y(n_176) );
AOI21x1_ASAP7_75t_L g526 ( .A1(n_168), .A2(n_527), .B(n_533), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_174), .Y(n_169) );
INVx3_ASAP7_75t_L g188 ( .A(n_176), .Y(n_188) );
AOI211xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_196), .B(n_216), .C(n_223), .Y(n_177) );
INVx2_ASAP7_75t_SL g318 ( .A(n_178), .Y(n_318) );
AND2x2_ASAP7_75t_L g324 ( .A(n_178), .B(n_197), .Y(n_324) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_187), .Y(n_178) );
INVx1_ASAP7_75t_L g220 ( .A(n_179), .Y(n_220) );
INVx1_ASAP7_75t_L g226 ( .A(n_179), .Y(n_226) );
INVx2_ASAP7_75t_L g251 ( .A(n_179), .Y(n_251) );
AND2x2_ASAP7_75t_L g275 ( .A(n_179), .B(n_199), .Y(n_275) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_179), .Y(n_304) );
OR2x2_ASAP7_75t_L g384 ( .A(n_179), .B(n_207), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_186), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_186), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_186), .A2(n_461), .B(n_462), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_186), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_186), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_186), .B(n_513), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_186), .B(n_515), .C(n_516), .Y(n_514) );
AND2x2_ASAP7_75t_L g250 ( .A(n_187), .B(n_251), .Y(n_250) );
NOR2x1_ASAP7_75t_SL g282 ( .A(n_187), .B(n_207), .Y(n_282) );
AO21x1_ASAP7_75t_SL g187 ( .A1(n_188), .A2(n_189), .B(n_195), .Y(n_187) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_188), .A2(n_189), .B(n_195), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_194), .Y(n_189) );
INVxp67_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g296 ( .A(n_197), .B(n_219), .Y(n_296) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_207), .Y(n_197) );
OR2x2_ASAP7_75t_L g228 ( .A(n_198), .B(n_207), .Y(n_228) );
BUFx2_ASAP7_75t_L g252 ( .A(n_198), .Y(n_252) );
NOR2xp67_ASAP7_75t_L g303 ( .A(n_198), .B(n_304), .Y(n_303) );
INVx4_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_199), .Y(n_255) );
AND2x2_ASAP7_75t_L g281 ( .A(n_199), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g291 ( .A(n_199), .Y(n_291) );
NAND2x1_ASAP7_75t_L g329 ( .A(n_199), .B(n_207), .Y(n_329) );
OR2x2_ASAP7_75t_L g404 ( .A(n_199), .B(n_221), .Y(n_404) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx2_ASAP7_75t_SL g217 ( .A(n_207), .Y(n_217) );
AND2x2_ASAP7_75t_L g276 ( .A(n_207), .B(n_221), .Y(n_276) );
AND2x2_ASAP7_75t_L g347 ( .A(n_207), .B(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g368 ( .A(n_207), .Y(n_368) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_215), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx1_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g290 ( .A(n_219), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
BUFx2_ASAP7_75t_L g285 ( .A(n_220), .Y(n_285) );
AND2x2_ASAP7_75t_L g257 ( .A(n_221), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g348 ( .A(n_221), .Y(n_348) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
OR2x2_ASAP7_75t_L g294 ( .A(n_225), .B(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_SL g336 ( .A(n_225), .B(n_337), .Y(n_336) );
AOI322xp5_ASAP7_75t_L g373 ( .A1(n_225), .A2(n_252), .A3(n_374), .B1(n_376), .B2(n_379), .C1(n_381), .C2(n_383), .Y(n_373) );
AND2x2_ASAP7_75t_L g438 ( .A(n_225), .B(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_226), .B(n_252), .Y(n_262) );
AOI322xp5_ASAP7_75t_L g313 ( .A1(n_227), .A2(n_314), .A3(n_318), .B1(n_319), .B2(n_322), .C1(n_324), .C2(n_325), .Y(n_313) );
INVx2_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g365 ( .A(n_228), .B(n_318), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_228), .A2(n_425), .B1(n_427), .B2(n_430), .Y(n_424) );
OR2x2_ASAP7_75t_L g442 ( .A(n_228), .B(n_391), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_252), .B(n_253), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
AOI221xp5_ASAP7_75t_SL g292 ( .A1(n_231), .A2(n_268), .B1(n_293), .B2(n_296), .C(n_297), .Y(n_292) );
AND2x2_ASAP7_75t_L g319 ( .A(n_231), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_232), .B(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g361 ( .A(n_232), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g390 ( .A(n_233), .Y(n_390) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_250), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_234), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g332 ( .A(n_234), .Y(n_332) );
OR2x2_ASAP7_75t_L g339 ( .A(n_234), .B(n_340), .Y(n_339) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g382 ( .A(n_235), .B(n_344), .Y(n_382) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
AND2x4_ASAP7_75t_L g261 ( .A(n_236), .B(n_237), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_239), .A2(n_245), .B1(n_507), .B2(n_509), .Y(n_506) );
AND2x4_ASAP7_75t_L g239 ( .A(n_240), .B(n_243), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
NOR2x1p5_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_250), .B(n_311), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_250), .B(n_291), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_250), .Y(n_391) );
INVx1_ASAP7_75t_L g258 ( .A(n_251), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_259), .B1(n_262), .B2(n_263), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
BUFx2_ASAP7_75t_SL g369 ( .A(n_257), .Y(n_369) );
AND2x2_ASAP7_75t_L g426 ( .A(n_258), .B(n_282), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_260), .B(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_SL g298 ( .A(n_260), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_260), .B(n_419), .Y(n_418) );
BUFx3_ASAP7_75t_L g286 ( .A(n_261), .Y(n_286) );
INVx2_ASAP7_75t_L g316 ( .A(n_261), .Y(n_316) );
AND2x2_ASAP7_75t_L g359 ( .A(n_261), .B(n_343), .Y(n_359) );
INVx1_ASAP7_75t_L g273 ( .A(n_263), .Y(n_273) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI21xp5_ASAP7_75t_SL g267 ( .A1(n_268), .A2(n_273), .B(n_274), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g352 ( .A(n_271), .Y(n_352) );
INVx2_ASAP7_75t_L g340 ( .A(n_272), .Y(n_340) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x2_ASAP7_75t_L g337 ( .A(n_276), .B(n_291), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_276), .A2(n_374), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_278), .B(n_292), .Y(n_277) );
AOI32xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_281), .A3(n_283), .B1(n_287), .B2(n_290), .Y(n_278) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_279), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_279), .A2(n_368), .B1(n_386), .B2(n_388), .C(n_394), .Y(n_385) );
AND2x2_ASAP7_75t_L g405 ( .A(n_279), .B(n_286), .Y(n_405) );
BUFx2_ASAP7_75t_L g289 ( .A(n_280), .Y(n_289) );
INVx1_ASAP7_75t_L g414 ( .A(n_280), .Y(n_414) );
INVx1_ASAP7_75t_L g419 ( .A(n_280), .Y(n_419) );
INVx1_ASAP7_75t_SL g412 ( .A(n_281), .Y(n_412) );
INVx2_ASAP7_75t_L g295 ( .A(n_282), .Y(n_295) );
AND2x2_ASAP7_75t_L g407 ( .A(n_283), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g379 ( .A(n_285), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g351 ( .A(n_286), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_286), .B(n_377), .Y(n_399) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g311 ( .A(n_291), .Y(n_311) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g301 ( .A(n_295), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g310 ( .A(n_295), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g415 ( .A(n_296), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .B1(n_305), .B2(n_310), .Y(n_297) );
INVx2_ASAP7_75t_SL g389 ( .A(n_299), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_299), .B(n_428), .Y(n_430) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_301), .A2(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g346 ( .A(n_303), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g374 ( .A(n_306), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g321 ( .A(n_307), .Y(n_321) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g363 ( .A(n_309), .Y(n_363) );
INVx1_ASAP7_75t_L g408 ( .A(n_310), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_326), .C(n_349), .Y(n_312) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx2_ASAP7_75t_L g375 ( .A(n_315), .Y(n_375) );
AND2x2_ASAP7_75t_L g393 ( .A(n_315), .B(n_334), .Y(n_393) );
OR2x2_ASAP7_75t_L g432 ( .A(n_315), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_316), .B(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g328 ( .A(n_318), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g395 ( .A(n_321), .B(n_332), .Y(n_395) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_324), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g436 ( .A(n_324), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .B1(n_334), .B2(n_336), .C(n_338), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g349 ( .A1(n_327), .A2(n_350), .B(n_353), .Y(n_349) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx3_ASAP7_75t_L g380 ( .A(n_329), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_329), .B(n_423), .Y(n_422) );
INVxp33_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g341 ( .A(n_337), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B1(n_342), .B2(n_345), .Y(n_338) );
INVx2_ASAP7_75t_L g444 ( .A(n_340), .Y(n_444) );
BUFx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVxp67_ASAP7_75t_L g423 ( .A(n_348), .Y(n_423) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NOR2x1_ASAP7_75t_L g354 ( .A(n_355), .B(n_400), .Y(n_354) );
NAND4xp25_ASAP7_75t_L g355 ( .A(n_356), .B(n_373), .C(n_385), .D(n_397), .Y(n_355) );
O2A1O1Ixp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B(n_364), .C(n_366), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g396 ( .A(n_359), .Y(n_396) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g366 ( .A1(n_361), .A2(n_367), .B(n_370), .Y(n_366) );
INVx2_ASAP7_75t_L g445 ( .A(n_362), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_363), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g378 ( .A(n_363), .Y(n_378) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
OR2x2_ASAP7_75t_L g440 ( .A(n_368), .B(n_404), .Y(n_440) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_375), .Y(n_411) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND2x2_ASAP7_75t_L g381 ( .A(n_377), .B(n_382), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_377), .A2(n_407), .B(n_409), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_377), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_SL g435 ( .A(n_377), .Y(n_435) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI22xp33_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_390), .B1(n_391), .B2(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND4xp25_ASAP7_75t_L g400 ( .A(n_401), .B(n_406), .C(n_416), .D(n_437), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B1(n_413), .B2(n_415), .Y(n_409) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI211xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_420), .B(n_424), .C(n_431), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_435), .B(n_436), .Y(n_431) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
OAI21xp5_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_441), .B(n_443), .Y(n_437) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
CKINVDCx11_ASAP7_75t_R g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx2_ASAP7_75t_L g729 ( .A(n_451), .Y(n_729) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_649), .Y(n_451) );
NOR3xp33_ASAP7_75t_SL g452 ( .A(n_453), .B(n_573), .C(n_623), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_553), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_494), .B(n_534), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_484), .Y(n_456) );
INVx1_ASAP7_75t_SL g659 ( .A(n_457), .Y(n_659) );
AOI32xp33_ASAP7_75t_L g690 ( .A1(n_457), .A2(n_672), .A3(n_691), .B1(n_692), .B2(n_693), .Y(n_690) );
AND2x2_ASAP7_75t_L g692 ( .A(n_457), .B(n_549), .Y(n_692) );
AND2x4_ASAP7_75t_SL g457 ( .A(n_458), .B(n_466), .Y(n_457) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_458), .Y(n_485) );
INVx5_ASAP7_75t_L g552 ( .A(n_458), .Y(n_552) );
OR2x2_ASAP7_75t_L g559 ( .A(n_458), .B(n_551), .Y(n_559) );
INVx2_ASAP7_75t_L g564 ( .A(n_458), .Y(n_564) );
AND2x2_ASAP7_75t_L g576 ( .A(n_458), .B(n_467), .Y(n_576) );
AND2x2_ASAP7_75t_L g581 ( .A(n_458), .B(n_475), .Y(n_581) );
OR2x2_ASAP7_75t_L g588 ( .A(n_458), .B(n_487), .Y(n_588) );
AND2x4_ASAP7_75t_L g597 ( .A(n_458), .B(n_476), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_SL g639 ( .A1(n_458), .A2(n_555), .B(n_590), .C(n_628), .Y(n_639) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx3_ASAP7_75t_SL g589 ( .A(n_466), .Y(n_589) );
AND2x2_ASAP7_75t_L g635 ( .A(n_466), .B(n_552), .Y(n_635) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_475), .Y(n_466) );
AND2x2_ASAP7_75t_L g486 ( .A(n_467), .B(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g566 ( .A(n_467), .B(n_476), .Y(n_566) );
AND2x2_ASAP7_75t_L g570 ( .A(n_467), .B(n_549), .Y(n_570) );
INVx1_ASAP7_75t_L g596 ( .A(n_467), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_467), .B(n_476), .Y(n_618) );
INVx2_ASAP7_75t_L g622 ( .A(n_467), .Y(n_622) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_467), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_467), .B(n_552), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g633 ( .A(n_476), .B(n_487), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_482), .Y(n_477) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g643 ( .A(n_485), .Y(n_643) );
NAND2xp33_ASAP7_75t_SL g668 ( .A(n_485), .B(n_560), .Y(n_668) );
AND2x2_ASAP7_75t_L g710 ( .A(n_486), .B(n_552), .Y(n_710) );
AND2x2_ASAP7_75t_L g621 ( .A(n_487), .B(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g684 ( .A(n_487), .Y(n_684) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_488), .Y(n_549) );
AOI21x1_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_493), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_494), .A2(n_575), .B1(n_677), .B2(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_517), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_495), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_495), .B(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_504), .Y(n_495) );
INVx2_ASAP7_75t_L g540 ( .A(n_496), .Y(n_540) );
OR2x2_ASAP7_75t_L g544 ( .A(n_496), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_496), .B(n_557), .Y(n_562) );
AND2x4_ASAP7_75t_SL g572 ( .A(n_496), .B(n_505), .Y(n_572) );
OR2x2_ASAP7_75t_L g579 ( .A(n_496), .B(n_519), .Y(n_579) );
OR2x2_ASAP7_75t_L g591 ( .A(n_496), .B(n_505), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_496), .B(n_519), .Y(n_605) );
INVx1_ASAP7_75t_L g610 ( .A(n_496), .Y(n_610) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_496), .Y(n_628) );
AND2x2_ASAP7_75t_L g691 ( .A(n_496), .B(n_611), .Y(n_691) );
INVx2_ASAP7_75t_L g695 ( .A(n_496), .Y(n_695) );
OR2x2_ASAP7_75t_L g702 ( .A(n_496), .B(n_592), .Y(n_702) );
OR2x2_ASAP7_75t_L g724 ( .A(n_496), .B(n_725), .Y(n_724) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
AND2x2_ASAP7_75t_L g541 ( .A(n_504), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_504), .B(n_525), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_504), .B(n_601), .Y(n_663) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g560 ( .A(n_505), .Y(n_560) );
AND2x4_ASAP7_75t_L g611 ( .A(n_505), .B(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_505), .B(n_556), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_505), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_505), .B(n_545), .Y(n_704) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_511), .Y(n_505) );
AND2x2_ASAP7_75t_L g571 ( .A(n_517), .B(n_572), .Y(n_571) );
AO221x1_ASAP7_75t_L g645 ( .A1(n_517), .A2(n_560), .B1(n_591), .B2(n_646), .C(n_647), .Y(n_645) );
OAI322xp33_ASAP7_75t_L g697 ( .A1(n_517), .A2(n_617), .A3(n_698), .B1(n_700), .B2(n_701), .C1(n_702), .C2(n_703), .Y(n_697) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_525), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx3_ASAP7_75t_L g539 ( .A(n_519), .Y(n_539) );
INVx2_ASAP7_75t_L g545 ( .A(n_519), .Y(n_545) );
AND2x2_ASAP7_75t_L g557 ( .A(n_519), .B(n_525), .Y(n_557) );
INVx1_ASAP7_75t_L g602 ( .A(n_519), .Y(n_602) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_519), .Y(n_658) );
INVx1_ASAP7_75t_L g542 ( .A(n_525), .Y(n_542) );
OR2x2_ASAP7_75t_L g592 ( .A(n_525), .B(n_545), .Y(n_592) );
INVx2_ASAP7_75t_L g612 ( .A(n_525), .Y(n_612) );
INVx1_ASAP7_75t_L g665 ( .A(n_525), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_525), .B(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_532), .Y(n_527) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI21xp33_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_543), .B(n_546), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_536), .A2(n_575), .B1(n_577), .B2(n_581), .C(n_582), .Y(n_574) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_541), .Y(n_537) );
NOR2x1p5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g661 ( .A(n_540), .Y(n_661) );
INVx1_ASAP7_75t_SL g580 ( .A(n_541), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_541), .A2(n_686), .B(n_688), .Y(n_685) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_542), .Y(n_585) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_545), .Y(n_648) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
OAI211xp5_ASAP7_75t_L g623 ( .A1(n_548), .A2(n_624), .B(n_629), .C(n_640), .Y(n_623) );
OR2x2_ASAP7_75t_L g713 ( .A(n_548), .B(n_618), .Y(n_713) );
AND2x2_ASAP7_75t_L g715 ( .A(n_548), .B(n_581), .Y(n_715) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g555 ( .A(n_549), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g617 ( .A(n_549), .B(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g655 ( .A(n_549), .B(n_622), .Y(n_655) );
OA33x2_ASAP7_75t_L g662 ( .A1(n_549), .A2(n_579), .A3(n_663), .B1(n_664), .B2(n_666), .B3(n_668), .Y(n_662) );
OR2x2_ASAP7_75t_L g673 ( .A(n_549), .B(n_658), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_549), .B(n_597), .Y(n_687) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AND2x2_ASAP7_75t_L g575 ( .A(n_551), .B(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_551), .A2(n_581), .B1(n_625), .B2(n_626), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_552), .B(n_632), .C(n_665), .Y(n_664) );
AOI322xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_558), .A3(n_560), .B1(n_561), .B2(n_563), .C1(n_567), .C2(n_571), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g660 ( .A(n_556), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g615 ( .A1(n_557), .A2(n_572), .B(n_616), .C(n_619), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_558), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
NAND4xp25_ASAP7_75t_SL g679 ( .A(n_559), .B(n_588), .C(n_680), .D(n_682), .Y(n_679) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g569 ( .A(n_564), .Y(n_569) );
OR2x2_ASAP7_75t_L g614 ( .A(n_564), .B(n_566), .Y(n_614) );
AND2x2_ASAP7_75t_L g683 ( .A(n_565), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_L g688 ( .A(n_569), .B(n_683), .Y(n_688) );
BUFx2_ASAP7_75t_L g681 ( .A(n_570), .Y(n_681) );
INVx1_ASAP7_75t_SL g711 ( .A(n_571), .Y(n_711) );
AND2x4_ASAP7_75t_L g647 ( .A(n_572), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g700 ( .A(n_572), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_593), .C(n_615), .Y(n_573) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_SL g637 ( .A(n_579), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g705 ( .A1(n_579), .A2(n_706), .B(n_707), .C(n_716), .Y(n_705) );
OR2x2_ASAP7_75t_L g627 ( .A(n_580), .B(n_628), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_586), .B1(n_589), .B2(n_590), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_584), .B(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_587), .B(n_644), .Y(n_726) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g701 ( .A(n_588), .B(n_589), .Y(n_701) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g646 ( .A(n_592), .Y(n_646) );
AOI222xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_598), .B1(n_603), .B2(n_607), .C1(n_608), .C2(n_613), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_596), .Y(n_607) );
AND2x2_ASAP7_75t_L g654 ( .A(n_597), .B(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_597), .A2(n_670), .B1(n_675), .B2(n_679), .Y(n_669) );
INVx2_ASAP7_75t_SL g722 ( .A(n_597), .Y(n_722) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVxp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g678 ( .A(n_602), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_602), .B(n_665), .Y(n_725) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g638 ( .A(n_606), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_608), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g676 ( .A(n_610), .Y(n_676) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_611), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g719 ( .A(n_611), .B(n_648), .Y(n_719) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g644 ( .A(n_618), .Y(n_644) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g723 ( .A(n_621), .Y(n_723) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_622), .Y(n_667) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_634), .B(n_636), .C(n_639), .Y(n_629) );
AND2x2_ASAP7_75t_SL g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g674 ( .A(n_636), .Y(n_674) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_645), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_689), .C(n_705), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_669), .C(n_685), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B1(n_659), .B2(n_660), .C(n_662), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_671), .B(n_674), .Y(n_670) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g698 ( .A(n_684), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g706 ( .A(n_688), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_696), .Y(n_689) );
INVx2_ASAP7_75t_L g712 ( .A(n_691), .Y(n_712) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OR2x2_ASAP7_75t_L g703 ( .A(n_694), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_711), .B1(n_712), .B2(n_713), .C(n_714), .Y(n_708) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B1(n_724), .B2(n_726), .Y(n_717) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g744 ( .A(n_729), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_741), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx2_ASAP7_75t_L g753 ( .A(n_740), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_742), .B(n_745), .Y(n_741) );
CKINVDCx11_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
CKINVDCx11_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
CKINVDCx8_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
endmodule