module fake_jpeg_11519_n_589 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_589);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_589;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_58),
.B(n_101),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_59),
.Y(n_165)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_9),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_64),
.B(n_42),
.Y(n_150)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_23),
.Y(n_71)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_72),
.Y(n_168)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_78),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_20),
.B(n_9),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_111),
.Y(n_128)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_98),
.B(n_108),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_21),
.B(n_9),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_102),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_110),
.Y(n_132)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_26),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_37),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_67),
.A2(n_52),
.B1(n_24),
.B2(n_31),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_120),
.A2(n_130),
.B1(n_137),
.B2(n_148),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_70),
.A2(n_52),
.B1(n_24),
.B2(n_31),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_53),
.B(n_28),
.C(n_29),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_135),
.B(n_66),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_57),
.A2(n_52),
.B1(n_51),
.B2(n_53),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_81),
.B(n_28),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_150),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_25),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_141),
.B(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_25),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_59),
.A2(n_51),
.B1(n_36),
.B2(n_29),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_42),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_99),
.A2(n_51),
.B1(n_37),
.B2(n_36),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_159),
.B1(n_163),
.B2(n_56),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_102),
.A2(n_51),
.B1(n_50),
.B2(n_39),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_103),
.A2(n_51),
.B1(n_50),
.B2(n_39),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_79),
.B(n_34),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_164),
.B(n_109),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_69),
.A2(n_33),
.B1(n_35),
.B2(n_34),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_167),
.A2(n_130),
.B1(n_137),
.B2(n_158),
.Y(n_218)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_180),
.Y(n_266)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_181),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_183),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_185),
.A2(n_1),
.B(n_4),
.Y(n_298)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_186),
.Y(n_271)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_188),
.Y(n_264)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_189),
.Y(n_283)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_128),
.A2(n_61),
.B1(n_62),
.B2(n_68),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_191),
.A2(n_198),
.B1(n_228),
.B2(n_241),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_192),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_193),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_56),
.B1(n_66),
.B2(n_91),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_194),
.A2(n_241),
.B(n_169),
.Y(n_252)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_195),
.Y(n_269)
);

BUFx2_ASAP7_75t_SL g196 ( 
.A(n_178),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_196),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_197),
.B(n_216),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_135),
.A2(n_72),
.B1(n_97),
.B2(n_75),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_199),
.Y(n_282)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_200),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_169),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_209),
.Y(n_244)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_134),
.Y(n_202)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_202),
.Y(n_276)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_203),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_140),
.B(n_35),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_204),
.B(n_222),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_205),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_167),
.A2(n_107),
.B1(n_105),
.B2(n_90),
.Y(n_206)
);

AO22x1_ASAP7_75t_L g248 ( 
.A1(n_206),
.A2(n_143),
.B1(n_126),
.B2(n_162),
.Y(n_248)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_207),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_120),
.A2(n_83),
.B1(n_93),
.B2(n_85),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_208),
.A2(n_123),
.B1(n_171),
.B2(n_113),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_210),
.Y(n_274)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_211),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_226),
.Y(n_251)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_213),
.Y(n_291)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_214),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_156),
.A2(n_84),
.B1(n_71),
.B2(n_60),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_215),
.A2(n_118),
.B1(n_114),
.B2(n_30),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_133),
.B(n_11),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_242),
.B1(n_224),
.B2(n_205),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_219),
.Y(n_280)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_146),
.Y(n_220)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_220),
.Y(n_288)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_116),
.Y(n_221)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_145),
.B(n_0),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_146),
.Y(n_223)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_225),
.B(n_229),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_132),
.A2(n_30),
.B1(n_27),
.B2(n_11),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_227),
.A2(n_234),
.B1(n_236),
.B2(n_239),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_151),
.A2(n_30),
.B1(n_27),
.B2(n_10),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_155),
.Y(n_229)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_230),
.B(n_231),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_119),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_123),
.B(n_0),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_136),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_235),
.Y(n_245)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_154),
.B(n_10),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_172),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_238),
.Y(n_260)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_126),
.Y(n_238)
);

INVx13_ASAP7_75t_L g239 ( 
.A(n_143),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_12),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_165),
.A2(n_30),
.B1(n_27),
.B2(n_12),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_148),
.A2(n_27),
.B1(n_30),
.B2(n_2),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_182),
.B(n_163),
.C(n_159),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_243),
.B(n_273),
.C(n_206),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_198),
.A2(n_151),
.B1(n_125),
.B2(n_168),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_246),
.A2(n_265),
.B1(n_279),
.B2(n_290),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_248),
.A2(n_249),
.B1(n_253),
.B2(n_258),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_252),
.B(n_270),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_218),
.A2(n_171),
.B1(n_168),
.B2(n_125),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_242),
.A2(n_117),
.B1(n_162),
.B2(n_139),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_204),
.B(n_118),
.C(n_114),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_184),
.B(n_8),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_278),
.B(n_228),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_191),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_205),
.A2(n_8),
.B1(n_18),
.B2(n_17),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_L g290 ( 
.A1(n_206),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_222),
.A2(n_194),
.B(n_232),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_296),
.A2(n_281),
.B(n_299),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_206),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_297),
.A2(n_230),
.B1(n_234),
.B2(n_183),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_298),
.A2(n_202),
.B(n_236),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_180),
.B(n_4),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_5),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_262),
.B(n_213),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_300),
.B(n_307),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_200),
.C(n_179),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_302),
.B(n_306),
.Y(n_358)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_303),
.Y(n_362)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_259),
.Y(n_305)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_305),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_289),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_308),
.B(n_317),
.Y(n_356)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_310),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_265),
.A2(n_231),
.B1(n_223),
.B2(n_211),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_311),
.A2(n_339),
.B1(n_340),
.B2(n_346),
.Y(n_357)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_312),
.Y(n_384)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_314),
.B(n_319),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_262),
.B(n_229),
.C(n_190),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_315),
.B(n_323),
.C(n_335),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_289),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_316),
.B(n_328),
.Y(n_359)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_320),
.Y(n_355)
);

AOI32xp33_ASAP7_75t_L g321 ( 
.A1(n_296),
.A2(n_220),
.A3(n_199),
.B1(n_186),
.B2(n_221),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_321),
.A2(n_327),
.B(n_338),
.Y(n_367)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_250),
.B(n_195),
.C(n_225),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_324),
.B(n_330),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_249),
.A2(n_203),
.B1(n_217),
.B2(n_210),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_325),
.A2(n_344),
.B1(n_283),
.B2(n_264),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_247),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_289),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_252),
.B(n_187),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_329),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_272),
.B(n_226),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_272),
.B(n_238),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_331),
.B(n_334),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_332),
.A2(n_341),
.B1(n_342),
.B2(n_283),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_343),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_273),
.B(n_219),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_243),
.B(n_193),
.C(n_192),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_244),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_336),
.B(n_337),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_251),
.B(n_245),
.Y(n_337)
);

NOR3xp33_ASAP7_75t_SL g338 ( 
.A(n_278),
.B(n_239),
.C(n_14),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_286),
.Y(n_339)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_254),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_297),
.A2(n_13),
.B1(n_17),
.B2(n_7),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_279),
.A2(n_13),
.B1(n_15),
.B2(n_7),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_5),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_253),
.A2(n_8),
.B1(n_13),
.B2(n_14),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_290),
.B(n_5),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_345),
.A2(n_288),
.B(n_291),
.Y(n_371)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_248),
.A2(n_8),
.B1(n_13),
.B2(n_19),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_347),
.A2(n_295),
.B(n_263),
.Y(n_366)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_292),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_348),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_284),
.B(n_19),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_349),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_260),
.B(n_5),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_274),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_352),
.A2(n_353),
.B1(n_361),
.B2(n_379),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_313),
.A2(n_298),
.B1(n_248),
.B2(n_261),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_354),
.A2(n_360),
.B1(n_377),
.B2(n_394),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_325),
.A2(n_264),
.B1(n_287),
.B2(n_293),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_313),
.A2(n_275),
.B1(n_276),
.B2(n_254),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_327),
.A2(n_295),
.B(n_294),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_363),
.A2(n_370),
.B(n_374),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_366),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_329),
.A2(n_288),
.B(n_275),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_312),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_372),
.B(n_317),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_343),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_373),
.B(n_324),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_329),
.A2(n_268),
.B(n_291),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_309),
.A2(n_276),
.B1(n_280),
.B2(n_247),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_308),
.A2(n_280),
.B1(n_255),
.B2(n_277),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_304),
.A2(n_294),
.B(n_257),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_380),
.A2(n_301),
.B(n_326),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_334),
.B(n_266),
.C(n_269),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_382),
.B(n_387),
.C(n_350),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_335),
.A2(n_277),
.B1(n_255),
.B2(n_257),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_383),
.A2(n_385),
.B1(n_390),
.B2(n_391),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_332),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_315),
.B(n_6),
.C(n_19),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_333),
.A2(n_6),
.B1(n_331),
.B2(n_304),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_306),
.A2(n_6),
.B1(n_328),
.B2(n_316),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_301),
.A2(n_6),
.B1(n_345),
.B2(n_318),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_395),
.Y(n_438)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_365),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_396),
.B(n_398),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_393),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_356),
.B(n_323),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_406),
.C(n_412),
.Y(n_433)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_393),
.Y(n_401)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_368),
.A2(n_318),
.B1(n_341),
.B2(n_301),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_402),
.A2(n_408),
.B1(n_430),
.B2(n_391),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_403),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_404),
.B(n_417),
.Y(n_441)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_393),
.Y(n_405)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_405),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_337),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_393),
.Y(n_407)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_368),
.A2(n_342),
.B1(n_345),
.B2(n_305),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_362),
.Y(n_409)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_409),
.Y(n_451)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_410),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_307),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_411),
.B(n_418),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_356),
.B(n_336),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_375),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_413),
.B(n_425),
.Y(n_446)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_364),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_414),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_416),
.C(n_419),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_378),
.B(n_351),
.C(n_382),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_351),
.B(n_338),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_303),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_314),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_378),
.B(n_319),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_431),
.C(n_370),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_377),
.A2(n_320),
.B1(n_346),
.B2(n_322),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_422),
.A2(n_429),
.B1(n_360),
.B2(n_405),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_426),
.B(n_432),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_375),
.B(n_339),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_427),
.B(n_388),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_359),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_428),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_353),
.A2(n_348),
.B1(n_340),
.B2(n_326),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_394),
.A2(n_6),
.B1(n_310),
.B2(n_359),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_382),
.B(n_372),
.C(n_379),
.Y(n_431)
);

BUFx24_ASAP7_75t_SL g432 ( 
.A(n_358),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_434),
.B(n_460),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_420),
.A2(n_386),
.B(n_363),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_459),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_372),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_440),
.B(n_444),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_418),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_392),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_388),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_453),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_454),
.C(n_456),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_423),
.A2(n_357),
.B1(n_354),
.B2(n_358),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_452),
.A2(n_458),
.B1(n_400),
.B2(n_402),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_419),
.B(n_367),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_421),
.B(n_383),
.C(n_387),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_406),
.B(n_355),
.C(n_374),
.Y(n_456)
);

OAI21xp33_ASAP7_75t_L g457 ( 
.A1(n_428),
.A2(n_367),
.B(n_386),
.Y(n_457)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_457),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_423),
.A2(n_424),
.B1(n_429),
.B2(n_420),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_395),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_403),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_431),
.B(n_389),
.C(n_384),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_415),
.C(n_427),
.Y(n_474)
);

AO21x2_ASAP7_75t_L g466 ( 
.A1(n_401),
.A2(n_366),
.B(n_357),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_380),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_462),
.B(n_376),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_468),
.B(n_470),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_446),
.B(n_376),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_474),
.B(n_476),
.C(n_480),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_475),
.A2(n_479),
.B1(n_485),
.B2(n_490),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_435),
.B(n_407),
.C(n_411),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_477),
.B(n_456),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_452),
.A2(n_390),
.B1(n_361),
.B2(n_397),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_435),
.B(n_397),
.C(n_417),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_465),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_481),
.B(n_484),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_440),
.B(n_424),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_483),
.B(n_489),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_444),
.B(n_450),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_458),
.A2(n_408),
.B1(n_430),
.B2(n_352),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_450),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_488),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_447),
.B(n_369),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_487),
.B(n_445),
.Y(n_502)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_436),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_433),
.B(n_453),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_438),
.A2(n_385),
.B1(n_410),
.B2(n_409),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_491),
.A2(n_460),
.B(n_439),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_438),
.A2(n_414),
.B1(n_369),
.B2(n_396),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_492),
.A2(n_466),
.B1(n_439),
.B2(n_464),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_448),
.B(n_364),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_493),
.B(n_454),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_461),
.B(n_384),
.C(n_381),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_494),
.B(n_495),
.C(n_464),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_433),
.B(n_381),
.C(n_371),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_497),
.B(n_499),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_469),
.A2(n_455),
.B1(n_437),
.B2(n_442),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_498),
.A2(n_514),
.B1(n_515),
.B2(n_516),
.Y(n_535)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_500),
.Y(n_537)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_502),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_503),
.B(n_511),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_504),
.A2(n_483),
.B1(n_482),
.B2(n_495),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_443),
.C(n_441),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_507),
.B(n_518),
.Y(n_528)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_492),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_513),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_441),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_449),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_512),
.B(n_517),
.Y(n_534)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_490),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_SL g514 ( 
.A1(n_472),
.A2(n_451),
.B1(n_463),
.B2(n_466),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_472),
.A2(n_466),
.B1(n_464),
.B2(n_426),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_471),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_488),
.A2(n_466),
.B(n_365),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_475),
.A2(n_485),
.B1(n_479),
.B2(n_467),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_494),
.B(n_478),
.C(n_474),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_519),
.B(n_478),
.C(n_473),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_506),
.B(n_480),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_520),
.B(n_524),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_521),
.B(n_508),
.Y(n_543)
);

INVx11_ASAP7_75t_L g523 ( 
.A(n_502),
.Y(n_523)
);

INVx11_ASAP7_75t_L g540 ( 
.A(n_523),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_510),
.B(n_473),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_526),
.A2(n_530),
.B1(n_505),
.B2(n_500),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_503),
.B(n_482),
.C(n_477),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_527),
.B(n_531),
.C(n_538),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_496),
.A2(n_504),
.B1(n_509),
.B2(n_513),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_519),
.B(n_497),
.C(n_512),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_516),
.B(n_501),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_528),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_515),
.A2(n_517),
.B1(n_498),
.B2(n_505),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_536),
.B(n_507),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_501),
.B(n_508),
.C(n_499),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_539),
.B(n_552),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_543),
.B(n_551),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_531),
.B(n_496),
.C(n_511),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_544),
.B(n_548),
.Y(n_562)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_536),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_545),
.B(n_546),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_526),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_547),
.B(n_550),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_530),
.A2(n_537),
.B1(n_523),
.B2(n_525),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_537),
.A2(n_522),
.B(n_535),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_549),
.A2(n_540),
.B(n_545),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_533),
.Y(n_550)
);

MAJx2_ASAP7_75t_L g551 ( 
.A(n_538),
.B(n_527),
.C(n_529),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_522),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_553),
.B(n_555),
.Y(n_567)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_529),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_554),
.B(n_546),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_521),
.A2(n_530),
.B1(n_514),
.B2(n_515),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_541),
.B(n_553),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_560),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_561),
.B(n_548),
.Y(n_568)
);

INVx11_ASAP7_75t_L g564 ( 
.A(n_540),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_564),
.B(n_565),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_542),
.B(n_541),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_542),
.B(n_552),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_566),
.B(n_550),
.C(n_551),
.Y(n_570)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_568),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_570),
.B(n_573),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_562),
.A2(n_544),
.B(n_549),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_572),
.A2(n_574),
.B(n_573),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_557),
.B(n_547),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_557),
.B(n_555),
.C(n_554),
.Y(n_574)
);

INVx6_ASAP7_75t_L g575 ( 
.A(n_564),
.Y(n_575)
);

AOI31xp67_ASAP7_75t_L g576 ( 
.A1(n_575),
.A2(n_561),
.A3(n_567),
.B(n_556),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_576),
.B(n_578),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_574),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_580),
.B(n_571),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_582),
.B(n_583),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_579),
.A2(n_556),
.B(n_568),
.Y(n_583)
);

NOR3xp33_ASAP7_75t_L g585 ( 
.A(n_581),
.B(n_569),
.C(n_577),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_585),
.B(n_560),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_586),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_587),
.B(n_584),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_588),
.A2(n_563),
.B(n_559),
.Y(n_589)
);


endmodule