module fake_jpeg_29665_n_438 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_438);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_438;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_46),
.B(n_53),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_65),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_69),
.B(n_24),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_36),
.B(n_17),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_74),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_80),
.Y(n_109)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_39),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_39),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_84),
.Y(n_117)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_86),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_32),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_89),
.B(n_96),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_97),
.B(n_102),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_35),
.B1(n_26),
.B2(n_34),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_103),
.A2(n_127),
.B1(n_32),
.B2(n_22),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_64),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_47),
.B(n_24),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_55),
.A2(n_35),
.B1(n_34),
.B2(n_40),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_47),
.B(n_27),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_109),
.Y(n_151)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_48),
.B(n_59),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_95),
.B(n_129),
.Y(n_170)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_45),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_144),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_88),
.A2(n_85),
.B1(n_52),
.B2(n_79),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_164),
.B1(n_123),
.B2(n_110),
.Y(n_175)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_44),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_146),
.A2(n_147),
.B1(n_156),
.B2(n_161),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_104),
.A2(n_57),
.B1(n_42),
.B2(n_49),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_50),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_165),
.Y(n_180)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_163),
.Y(n_172)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_108),
.A2(n_23),
.B(n_19),
.C(n_41),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_162),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_104),
.A2(n_42),
.B1(n_72),
.B2(n_76),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_116),
.A2(n_42),
.B1(n_35),
.B2(n_82),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_78),
.C(n_58),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_88),
.A2(n_63),
.B1(n_75),
.B2(n_56),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_41),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_116),
.A2(n_42),
.B1(n_40),
.B2(n_22),
.Y(n_167)
);

BUFx24_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_169),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_113),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_174),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_113),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_185),
.B1(n_188),
.B2(n_170),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_140),
.A2(n_164),
.B1(n_166),
.B2(n_123),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_190),
.B1(n_94),
.B2(n_107),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_134),
.A2(n_95),
.B(n_125),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_SL g216 ( 
.A(n_188),
.B(n_130),
.C(n_111),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_110),
.B1(n_91),
.B2(n_132),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_119),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_162),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_179),
.B(n_154),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_193),
.C(n_186),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_SL g204 ( 
.A(n_198),
.B(n_157),
.C(n_152),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_204),
.B(n_208),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_165),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_151),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_212),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_155),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_194),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_133),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_180),
.B(n_27),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_215),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_111),
.B(n_193),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_198),
.B1(n_197),
.B2(n_168),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_173),
.B(n_141),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_189),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_174),
.B(n_14),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_219),
.Y(n_234)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_220),
.A2(n_222),
.B1(n_169),
.B2(n_191),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_153),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_221),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_181),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_173),
.A2(n_137),
.B1(n_160),
.B2(n_119),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_195),
.B1(n_187),
.B2(n_192),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_235),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_175),
.B1(n_198),
.B2(n_197),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_238),
.B1(n_242),
.B2(n_191),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_228),
.A2(n_199),
.B1(n_219),
.B2(n_209),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_216),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_198),
.B(n_182),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_247),
.B(n_221),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_217),
.A2(n_159),
.B1(n_94),
.B2(n_128),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_233),
.A2(n_220),
.B1(n_202),
.B2(n_169),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_132),
.B1(n_107),
.B2(n_128),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_195),
.C(n_187),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_218),
.C(n_200),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_201),
.A2(n_111),
.B(n_192),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_212),
.Y(n_248)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_230),
.B(n_243),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_249),
.B(n_224),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_138),
.Y(n_294)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_205),
.Y(n_255)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_256),
.Y(n_287)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_261),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_258),
.A2(n_239),
.B1(n_177),
.B2(n_87),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_266),
.C(n_225),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_211),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_229),
.B(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_222),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_264),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_210),
.B1(n_208),
.B2(n_200),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_263),
.A2(n_273),
.B1(n_246),
.B2(n_247),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_215),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_233),
.B1(n_231),
.B2(n_245),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_267),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_208),
.C(n_223),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_269),
.Y(n_298)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_234),
.B(n_207),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_272),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_239),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_271),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_236),
.B(n_206),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_231),
.A2(n_220),
.B1(n_202),
.B2(n_91),
.Y(n_273)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_276),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_291),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_279),
.A2(n_286),
.B1(n_302),
.B2(n_273),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_241),
.C(n_235),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_304),
.C(n_176),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_284),
.B(n_289),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_275),
.A2(n_245),
.B1(n_238),
.B2(n_229),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_225),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_235),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_224),
.Y(n_292)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

A2O1A1O1Ixp25_ASAP7_75t_L g293 ( 
.A1(n_255),
.A2(n_242),
.B(n_232),
.C(n_245),
.D(n_19),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_301),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_294),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_171),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_279),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_130),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_249),
.B(n_171),
.C(n_184),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_297),
.A2(n_275),
.B1(n_265),
.B2(n_254),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_305),
.A2(n_309),
.B1(n_320),
.B2(n_323),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_306),
.A2(n_310),
.B1(n_322),
.B2(n_298),
.Y(n_330)
);

XNOR2x1_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_250),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_308),
.B(n_293),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_297),
.A2(n_251),
.B1(n_269),
.B2(n_261),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_257),
.B1(n_256),
.B2(n_253),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_252),
.Y(n_311)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_311),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_314),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_289),
.B(n_251),
.CI(n_268),
.CON(n_314),
.SN(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_271),
.Y(n_315)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_315),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_105),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_325),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_303),
.A2(n_239),
.B1(n_87),
.B2(n_60),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_321),
.B(n_328),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_303),
.A2(n_145),
.B1(n_184),
.B2(n_176),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_280),
.B(n_105),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_277),
.C(n_284),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_278),
.A2(n_40),
.B1(n_34),
.B2(n_142),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_327),
.A2(n_287),
.B1(n_295),
.B2(n_282),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_143),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_283),
.B(n_136),
.Y(n_329)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_330),
.A2(n_331),
.B1(n_345),
.B2(n_348),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g331 ( 
.A(n_315),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_331),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_311),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_332),
.A2(n_333),
.B1(n_335),
.B2(n_307),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_329),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_341),
.C(n_342),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_322),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_339),
.A2(n_353),
.B1(n_150),
.B2(n_158),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_301),
.C(n_294),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_294),
.C(n_290),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_312),
.B(n_290),
.C(n_283),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_348),
.C(n_349),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_317),
.B(n_296),
.Y(n_344)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_344),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_347),
.A2(n_319),
.B1(n_135),
.B2(n_163),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_318),
.B(n_276),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_282),
.C(n_298),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_351),
.C(n_307),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_149),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_309),
.Y(n_352)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_352),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_305),
.A2(n_125),
.B1(n_112),
.B2(n_114),
.Y(n_353)
);

AOI322xp5_ASAP7_75t_L g356 ( 
.A1(n_337),
.A2(n_324),
.A3(n_316),
.B1(n_306),
.B2(n_314),
.C1(n_308),
.C2(n_320),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_356),
.B(n_340),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_314),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_365),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_358),
.A2(n_364),
.B1(n_366),
.B2(n_368),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_359),
.A2(n_360),
.B1(n_43),
.B2(n_1),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_121),
.Y(n_387)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_346),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_339),
.A2(n_71),
.B1(n_83),
.B2(n_67),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_373),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_351),
.A2(n_68),
.B1(n_61),
.B2(n_112),
.Y(n_368)
);

OAI322xp33_ASAP7_75t_L g369 ( 
.A1(n_334),
.A2(n_105),
.A3(n_149),
.B1(n_121),
.B2(n_15),
.C1(n_17),
.C2(n_16),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_372),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_341),
.C(n_342),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_41),
.C(n_23),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_16),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_340),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_349),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_377),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_353),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_381),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_363),
.A2(n_114),
.B1(n_34),
.B2(n_19),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_23),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_383),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_15),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_14),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_384),
.B(n_385),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_354),
.B(n_14),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_386),
.B(n_0),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_388),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_361),
.B(n_121),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_389),
.B(n_387),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_357),
.Y(n_391)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_391),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_374),
.A2(n_354),
.B(n_370),
.Y(n_393)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_393),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_395),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_371),
.C(n_368),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_397),
.B(n_400),
.C(n_401),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_359),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_399),
.B(n_22),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_366),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_371),
.Y(n_401)
);

OA21x2_ASAP7_75t_SL g403 ( 
.A1(n_390),
.A2(n_375),
.B(n_385),
.Y(n_403)
);

NAND3xp33_ASAP7_75t_SL g419 ( 
.A(n_403),
.B(n_32),
.C(n_7),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_397),
.B(n_389),
.C(n_388),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_409),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_400),
.A2(n_396),
.B1(n_391),
.B2(n_401),
.Y(n_407)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_407),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_392),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_402),
.A2(n_43),
.B1(n_22),
.B2(n_32),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_394),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_410),
.B(n_4),
.Y(n_416)
);

OAI221xp5_ASAP7_75t_L g412 ( 
.A1(n_398),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_412),
.A2(n_3),
.B(n_4),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_414),
.B(n_415),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_417),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_407),
.B(n_32),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g418 ( 
.A1(n_411),
.A2(n_5),
.B(n_6),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_410),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_6),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_413),
.A2(n_406),
.B(n_404),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_421),
.A2(n_420),
.B(n_422),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_425),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_427),
.A2(n_428),
.B(n_7),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_404),
.Y(n_428)
);

AOI322xp5_ASAP7_75t_L g429 ( 
.A1(n_426),
.A2(n_405),
.A3(n_22),
.B1(n_43),
.B2(n_10),
.C1(n_7),
.C2(n_12),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_430),
.Y(n_434)
);

AOI322xp5_ASAP7_75t_L g431 ( 
.A1(n_423),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_431),
.A2(n_8),
.B(n_9),
.Y(n_433)
);

AOI31xp67_ASAP7_75t_SL g435 ( 
.A1(n_433),
.A2(n_432),
.A3(n_9),
.B(n_10),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_435),
.B(n_434),
.C(n_8),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_436),
.A2(n_8),
.B(n_11),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_11),
.Y(n_438)
);


endmodule