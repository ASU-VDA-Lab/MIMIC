module real_jpeg_15431_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_525;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_16),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_17),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_1),
.Y(n_154)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_2),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_2),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_2),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g275 ( 
.A(n_2),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_3),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_3),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_3),
.A2(n_222),
.B1(n_380),
.B2(n_383),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g444 ( 
.A1(n_3),
.A2(n_222),
.B1(n_228),
.B2(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_3),
.A2(n_222),
.B1(n_496),
.B2(n_498),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_4),
.Y(n_117)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_4),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_5),
.A2(n_23),
.B1(n_118),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_5),
.A2(n_23),
.B1(n_173),
.B2(n_176),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_5),
.A2(n_260),
.A3(n_263),
.B1(n_264),
.B2(n_269),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_5),
.B(n_84),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_5),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_5),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_5),
.B(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_6),
.Y(n_90)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_6),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_6),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_6),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_6),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_6),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_6),
.Y(n_303)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_8),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_8),
.A2(n_50),
.B1(n_78),
.B2(n_82),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_8),
.B(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_8),
.A2(n_50),
.B1(n_296),
.B2(n_300),
.Y(n_295)
);

OAI22x1_ASAP7_75t_L g94 ( 
.A1(n_9),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_9),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_9),
.A2(n_98),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_9),
.A2(n_98),
.B1(n_242),
.B2(n_245),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_9),
.A2(n_98),
.B1(n_286),
.B2(n_289),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_12),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_12),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_12),
.Y(n_133)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_13),
.Y(n_244)
);

BUFx8_ASAP7_75t_L g502 ( 
.A(n_13),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_525),
.Y(n_17)
);

OAI221xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_65),
.B1(n_69),
.B2(n_468),
.C(n_519),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_19),
.B(n_65),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_20),
.B(n_517),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_20),
.B(n_517),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_43),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_31),
.Y(n_21)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_22),
.B(n_54),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B(n_28),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_23),
.B(n_32),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_23),
.B(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_23),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_23),
.B(n_265),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_28),
.A2(n_144),
.B1(n_227),
.B2(n_231),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_31),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_31),
.B(n_45),
.Y(n_372)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_55),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_32),
.A2(n_66),
.B1(n_68),
.B2(n_429),
.Y(n_428)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_34),
.Y(n_347)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_35),
.Y(n_230)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_38),
.Y(n_237)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_40),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_42),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g448 ( 
.A(n_42),
.Y(n_448)
);

OAI21xp33_ASAP7_75t_SL g494 ( 
.A1(n_43),
.A2(n_67),
.B(n_495),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_44),
.B(n_240),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_54),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g497 ( 
.A(n_49),
.Y(n_497)
);

O2A1O1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_50),
.A2(n_127),
.B(n_129),
.C(n_134),
.Y(n_126)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_53),
.Y(n_245)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_54),
.B(n_241),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_59),
.B1(n_62),
.B2(n_64),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_58),
.Y(n_233)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_65),
.A2(n_162),
.B1(n_350),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_65),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_65),
.A2(n_350),
.B(n_458),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_68),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_66),
.A2(n_372),
.B(n_495),
.Y(n_512)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AO221x1_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_362),
.B1(n_461),
.B2(n_466),
.C(n_467),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_254),
.B(n_361),
.Y(n_71)
);

NOR2xp67_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_211),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_73),
.B(n_211),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_141),
.C(n_167),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_74),
.B(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_110),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_75),
.B(n_111),
.C(n_140),
.Y(n_214)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_93),
.Y(n_75)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_76),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_76),
.A2(n_348),
.B(n_444),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_84),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_77),
.B(n_102),
.Y(n_253)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2x1p5_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_84),
.B(n_94),
.Y(n_252)
);

NAND2xp33_ASAP7_75t_SL g369 ( 
.A(n_84),
.B(n_344),
.Y(n_369)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_84),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_84),
.A2(n_443),
.B(n_449),
.Y(n_442)
);

AO22x2_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_103)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_93),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_102),
.Y(n_348)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_139),
.B2(n_140),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_126),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_113),
.B(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_114),
.B(n_129),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_114),
.B(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_114),
.A2(n_218),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_120),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_125),
.Y(n_187)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_125),
.Y(n_268)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_125),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_126),
.B(n_284),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_126),
.Y(n_391)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_133),
.Y(n_221)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_133),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_SL g217 ( 
.A1(n_134),
.A2(n_218),
.B(n_224),
.Y(n_217)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_137),
.Y(n_283)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_141),
.A2(n_167),
.B1(n_168),
.B2(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_141),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_162),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_142),
.A2(n_162),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_142),
.Y(n_351)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.A3(n_149),
.B1(n_155),
.B2(n_159),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_147),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_159),
.B(n_345),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_162),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_162),
.A2(n_350),
.B1(n_419),
.B2(n_420),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_162),
.B(n_420),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_165),
.B(n_166),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_163),
.A2(n_166),
.B(n_225),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_166),
.A2(n_281),
.B(n_284),
.Y(n_280)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_192),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_170),
.B(n_338),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_180),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g249 ( 
.A1(n_172),
.A2(n_181),
.B(n_193),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_172),
.B(n_193),
.Y(n_278)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_179),
.Y(n_385)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_180),
.Y(n_324)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_181),
.B(n_207),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_181),
.B(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_187),
.B1(n_188),
.B2(n_191),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_192),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_207),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_193),
.B(n_295),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_193),
.Y(n_422)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_197),
.B1(n_200),
.B2(n_204),
.Y(n_194)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_196),
.Y(n_382)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_205),
.Y(n_262)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_238),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_213),
.B(n_216),
.C(n_238),
.Y(n_407)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_226),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_217),
.B(n_226),
.Y(n_367)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_224),
.B(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_247),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_239),
.B(n_248),
.C(n_251),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_246),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_241),
.Y(n_429)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_246),
.B(n_372),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_248),
.A2(n_249),
.B1(n_477),
.B2(n_478),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_248),
.A2(n_249),
.B1(n_491),
.B2(n_492),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_249),
.B(n_477),
.C(n_479),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_249),
.B(n_492),
.C(n_493),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_252),
.B(n_341),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_253),
.Y(n_449)
);

AND2x2_ASAP7_75t_SL g492 ( 
.A(n_253),
.B(n_369),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_355),
.B(n_360),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_332),
.B(n_354),
.Y(n_255)
);

AOI21x1_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_307),
.B(n_331),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_279),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_258),
.B(n_279),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_276),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_259),
.B(n_276),
.Y(n_329)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

NAND2xp67_ASAP7_75t_L g389 ( 
.A(n_278),
.B(n_294),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_292),
.Y(n_279)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_280),
.Y(n_353)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_285),
.Y(n_320)
);

INVx4_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_292)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_294),
.A2(n_421),
.B(n_422),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_304),
.B(n_305),
.C(n_353),
.Y(n_352)
);

OAI21x1_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_326),
.B(n_330),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_321),
.B(n_325),
.Y(n_308)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_319),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_315),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_323),
.Y(n_325)
);

NAND2xp33_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_379),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_329),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_352),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_352),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_349),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_339),
.B2(n_340),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_340),
.C(n_349),
.Y(n_359)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_338),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2x1_ASAP7_75t_L g426 ( 
.A(n_342),
.B(n_427),
.Y(n_426)
);

NOR2x1_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_348),
.Y(n_342)
);

AOI21x1_ASAP7_75t_L g394 ( 
.A1(n_343),
.A2(n_348),
.B(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_359),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_356),
.B(n_359),
.Y(n_360)
);

NOR3xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_410),
.C(n_432),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_406),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_364),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_398),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_365),
.B(n_398),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_374),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_375),
.C(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.C(n_370),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_368),
.A2(n_370),
.B1(n_371),
.B2(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_368),
.Y(n_402)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_387),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_376),
.A2(n_378),
.B(n_386),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_386),
.Y(n_377)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

XNOR2x1_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_392),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_388),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_389),
.B(n_390),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_393),
.A2(n_394),
.B1(n_396),
.B2(n_397),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_394),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_394),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_511)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_394),
.Y(n_514)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_396),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_415),
.C(n_416),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_403),
.C(n_405),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_409),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_405),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_407),
.B(n_408),
.Y(n_464)
);

A2O1A1Ixp33_ASAP7_75t_L g461 ( 
.A1(n_410),
.A2(n_462),
.B(n_463),
.C(n_465),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_411),
.B(n_413),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_417),
.Y(n_413)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_414),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_423),
.B1(n_430),
.B2(n_431),
.Y(n_417)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_434),
.C(n_435),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_423),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_424),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_426),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_428),
.B(n_438),
.C(n_439),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_431),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_432),
.Y(n_466)
);

NOR2x1_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_436),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_436),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_440),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_437),
.B(n_441),
.C(n_484),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_453),
.B1(n_459),
.B2(n_460),
.Y(n_440)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_441),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_450),
.B(n_452),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_451),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx3_ASAP7_75t_SL g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_452),
.A2(n_473),
.B1(n_474),
.B2(n_481),
.Y(n_472)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_452),
.Y(n_481)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_453),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_455),
.B1(n_457),
.B2(n_458),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_457),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_460),
.Y(n_484)
);

NAND3xp33_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_507),
.C(n_516),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_485),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_483),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_471),
.B(n_483),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_482),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_474),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_475),
.A2(n_476),
.B1(n_479),
.B2(n_480),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_477),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_479),
.A2(n_480),
.B1(n_489),
.B2(n_504),
.Y(n_488)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_489),
.C(n_509),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_482),
.C(n_506),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_485),
.A2(n_521),
.B(n_522),
.Y(n_520)
);

NOR2x1_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_505),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_486),
.B(n_505),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_487),
.Y(n_509)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_489),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_490),
.A2(n_493),
.B1(n_494),
.B2(n_503),
.Y(n_489)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_490),
.Y(n_503)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVxp33_ASAP7_75t_SL g493 ( 
.A(n_494),
.Y(n_493)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g519 ( 
.A1(n_507),
.A2(n_516),
.B(n_520),
.C(n_523),
.D(n_524),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_508),
.B(n_510),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_510),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_515),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_512),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_512),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_514),
.B(n_515),
.C(n_518),
.Y(n_517)
);


endmodule