module fake_ibex_719_n_5648 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_974, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_854, n_1008, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_993, n_1012, n_689, n_960, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_1004, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_5648);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_974;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_689;
input n_960;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_1004;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_5648;

wire n_4557;
wire n_5285;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_4204;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3472;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_4801;
wire n_3639;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_1070;
wire n_4510;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_3565;
wire n_5304;
wire n_3883;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_4854;
wire n_3769;
wire n_1445;
wire n_2147;
wire n_5591;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_5261;
wire n_1078;
wire n_4422;
wire n_1865;
wire n_5033;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_1118;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_2550;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_5612;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_4290;
wire n_1549;
wire n_1531;
wire n_2919;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_1121;
wire n_4823;
wire n_5195;
wire n_5541;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_5609;
wire n_4757;
wire n_5254;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_3950;
wire n_1042;
wire n_5252;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_5238;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_1932;
wire n_3775;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_4374;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3529;
wire n_3222;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_5199;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_5099;
wire n_1210;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_2361;
wire n_4128;
wire n_5213;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_5163;
wire n_1408;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_2046;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_4674;
wire n_1232;
wire n_2715;
wire n_4679;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_3796;
wire n_5157;
wire n_1836;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_5216;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_1448;
wire n_3034;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_5083;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_1967;
wire n_1095;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_3428;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_3339;
wire n_3673;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_3269;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_1025;
wire n_2679;
wire n_4028;
wire n_1517;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_1763;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1021;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_4729;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_3099;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_1017;
wire n_2049;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_5566;
wire n_5342;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_4417;
wire n_1550;
wire n_1169;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_2194;
wire n_1072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_5332;
wire n_3096;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_5227;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_5472;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_5546;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_4919;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_1047;
wire n_1878;
wire n_4803;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_2871;
wire n_2764;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_5403;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_1459;
wire n_4032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_1303;
wire n_1994;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4789;
wire n_4778;
wire n_2703;
wire n_2574;
wire n_5492;
wire n_1887;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_5260;
wire n_5069;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_5309;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_3742;
wire n_3532;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_4686;
wire n_4682;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_5186;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_5180;
wire n_4733;
wire n_5368;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_1166;
wire n_5267;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_4962;
wire n_5397;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_4644;
wire n_4412;
wire n_4266;
wire n_5605;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_5384;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_1230;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_5107;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_2961;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1033;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_5506;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_5253;
wire n_3789;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_5390;
wire n_4926;
wire n_5043;
wire n_5097;
wire n_4688;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_3904;
wire n_4378;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_3726;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4970;
wire n_4652;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5551;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5319;
wire n_5543;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_5621;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_3030;
wire n_5631;
wire n_4503;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_3210;
wire n_3221;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5221;
wire n_1301;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_4610;
wire n_4067;
wire n_4997;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_5357;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5619;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_1312;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_5294;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_5089;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_1711;
wire n_3069;
wire n_5465;
wire n_3107;
wire n_5488;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_1053;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_3757;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5514;
wire n_2554;
wire n_1676;
wire n_1013;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_1014;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_3394;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_3488;
wire n_2832;
wire n_4991;
wire n_1028;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_3703;
wire n_5116;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_5194;
wire n_4579;
wire n_5628;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_2398;
wire n_1593;
wire n_1775;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_3074;
wire n_4640;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_5193;
wire n_2170;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_5153;
wire n_5369;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_2463;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_3350;
wire n_5399;
wire n_4873;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_4636;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_4609;
wire n_5148;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_1067;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_1331;
wire n_1223;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_1294;
wire n_1351;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_3336;
wire n_1291;
wire n_3763;
wire n_4284;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_1662;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_1962;
wire n_5296;
wire n_5159;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_2309;
wire n_2274;
wire n_5096;
wire n_3712;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_4643;
wire n_5217;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_2214;
wire n_1066;
wire n_1726;
wire n_1241;
wire n_2589;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_1238;
wire n_3959;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_3044;
wire n_2868;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_4905;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_5277;
wire n_3647;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_5569;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1018;
wire n_1669;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_1175;
wire n_4408;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_5645;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_1507;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_5114;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_5395;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_1798;
wire n_5559;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_5295;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_5047;
wire n_5504;
wire n_5076;
wire n_3543;
wire n_3655;
wire n_3791;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_3898;
wire n_3366;
wire n_1024;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_4961;
wire n_5013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_3207;
wire n_5450;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_3036;
wire n_5012;
wire n_5376;
wire n_4207;
wire n_1022;
wire n_1760;
wire n_5208;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_5503;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_5644;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_5324;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5022;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_5245;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_5329;
wire n_5510;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_1780;
wire n_1091;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_5061;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_5132;
wire n_4883;
wire n_1079;
wire n_3559;
wire n_5184;
wire n_4943;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_3838;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_5618;
wire n_4159;
wire n_4372;
wire n_5528;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_5464;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_1829;
wire n_1338;
wire n_1327;
wire n_5204;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_2565;
wire n_4201;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_3996;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_1841;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_3802;
wire n_5343;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_3765;
wire n_2216;
wire n_4259;
wire n_1620;
wire n_5196;
wire n_5086;
wire n_3518;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_2899;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_2564;
wire n_5110;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_1764;
wire n_1019;
wire n_1250;
wire n_1190;
wire n_4598;
wire n_3259;
wire n_5483;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_1803;
wire n_5264;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_4604;
wire n_5123;
wire n_3467;
wire n_4240;
wire n_2219;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_2539;
wire n_1701;
wire n_5236;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4126;
wire n_4103;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_2748;
wire n_5359;
wire n_2224;
wire n_5526;
wire n_2233;
wire n_2499;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_5147;
wire n_5407;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_5389;
wire n_3171;
wire n_1733;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_1189;
wire n_4995;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_4205;
wire n_3790;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_5435;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_2063;
wire n_1076;
wire n_3082;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_1712;
wire n_4537;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_3248;
wire n_2606;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_5084;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_4876;
wire n_5322;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_1264;
wire n_2808;
wire n_5010;
wire n_3396;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_3599;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_4587;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_1115;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_2419;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_5170;
wire n_1523;
wire n_1086;
wire n_1756;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_4496;
wire n_1528;
wire n_3840;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_1413;
wire n_2464;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_1706;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_2414;
wire n_5642;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_2684;
wire n_2205;
wire n_1104;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_5136;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_1920;
wire n_4306;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_5634;
wire n_3028;
wire n_3228;
wire n_5079;
wire n_3706;
wire n_1432;
wire n_3322;
wire n_1174;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_2694;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_5606;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_2180;
wire n_3376;
wire n_2617;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_4832;
wire n_5229;
wire n_3666;
wire n_1839;
wire n_5160;
wire n_1587;
wire n_2555;
wire n_2330;
wire n_5313;
wire n_2108;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_2196;
wire n_1538;
wire n_3773;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_1889;
wire n_1124;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_1054;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_1642;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_2587;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_3410;
wire n_4900;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_2299;
wire n_2078;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_2315;
wire n_3623;
wire n_5558;
wire n_2157;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5223;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_4334;
wire n_2211;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_1501;
wire n_5636;
wire n_5106;
wire n_5257;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_2893;
wire n_2009;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_5623;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_5178;
wire n_1105;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_5592;
wire n_5484;
wire n_4982;
wire n_5418;
wire n_5432;
wire n_1769;
wire n_1060;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_5156;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_5139;
wire n_4555;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_3989;
wire n_5565;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_3191;
wire n_1029;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_5500;
wire n_5293;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_1336;
wire n_1358;
wire n_3318;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_1074;
wire n_5059;
wire n_1462;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_1692;
wire n_4796;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_5038;
wire n_3837;
wire n_4841;
wire n_3076;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_1027;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_2331;
wire n_1600;
wire n_4701;
wire n_5248;
wire n_4088;
wire n_2136;
wire n_5443;
wire n_1913;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_5533;
wire n_1822;
wire n_1804;
wire n_1581;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_4329;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_4327;
wire n_5412;
wire n_2656;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_1016;
wire n_4465;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_4224;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_2368;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_1080;
wire n_5377;
wire n_2290;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_4912;
wire n_1971;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_2571;
wire n_5479;
wire n_5598;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_5211;
wire n_1668;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_4311;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_3881;
wire n_1030;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_5279;
wire n_4650;
wire n_1038;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_5613;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_5063;
wire n_4671;
wire n_1326;
wire n_4981;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_2723;
wire n_4054;
wire n_1569;
wire n_4012;
wire n_5582;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_3560;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_5467;
wire n_2646;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_4755;
wire n_3827;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_2416;
wire n_2962;
wire n_1031;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_1036;
wire n_5331;
wire n_1106;
wire n_4655;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_5456;
wire n_5523;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_5512;
wire n_3436;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_4527;
wire n_2877;
wire n_1996;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5077;
wire n_5214;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_3624;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_3145;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_1464;
wire n_1566;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_2252;
wire n_1982;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2991;
wire n_2699;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_4042;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_4764;
wire n_4899;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_1357;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_5604;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_2117;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_3638;
wire n_2106;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_5105;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_4133;
wire n_3985;
wire n_5481;
wire n_5187;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_3747;
wire n_1323;
wire n_3710;
wire n_1429;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_5200;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_2271;
wire n_2356;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_2642;
wire n_5485;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_5355;
wire n_4048;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_5185;
wire n_2849;
wire n_5091;
wire n_1177;
wire n_3292;
wire n_3940;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_3047;
wire n_2610;
wire n_5306;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_4383;
wire n_2709;
wire n_5074;
wire n_2244;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5409;
wire n_2581;
wire n_5540;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_2137;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_4222;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_1167;
wire n_3231;
wire n_3138;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_1788;
wire n_2348;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_5082;
wire n_1907;
wire n_3994;
wire n_5118;
wire n_2135;
wire n_1088;
wire n_1102;
wire n_5145;
wire n_4487;
wire n_1165;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_2869;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_2667;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_1542;
wire n_1547;
wire n_1362;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_1951;
wire n_1330;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_4761;
wire n_2021;
wire n_2713;
wire n_3227;
wire n_2938;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_2061;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_2827;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_2491;
wire n_5298;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_4147;
wire n_3992;
wire n_4811;
wire n_5093;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_2296;
wire n_1911;
wire n_2870;
wire n_4869;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_5283;
wire n_1419;
wire n_4738;
wire n_1193;
wire n_2928;
wire n_3380;
wire n_3557;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_1499;
wire n_2155;
wire n_3938;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_3053;
wire n_1039;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1026;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_1791;
wire n_5301;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_5507;
wire n_1164;
wire n_3749;
wire n_5470;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_4280;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_5393;
wire n_4978;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_1417;
wire n_5455;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_1410;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_717),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_273),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_630),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_180),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_806),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_525),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_964),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_69),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_48),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_1005),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_425),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_133),
.Y(n_1024)
);

CKINVDCx16_ASAP7_75t_R g1025 ( 
.A(n_718),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_907),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_593),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_497),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_282),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_851),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_873),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_709),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_607),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_19),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_785),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_190),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_991),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_258),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_138),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_284),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_371),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_933),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_878),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_757),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_449),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_802),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_165),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_877),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_167),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_32),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_554),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_31),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_543),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_138),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_201),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_36),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_169),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_896),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_783),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_982),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_513),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_76),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_490),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_651),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_992),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_909),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_116),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_633),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_840),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_962),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_730),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_820),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_942),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_781),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_446),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_881),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_476),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_798),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_506),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_716),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_590),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_679),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_193),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_296),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_961),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_729),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_887),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_870),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_21),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_780),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_993),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_772),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_196),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_353),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_89),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_501),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_458),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_957),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_443),
.Y(n_1099)
);

CKINVDCx16_ASAP7_75t_R g1100 ( 
.A(n_776),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_929),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_293),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_840),
.Y(n_1103)
);

BUFx10_ASAP7_75t_L g1104 ( 
.A(n_928),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_934),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_869),
.Y(n_1106)
);

BUFx5_ASAP7_75t_L g1107 ( 
.A(n_142),
.Y(n_1107)
);

CKINVDCx16_ASAP7_75t_R g1108 ( 
.A(n_614),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_870),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_568),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_174),
.Y(n_1111)
);

BUFx10_ASAP7_75t_L g1112 ( 
.A(n_735),
.Y(n_1112)
);

BUFx8_ASAP7_75t_SL g1113 ( 
.A(n_703),
.Y(n_1113)
);

CKINVDCx14_ASAP7_75t_R g1114 ( 
.A(n_493),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_469),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_774),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_473),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_553),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_959),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_692),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_901),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_756),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_711),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_385),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_276),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_121),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_876),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_613),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_431),
.Y(n_1129)
);

CKINVDCx20_ASAP7_75t_R g1130 ( 
.A(n_868),
.Y(n_1130)
);

BUFx10_ASAP7_75t_L g1131 ( 
.A(n_441),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_857),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_434),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_326),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_67),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_335),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_180),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_533),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_37),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_217),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_114),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_730),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_227),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_852),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_329),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_363),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_778),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_3),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_141),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_560),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_867),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_452),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_922),
.Y(n_1153)
);

BUFx5_ASAP7_75t_L g1154 ( 
.A(n_998),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_247),
.Y(n_1155)
);

CKINVDCx16_ASAP7_75t_R g1156 ( 
.A(n_240),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_602),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_29),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_291),
.Y(n_1159)
);

CKINVDCx14_ASAP7_75t_R g1160 ( 
.A(n_613),
.Y(n_1160)
);

CKINVDCx16_ASAP7_75t_R g1161 ( 
.A(n_74),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_570),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_121),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_345),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_295),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_479),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_985),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_219),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_641),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_274),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_875),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_580),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_151),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_764),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_993),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_514),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_668),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_126),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_804),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1007),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_297),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_970),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_792),
.Y(n_1183)
);

CKINVDCx16_ASAP7_75t_R g1184 ( 
.A(n_249),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_72),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_991),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_592),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_20),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_115),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_60),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_624),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_917),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_467),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_79),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_122),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_254),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_144),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_584),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_167),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_4),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_880),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_559),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1011),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_921),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_127),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_383),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_938),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_843),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_463),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_621),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_524),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_545),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_168),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_905),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_974),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_75),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_89),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_522),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_925),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_608),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_914),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_851),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_94),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_970),
.Y(n_1224)
);

BUFx10_ASAP7_75t_L g1225 ( 
.A(n_168),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_100),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_521),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_3),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_249),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_277),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1007),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_893),
.Y(n_1232)
);

BUFx10_ASAP7_75t_L g1233 ( 
.A(n_27),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_400),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_188),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_421),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_302),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_830),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_546),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_969),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_49),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_72),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_571),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_684),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_667),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_676),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_254),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_569),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_285),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_454),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_923),
.Y(n_1251)
);

CKINVDCx16_ASAP7_75t_R g1252 ( 
.A(n_337),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_770),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_255),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_866),
.Y(n_1255)
);

BUFx8_ASAP7_75t_SL g1256 ( 
.A(n_272),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_281),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_237),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_360),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_588),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_662),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_576),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_172),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_131),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_14),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_95),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_691),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_973),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_969),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_362),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_788),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_729),
.Y(n_1272)
);

BUFx10_ASAP7_75t_L g1273 ( 
.A(n_904),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_986),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_348),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_950),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_974),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_996),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_562),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_871),
.Y(n_1280)
);

BUFx10_ASAP7_75t_L g1281 ( 
.A(n_982),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_877),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_659),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_277),
.Y(n_1284)
);

BUFx10_ASAP7_75t_L g1285 ( 
.A(n_393),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_959),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_416),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_997),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_723),
.Y(n_1289)
);

BUFx10_ASAP7_75t_L g1290 ( 
.A(n_733),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_916),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_828),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_900),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_397),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_177),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_891),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_674),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_921),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_919),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_848),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_777),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_630),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1008),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_995),
.Y(n_1304)
);

CKINVDCx16_ASAP7_75t_R g1305 ( 
.A(n_519),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_576),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_507),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_709),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_174),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_427),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1005),
.Y(n_1311)
);

CKINVDCx16_ASAP7_75t_R g1312 ( 
.A(n_487),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_715),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_183),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_395),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_958),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_911),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_750),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_275),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1009),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_977),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_979),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_946),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_968),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_308),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_327),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_491),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1006),
.Y(n_1328)
);

BUFx10_ASAP7_75t_L g1329 ( 
.A(n_937),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_515),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_696),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_265),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_908),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_932),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_625),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_209),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_116),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_294),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_935),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_221),
.Y(n_1340)
);

BUFx10_ASAP7_75t_L g1341 ( 
.A(n_390),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_388),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_30),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_975),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_158),
.Y(n_1345)
);

BUFx10_ASAP7_75t_L g1346 ( 
.A(n_214),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_898),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_459),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_930),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_586),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_965),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_931),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_673),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_357),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_349),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_260),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_918),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_939),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_366),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_536),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_894),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_994),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_593),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_237),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_42),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_903),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_828),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_772),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_569),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_279),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_563),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_622),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_952),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_109),
.Y(n_1374)
);

BUFx8_ASAP7_75t_SL g1375 ( 
.A(n_32),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_100),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_200),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_160),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_763),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_936),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_479),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_661),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_80),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_889),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_332),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_724),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_268),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_591),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_858),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_282),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_372),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_69),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_947),
.Y(n_1393)
);

BUFx5_ASAP7_75t_L g1394 ( 
.A(n_926),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_245),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_41),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_234),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_433),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_281),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_496),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_613),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_973),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_812),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_891),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_508),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_494),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_888),
.Y(n_1407)
);

BUFx2_ASAP7_75t_SL g1408 ( 
.A(n_936),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_595),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_35),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_886),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_163),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_372),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_949),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_714),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_749),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_890),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_5),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_415),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_948),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_964),
.Y(n_1421)
);

BUFx8_ASAP7_75t_SL g1422 ( 
.A(n_915),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_546),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_245),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_981),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_788),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_81),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_875),
.Y(n_1428)
);

BUFx2_ASAP7_75t_SL g1429 ( 
.A(n_897),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_616),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_52),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_631),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_147),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_879),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_76),
.Y(n_1435)
);

BUFx8_ASAP7_75t_SL g1436 ( 
.A(n_219),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_800),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_462),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_999),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_744),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_533),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_879),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_151),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_454),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_987),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_872),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_444),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_600),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_461),
.Y(n_1449)
);

BUFx10_ASAP7_75t_L g1450 ( 
.A(n_798),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_421),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_125),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_63),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_954),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_126),
.Y(n_1455)
);

BUFx5_ASAP7_75t_L g1456 ( 
.A(n_980),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_966),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_920),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_531),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_899),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_943),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_405),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_647),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_820),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_977),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_885),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_505),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_848),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_171),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_19),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_236),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_517),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_944),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_949),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_308),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_46),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_164),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_114),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_436),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_47),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_554),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_473),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1012),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_907),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_967),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_154),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_31),
.Y(n_1487)
);

BUFx5_ASAP7_75t_L g1488 ( 
.A(n_323),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_984),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_482),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_941),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_147),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_924),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_316),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_412),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_523),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_16),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_989),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_883),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_564),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_214),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_326),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_592),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_955),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_507),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_292),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_874),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_67),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_243),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_320),
.Y(n_1510)
);

CKINVDCx16_ASAP7_75t_R g1511 ( 
.A(n_990),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_895),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_301),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_825),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_773),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_600),
.Y(n_1516)
);

CKINVDCx16_ASAP7_75t_R g1517 ( 
.A(n_1003),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_135),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_648),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1009),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_963),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_534),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_41),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_566),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_56),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_836),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_884),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_899),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1000),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1010),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_763),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_474),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_686),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_902),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_839),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1004),
.Y(n_1536)
);

CKINVDCx16_ASAP7_75t_R g1537 ( 
.A(n_199),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_619),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_61),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_972),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_683),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_423),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_88),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_849),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_889),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_823),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1008),
.Y(n_1547)
);

CKINVDCx14_ASAP7_75t_R g1548 ( 
.A(n_429),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_961),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1001),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_912),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_99),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_146),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_892),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_902),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_179),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_634),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_422),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_315),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_927),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_593),
.Y(n_1561)
);

BUFx10_ASAP7_75t_L g1562 ( 
.A(n_906),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_189),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_910),
.Y(n_1564)
);

BUFx10_ASAP7_75t_L g1565 ( 
.A(n_15),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_766),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_956),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_951),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_647),
.Y(n_1569)
);

CKINVDCx16_ASAP7_75t_R g1570 ( 
.A(n_793),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_190),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_781),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_913),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_737),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_625),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_901),
.Y(n_1576)
);

BUFx10_ASAP7_75t_L g1577 ( 
.A(n_419),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_269),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_289),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_180),
.Y(n_1580)
);

CKINVDCx20_ASAP7_75t_R g1581 ( 
.A(n_927),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_832),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_960),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_540),
.Y(n_1584)
);

BUFx10_ASAP7_75t_L g1585 ( 
.A(n_983),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_648),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_222),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_7),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_500),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_953),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_945),
.Y(n_1591)
);

CKINVDCx16_ASAP7_75t_R g1592 ( 
.A(n_971),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_742),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_306),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_356),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_203),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_741),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_24),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_978),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_836),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_854),
.Y(n_1601)
);

BUFx10_ASAP7_75t_L g1602 ( 
.A(n_976),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_604),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_988),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_882),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1002),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_371),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_606),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1006),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_703),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_57),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_940),
.Y(n_1612)
);

BUFx5_ASAP7_75t_L g1613 ( 
.A(n_426),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1052),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1113),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1113),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1049),
.B(n_1),
.Y(n_1617)
);

INVxp33_ASAP7_75t_SL g1618 ( 
.A(n_1036),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1094),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1114),
.Y(n_1620)
);

CKINVDCx14_ASAP7_75t_R g1621 ( 
.A(n_1114),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1149),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1229),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1295),
.Y(n_1624)
);

INVxp33_ASAP7_75t_L g1625 ( 
.A(n_1050),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1160),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1160),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1195),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1348),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1376),
.Y(n_1630)
);

CKINVDCx14_ASAP7_75t_R g1631 ( 
.A(n_1548),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1533),
.Y(n_1632)
);

INVxp67_ASAP7_75t_SL g1633 ( 
.A(n_1021),
.Y(n_1633)
);

INVxp67_ASAP7_75t_SL g1634 ( 
.A(n_1021),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1256),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1022),
.B(n_0),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1548),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1220),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1226),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1283),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1451),
.Y(n_1641)
);

INVxp67_ASAP7_75t_SL g1642 ( 
.A(n_1034),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1496),
.Y(n_1643)
);

INVxp67_ASAP7_75t_SL g1644 ( 
.A(n_1034),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1103),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1016),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1256),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1375),
.Y(n_1648)
);

INVxp33_ASAP7_75t_L g1649 ( 
.A(n_1059),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1089),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1028),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1033),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1038),
.Y(n_1653)
);

INVxp67_ASAP7_75t_SL g1654 ( 
.A(n_1089),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1362),
.Y(n_1655)
);

INVxp33_ASAP7_75t_L g1656 ( 
.A(n_1612),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1055),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1118),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1067),
.Y(n_1659)
);

INVxp33_ASAP7_75t_SL g1660 ( 
.A(n_1013),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1082),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1118),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1093),
.Y(n_1663)
);

CKINVDCx16_ASAP7_75t_R g1664 ( 
.A(n_1025),
.Y(n_1664)
);

INVxp67_ASAP7_75t_L g1665 ( 
.A(n_1202),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1108),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1202),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1111),
.Y(n_1668)
);

CKINVDCx16_ASAP7_75t_R g1669 ( 
.A(n_1156),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1120),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1126),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1129),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1436),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1145),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1148),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1155),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1158),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1275),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1334),
.Y(n_1679)
);

INVxp33_ASAP7_75t_L g1680 ( 
.A(n_1436),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1164),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1176),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1181),
.Y(n_1683)
);

CKINVDCx20_ASAP7_75t_R g1684 ( 
.A(n_1040),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1422),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1190),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1191),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1422),
.Y(n_1688)
);

CKINVDCx16_ASAP7_75t_R g1689 ( 
.A(n_1161),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1275),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1194),
.Y(n_1691)
);

CKINVDCx14_ASAP7_75t_R g1692 ( 
.A(n_1131),
.Y(n_1692)
);

CKINVDCx16_ASAP7_75t_R g1693 ( 
.A(n_1184),
.Y(n_1693)
);

CKINVDCx20_ASAP7_75t_R g1694 ( 
.A(n_1045),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1205),
.Y(n_1695)
);

INVxp67_ASAP7_75t_SL g1696 ( 
.A(n_1310),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1252),
.Y(n_1697)
);

CKINVDCx16_ASAP7_75t_R g1698 ( 
.A(n_1305),
.Y(n_1698)
);

CKINVDCx16_ASAP7_75t_R g1699 ( 
.A(n_1312),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1334),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1210),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1211),
.Y(n_1702)
);

INVxp33_ASAP7_75t_L g1703 ( 
.A(n_1035),
.Y(n_1703)
);

INVxp67_ASAP7_75t_SL g1704 ( 
.A(n_1310),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1154),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1537),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1361),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1241),
.Y(n_1708)
);

INVxp67_ASAP7_75t_SL g1709 ( 
.A(n_1378),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1245),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1378),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1080),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1258),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1261),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1014),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1116),
.Y(n_1716)
);

CKINVDCx14_ASAP7_75t_R g1717 ( 
.A(n_1131),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1262),
.Y(n_1718)
);

CKINVDCx16_ASAP7_75t_R g1719 ( 
.A(n_1131),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1264),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1279),
.Y(n_1721)
);

CKINVDCx16_ASAP7_75t_R g1722 ( 
.A(n_1341),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1287),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1302),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1308),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1154),
.Y(n_1726)
);

INVxp67_ASAP7_75t_SL g1727 ( 
.A(n_1444),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1325),
.Y(n_1728)
);

INVxp67_ASAP7_75t_SL g1729 ( 
.A(n_1444),
.Y(n_1729)
);

CKINVDCx20_ASAP7_75t_R g1730 ( 
.A(n_1083),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1335),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_1015),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1343),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1154),
.Y(n_1734)
);

CKINVDCx20_ASAP7_75t_R g1735 ( 
.A(n_1110),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1355),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1359),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1360),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1364),
.Y(n_1739)
);

INVxp33_ASAP7_75t_SL g1740 ( 
.A(n_1023),
.Y(n_1740)
);

INVxp33_ASAP7_75t_SL g1741 ( 
.A(n_1024),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1369),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1341),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1371),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1388),
.Y(n_1745)
);

CKINVDCx20_ASAP7_75t_R g1746 ( 
.A(n_1115),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1154),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1027),
.Y(n_1748)
);

CKINVDCx20_ASAP7_75t_R g1749 ( 
.A(n_1166),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1390),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1029),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1395),
.Y(n_1752)
);

CKINVDCx14_ASAP7_75t_R g1753 ( 
.A(n_1346),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1398),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1399),
.Y(n_1755)
);

BUFx12f_ASAP7_75t_L g1756 ( 
.A(n_1647),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1625),
.B(n_1346),
.Y(n_1757)
);

OAI22x1_ASAP7_75t_L g1758 ( 
.A1(n_1666),
.A2(n_1032),
.B1(n_1053),
.B2(n_1047),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1679),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1658),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1626),
.B(n_1037),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1743),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1716),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1627),
.B(n_1373),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1618),
.A2(n_1054),
.B1(n_1057),
.B2(n_1056),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1692),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1700),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1717),
.B(n_1346),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1753),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1743),
.B(n_1061),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1719),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1662),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1707),
.Y(n_1773)
);

BUFx12f_ASAP7_75t_L g1774 ( 
.A(n_1648),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1706),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1614),
.B(n_1520),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1662),
.Y(n_1777)
);

INVx2_ASAP7_75t_SL g1778 ( 
.A(n_1722),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1665),
.B(n_1062),
.Y(n_1779)
);

OAI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1726),
.A2(n_1235),
.B(n_1051),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1665),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1621),
.A2(n_1064),
.B1(n_1068),
.B2(n_1063),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1667),
.B(n_1075),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1716),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1628),
.A2(n_1081),
.B1(n_1095),
.B2(n_1077),
.Y(n_1785)
);

OAI22x1_ASAP7_75t_L g1786 ( 
.A1(n_1673),
.A2(n_1097),
.B1(n_1099),
.B2(n_1096),
.Y(n_1786)
);

CKINVDCx8_ASAP7_75t_R g1787 ( 
.A(n_1664),
.Y(n_1787)
);

INVx6_ASAP7_75t_L g1788 ( 
.A(n_1669),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1619),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1638),
.B(n_1440),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1734),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1667),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1649),
.B(n_1225),
.Y(n_1793)
);

CKINVDCx8_ASAP7_75t_R g1794 ( 
.A(n_1689),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1631),
.A2(n_1102),
.B1(n_1124),
.B2(n_1123),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1622),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1660),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1645),
.A2(n_1125),
.B1(n_1133),
.B2(n_1128),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1747),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1711),
.B(n_1134),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1711),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1623),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1716),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1624),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1629),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1633),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1634),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1715),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1630),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1740),
.Y(n_1810)
);

BUFx6f_ASAP7_75t_L g1811 ( 
.A(n_1632),
.Y(n_1811)
);

INVx6_ASAP7_75t_L g1812 ( 
.A(n_1693),
.Y(n_1812)
);

AND2x2_ASAP7_75t_SL g1813 ( 
.A(n_1698),
.B(n_1100),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1642),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1655),
.B(n_1504),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1646),
.Y(n_1816)
);

OA21x2_ASAP7_75t_L g1817 ( 
.A1(n_1651),
.A2(n_1653),
.B(n_1652),
.Y(n_1817)
);

OA21x2_ASAP7_75t_L g1818 ( 
.A1(n_1755),
.A2(n_1659),
.B(n_1657),
.Y(n_1818)
);

INVx4_ASAP7_75t_L g1819 ( 
.A(n_1620),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1644),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1712),
.A2(n_1135),
.B1(n_1137),
.B2(n_1136),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1650),
.B(n_1138),
.Y(n_1822)
);

OA21x2_ASAP7_75t_L g1823 ( 
.A1(n_1661),
.A2(n_1239),
.B(n_1236),
.Y(n_1823)
);

OAI22x1_ASAP7_75t_L g1824 ( 
.A1(n_1685),
.A2(n_1140),
.B1(n_1141),
.B2(n_1139),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1699),
.A2(n_1146),
.B1(n_1152),
.B2(n_1143),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1663),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1654),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1656),
.A2(n_1157),
.B1(n_1162),
.B2(n_1159),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_SL g1829 ( 
.A1(n_1684),
.A2(n_1169),
.B1(n_1223),
.B2(n_1168),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1678),
.B(n_1163),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1741),
.B(n_1554),
.Y(n_1831)
);

INVx4_ASAP7_75t_L g1832 ( 
.A(n_1637),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1690),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1668),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1639),
.A2(n_1165),
.B1(n_1172),
.B2(n_1170),
.Y(n_1835)
);

INVx6_ASAP7_75t_L g1836 ( 
.A(n_1617),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1640),
.B(n_1225),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1696),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1670),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1704),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1709),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1671),
.Y(n_1842)
);

INVx3_ASAP7_75t_L g1843 ( 
.A(n_1672),
.Y(n_1843)
);

INVx5_ASAP7_75t_L g1844 ( 
.A(n_1727),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1729),
.B(n_1173),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1641),
.B(n_1643),
.Y(n_1846)
);

OAI22x1_ASAP7_75t_R g1847 ( 
.A1(n_1694),
.A2(n_1263),
.B1(n_1284),
.B2(n_1244),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1674),
.Y(n_1848)
);

BUFx2_ASAP7_75t_L g1849 ( 
.A(n_1732),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1748),
.B(n_1560),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1675),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1676),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1677),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1681),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1682),
.Y(n_1855)
);

BUFx6f_ASAP7_75t_L g1856 ( 
.A(n_1683),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1751),
.B(n_1574),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1686),
.Y(n_1858)
);

INVx4_ASAP7_75t_L g1859 ( 
.A(n_1697),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1687),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1691),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1695),
.B(n_1177),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1701),
.Y(n_1863)
);

AOI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1636),
.A2(n_1185),
.B1(n_1187),
.B2(n_1178),
.Y(n_1864)
);

OA21x2_ASAP7_75t_L g1865 ( 
.A1(n_1702),
.A2(n_1239),
.B(n_1236),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1708),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1710),
.Y(n_1867)
);

OA21x2_ASAP7_75t_L g1868 ( 
.A1(n_1754),
.A2(n_1248),
.B(n_1247),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1713),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1714),
.Y(n_1870)
);

INVx2_ASAP7_75t_SL g1871 ( 
.A(n_1718),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1720),
.Y(n_1872)
);

NAND2xp33_ASAP7_75t_L g1873 ( 
.A(n_1721),
.B(n_1107),
.Y(n_1873)
);

OA21x2_ASAP7_75t_L g1874 ( 
.A1(n_1752),
.A2(n_1248),
.B(n_1247),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1723),
.Y(n_1875)
);

CKINVDCx20_ASAP7_75t_R g1876 ( 
.A(n_1730),
.Y(n_1876)
);

BUFx6f_ASAP7_75t_L g1877 ( 
.A(n_1724),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1725),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1728),
.Y(n_1879)
);

BUFx8_ASAP7_75t_L g1880 ( 
.A(n_1616),
.Y(n_1880)
);

INVx6_ASAP7_75t_L g1881 ( 
.A(n_1703),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1731),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1733),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1736),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1737),
.Y(n_1885)
);

BUFx6f_ASAP7_75t_L g1886 ( 
.A(n_1738),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1739),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1742),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1744),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1745),
.Y(n_1890)
);

OAI21x1_ASAP7_75t_L g1891 ( 
.A1(n_1750),
.A2(n_1306),
.B(n_1249),
.Y(n_1891)
);

BUFx6f_ASAP7_75t_L g1892 ( 
.A(n_1688),
.Y(n_1892)
);

INVxp67_ASAP7_75t_L g1893 ( 
.A(n_1680),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1735),
.B(n_1361),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1746),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1635),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1749),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1679),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1743),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1658),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1679),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1679),
.Y(n_1902)
);

INVx3_ASAP7_75t_L g1903 ( 
.A(n_1743),
.Y(n_1903)
);

BUFx3_ASAP7_75t_L g1904 ( 
.A(n_1743),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1658),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1658),
.Y(n_1906)
);

BUFx3_ASAP7_75t_L g1907 ( 
.A(n_1743),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1679),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1626),
.B(n_1499),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1658),
.Y(n_1910)
);

BUFx6f_ASAP7_75t_L g1911 ( 
.A(n_1716),
.Y(n_1911)
);

BUFx12f_ASAP7_75t_L g1912 ( 
.A(n_1647),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1692),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1692),
.Y(n_1914)
);

OAI21x1_ASAP7_75t_L g1915 ( 
.A1(n_1705),
.A2(n_1306),
.B(n_1249),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1679),
.Y(n_1916)
);

AND2x6_ASAP7_75t_L g1917 ( 
.A(n_1743),
.B(n_1452),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1716),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1716),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1658),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_SL g1921 ( 
.A1(n_1684),
.A2(n_1309),
.B1(n_1319),
.B2(n_1294),
.Y(n_1921)
);

BUFx6f_ASAP7_75t_L g1922 ( 
.A(n_1716),
.Y(n_1922)
);

OA21x2_ASAP7_75t_L g1923 ( 
.A1(n_1705),
.A2(n_1381),
.B(n_1370),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1626),
.B(n_1188),
.Y(n_1924)
);

AND2x2_ASAP7_75t_SL g1925 ( 
.A(n_1719),
.B(n_1511),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1658),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1679),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1743),
.B(n_1517),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1692),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1743),
.Y(n_1930)
);

INVx2_ASAP7_75t_SL g1931 ( 
.A(n_1743),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1743),
.Y(n_1932)
);

BUFx6f_ASAP7_75t_L g1933 ( 
.A(n_1716),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1658),
.Y(n_1934)
);

OA21x2_ASAP7_75t_L g1935 ( 
.A1(n_1705),
.A2(n_1381),
.B(n_1370),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1743),
.B(n_1570),
.Y(n_1936)
);

INVx2_ASAP7_75t_SL g1937 ( 
.A(n_1743),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1658),
.Y(n_1938)
);

BUFx6f_ASAP7_75t_L g1939 ( 
.A(n_1716),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1692),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_1692),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1658),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1679),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1625),
.B(n_1233),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1626),
.B(n_1551),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1626),
.B(n_1551),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1679),
.Y(n_1947)
);

OA21x2_ASAP7_75t_L g1948 ( 
.A1(n_1705),
.A2(n_1387),
.B(n_1382),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1658),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1716),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1679),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1626),
.B(n_1193),
.Y(n_1952)
);

INVx5_ASAP7_75t_L g1953 ( 
.A(n_1743),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1658),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1658),
.Y(n_1955)
);

BUFx6f_ASAP7_75t_L g1956 ( 
.A(n_1716),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_L g1957 ( 
.A1(n_1705),
.A2(n_1387),
.B(n_1382),
.Y(n_1957)
);

CKINVDCx8_ASAP7_75t_R g1958 ( 
.A(n_1719),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1626),
.B(n_1196),
.Y(n_1959)
);

BUFx8_ASAP7_75t_SL g1960 ( 
.A(n_1615),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1658),
.Y(n_1961)
);

INVx4_ASAP7_75t_L g1962 ( 
.A(n_1719),
.Y(n_1962)
);

OA21x2_ASAP7_75t_L g1963 ( 
.A1(n_1705),
.A2(n_1508),
.B(n_1463),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1743),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1658),
.Y(n_1965)
);

INVx4_ASAP7_75t_L g1966 ( 
.A(n_1719),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1679),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_1716),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1716),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1626),
.B(n_1197),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1658),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1679),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1679),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1679),
.Y(n_1974)
);

BUFx2_ASAP7_75t_L g1975 ( 
.A(n_1692),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1881),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1960),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1914),
.Y(n_1978)
);

CKINVDCx20_ASAP7_75t_R g1979 ( 
.A(n_1876),
.Y(n_1979)
);

NOR2xp67_ASAP7_75t_L g1980 ( 
.A(n_1966),
.B(n_0),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1802),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_1929),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1940),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1804),
.Y(n_1984)
);

BUFx10_ASAP7_75t_L g1985 ( 
.A(n_1913),
.Y(n_1985)
);

INVx3_ASAP7_75t_L g1986 ( 
.A(n_1809),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1789),
.Y(n_1987)
);

INVx3_ASAP7_75t_L g1988 ( 
.A(n_1809),
.Y(n_1988)
);

CKINVDCx20_ASAP7_75t_R g1989 ( 
.A(n_1958),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1941),
.Y(n_1990)
);

CKINVDCx20_ASAP7_75t_R g1991 ( 
.A(n_1958),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1771),
.Y(n_1992)
);

CKINVDCx20_ASAP7_75t_R g1993 ( 
.A(n_1797),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1891),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1823),
.Y(n_1995)
);

CKINVDCx20_ASAP7_75t_R g1996 ( 
.A(n_1810),
.Y(n_1996)
);

CKINVDCx20_ASAP7_75t_R g1997 ( 
.A(n_1769),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1775),
.B(n_1592),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_R g1999 ( 
.A(n_1787),
.B(n_1327),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1975),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_1756),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1774),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1912),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1865),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1880),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1796),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1871),
.B(n_1150),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1805),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1868),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1816),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1903),
.B(n_1270),
.Y(n_2011)
);

BUFx10_ASAP7_75t_L g2012 ( 
.A(n_1778),
.Y(n_2012)
);

BUFx2_ASAP7_75t_L g2013 ( 
.A(n_1944),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1874),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1794),
.Y(n_2015)
);

CKINVDCx16_ASAP7_75t_R g2016 ( 
.A(n_1847),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1780),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1794),
.Y(n_2018)
);

INVxp67_ASAP7_75t_SL g2019 ( 
.A(n_1944),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_1757),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_R g2021 ( 
.A(n_1778),
.B(n_1338),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1915),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1843),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1849),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1957),
.Y(n_2025)
);

CKINVDCx16_ASAP7_75t_R g2026 ( 
.A(n_1768),
.Y(n_2026)
);

BUFx2_ASAP7_75t_L g2027 ( 
.A(n_1836),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1788),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_1793),
.Y(n_2029)
);

OAI22xp33_ASAP7_75t_SL g2030 ( 
.A1(n_1765),
.A2(n_1199),
.B1(n_1200),
.B2(n_1198),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1812),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1895),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1829),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1921),
.Y(n_2034)
);

CKINVDCx20_ASAP7_75t_R g2035 ( 
.A(n_1808),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_1925),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1923),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1813),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1825),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1859),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1892),
.Y(n_2041)
);

AO21x2_ASAP7_75t_L g2042 ( 
.A1(n_1873),
.A2(n_1415),
.B(n_1401),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1892),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1837),
.B(n_1233),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1828),
.Y(n_2045)
);

CKINVDCx20_ASAP7_75t_R g2046 ( 
.A(n_1821),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1896),
.Y(n_2047)
);

NOR2xp67_ASAP7_75t_L g2048 ( 
.A(n_1893),
.B(n_1),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1878),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1782),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1935),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_R g2052 ( 
.A(n_1897),
.B(n_1410),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1795),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1835),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1758),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1811),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_1837),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1785),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_1798),
.Y(n_2059)
);

CKINVDCx20_ASAP7_75t_R g2060 ( 
.A(n_1864),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1948),
.Y(n_2061)
);

CKINVDCx20_ASAP7_75t_R g2062 ( 
.A(n_1819),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1832),
.Y(n_2063)
);

CKINVDCx20_ASAP7_75t_R g2064 ( 
.A(n_1844),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1786),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1786),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1963),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1852),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1852),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1856),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_1824),
.Y(n_2071)
);

NOR2xp67_ASAP7_75t_L g2072 ( 
.A(n_1953),
.B(n_1),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1894),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1856),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_1846),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1860),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_1844),
.Y(n_2077)
);

INVx2_ASAP7_75t_SL g2078 ( 
.A(n_1953),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_1817),
.Y(n_2079)
);

CKINVDCx20_ASAP7_75t_R g2080 ( 
.A(n_1924),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1850),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1869),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_1857),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1877),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_R g2085 ( 
.A(n_1917),
.B(n_1438),
.Y(n_2085)
);

CKINVDCx5p33_ASAP7_75t_R g2086 ( 
.A(n_1762),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_1899),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1871),
.B(n_1372),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_1904),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1877),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1886),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1886),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_R g2093 ( 
.A(n_1917),
.B(n_1455),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_1907),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1779),
.B(n_1107),
.Y(n_2095)
);

INVx3_ASAP7_75t_L g2096 ( 
.A(n_1818),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1806),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1759),
.Y(n_2098)
);

CKINVDCx5p33_ASAP7_75t_R g2099 ( 
.A(n_1932),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1767),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_1831),
.Y(n_2101)
);

CKINVDCx20_ASAP7_75t_R g2102 ( 
.A(n_1952),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1807),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1928),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_1936),
.Y(n_2105)
);

NOR2xp67_ASAP7_75t_L g2106 ( 
.A(n_1930),
.B(n_2),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_1783),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_R g2108 ( 
.A(n_1917),
.B(n_1462),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1814),
.Y(n_2109)
);

CKINVDCx5p33_ASAP7_75t_R g2110 ( 
.A(n_1800),
.Y(n_2110)
);

CKINVDCx16_ASAP7_75t_R g2111 ( 
.A(n_1909),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_R g2112 ( 
.A(n_1964),
.B(n_1476),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1820),
.Y(n_2113)
);

HB1xp67_ASAP7_75t_L g2114 ( 
.A(n_1959),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_1770),
.B(n_1463),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_1970),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1773),
.Y(n_2117)
);

CKINVDCx20_ASAP7_75t_R g2118 ( 
.A(n_1822),
.Y(n_2118)
);

CKINVDCx5p33_ASAP7_75t_R g2119 ( 
.A(n_1790),
.Y(n_2119)
);

AOI21x1_ASAP7_75t_L g2120 ( 
.A1(n_1791),
.A2(n_1419),
.B(n_1418),
.Y(n_2120)
);

CKINVDCx5p33_ASAP7_75t_R g2121 ( 
.A(n_1815),
.Y(n_2121)
);

BUFx3_ASAP7_75t_L g2122 ( 
.A(n_1898),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1827),
.Y(n_2123)
);

CKINVDCx5p33_ASAP7_75t_R g2124 ( 
.A(n_1830),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1845),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_1931),
.B(n_1206),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_1764),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1833),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1838),
.Y(n_2129)
);

BUFx6f_ASAP7_75t_L g2130 ( 
.A(n_1901),
.Y(n_2130)
);

INVx1_ASAP7_75t_SL g2131 ( 
.A(n_1862),
.Y(n_2131)
);

CKINVDCx5p33_ASAP7_75t_R g2132 ( 
.A(n_1761),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1840),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_1841),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1826),
.Y(n_2135)
);

CKINVDCx20_ASAP7_75t_R g2136 ( 
.A(n_1760),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1834),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1902),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_1945),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_1946),
.Y(n_2140)
);

CKINVDCx5p33_ASAP7_75t_R g2141 ( 
.A(n_1937),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_1937),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1772),
.Y(n_2143)
);

NOR2xp33_ASAP7_75t_R g2144 ( 
.A(n_1777),
.B(n_1505),
.Y(n_2144)
);

CKINVDCx20_ASAP7_75t_R g2145 ( 
.A(n_1781),
.Y(n_2145)
);

OAI21x1_ASAP7_75t_L g2146 ( 
.A1(n_1851),
.A2(n_1518),
.B(n_1508),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_R g2147 ( 
.A(n_1792),
.B(n_1506),
.Y(n_2147)
);

NOR2x1p5_ASAP7_75t_L g2148 ( 
.A(n_1801),
.B(n_1209),
.Y(n_2148)
);

CKINVDCx20_ASAP7_75t_R g2149 ( 
.A(n_1900),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_1905),
.Y(n_2150)
);

NOR2xp33_ASAP7_75t_R g2151 ( 
.A(n_1906),
.B(n_1541),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1908),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_1910),
.Y(n_2153)
);

CKINVDCx20_ASAP7_75t_R g2154 ( 
.A(n_1920),
.Y(n_2154)
);

CKINVDCx5p33_ASAP7_75t_R g2155 ( 
.A(n_1926),
.Y(n_2155)
);

CKINVDCx16_ASAP7_75t_R g2156 ( 
.A(n_1934),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_R g2157 ( 
.A(n_1938),
.B(n_1543),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_1942),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1916),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_1949),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1839),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_1954),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_1955),
.B(n_1212),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_1961),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1842),
.Y(n_2165)
);

CKINVDCx5p33_ASAP7_75t_R g2166 ( 
.A(n_1965),
.Y(n_2166)
);

CKINVDCx5p33_ASAP7_75t_R g2167 ( 
.A(n_1971),
.Y(n_2167)
);

CKINVDCx20_ASAP7_75t_R g2168 ( 
.A(n_1853),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_R g2169 ( 
.A(n_1776),
.B(n_1579),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_1927),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1861),
.B(n_1107),
.Y(n_2171)
);

HB1xp67_ASAP7_75t_L g2172 ( 
.A(n_1848),
.Y(n_2172)
);

CKINVDCx16_ASAP7_75t_R g2173 ( 
.A(n_1863),
.Y(n_2173)
);

OAI22xp33_ASAP7_75t_SL g2174 ( 
.A1(n_1866),
.A2(n_1216),
.B1(n_1217),
.B2(n_1213),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_1943),
.Y(n_2175)
);

CKINVDCx5p33_ASAP7_75t_R g2176 ( 
.A(n_1947),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_R g2177 ( 
.A(n_1870),
.B(n_1580),
.Y(n_2177)
);

NOR2xp33_ASAP7_75t_R g2178 ( 
.A(n_1875),
.B(n_1584),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_1951),
.Y(n_2179)
);

NOR2xp67_ASAP7_75t_L g2180 ( 
.A(n_1967),
.B(n_2),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_1972),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1854),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1973),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_1855),
.B(n_1020),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1858),
.Y(n_2185)
);

BUFx6f_ASAP7_75t_L g2186 ( 
.A(n_1974),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_1867),
.B(n_1218),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1872),
.Y(n_2188)
);

CKINVDCx20_ASAP7_75t_R g2189 ( 
.A(n_1879),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1882),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1883),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_1884),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_1885),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1887),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1888),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_R g2196 ( 
.A(n_1889),
.B(n_1058),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_1890),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_1799),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_R g2199 ( 
.A(n_1763),
.B(n_1091),
.Y(n_2199)
);

CKINVDCx16_ASAP7_75t_R g2200 ( 
.A(n_1763),
.Y(n_2200)
);

CKINVDCx20_ASAP7_75t_R g2201 ( 
.A(n_1784),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_1784),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_1803),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_1803),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1911),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1911),
.Y(n_2206)
);

BUFx3_ASAP7_75t_L g2207 ( 
.A(n_1918),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_1918),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1919),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1919),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1922),
.Y(n_2211)
);

BUFx2_ASAP7_75t_L g2212 ( 
.A(n_1922),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1933),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_1933),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_1939),
.Y(n_2215)
);

CKINVDCx20_ASAP7_75t_R g2216 ( 
.A(n_1939),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1950),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_1956),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_1956),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_1968),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1968),
.Y(n_2221)
);

INVx3_ASAP7_75t_L g2222 ( 
.A(n_1969),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_1809),
.Y(n_2223)
);

HB1xp67_ASAP7_75t_L g2224 ( 
.A(n_1881),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_1881),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1802),
.Y(n_2226)
);

CKINVDCx5p33_ASAP7_75t_R g2227 ( 
.A(n_1881),
.Y(n_2227)
);

NOR2xp33_ASAP7_75t_R g2228 ( 
.A(n_1766),
.B(n_1119),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1802),
.Y(n_2229)
);

BUFx6f_ASAP7_75t_L g2230 ( 
.A(n_1891),
.Y(n_2230)
);

CKINVDCx5p33_ASAP7_75t_R g2231 ( 
.A(n_1881),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1802),
.Y(n_2232)
);

CKINVDCx5p33_ASAP7_75t_R g2233 ( 
.A(n_1881),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_R g2234 ( 
.A(n_1766),
.B(n_1130),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_1881),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_1881),
.Y(n_2236)
);

CKINVDCx20_ASAP7_75t_R g2237 ( 
.A(n_1876),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_1881),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_1881),
.Y(n_2239)
);

XNOR2x2_ASAP7_75t_L g2240 ( 
.A(n_1758),
.B(n_1041),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_R g2241 ( 
.A(n_1766),
.B(n_1174),
.Y(n_2241)
);

INVx2_ASAP7_75t_SL g2242 ( 
.A(n_1881),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_1881),
.Y(n_2243)
);

HB1xp67_ASAP7_75t_L g2244 ( 
.A(n_1881),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_1881),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_1881),
.Y(n_2246)
);

CKINVDCx16_ASAP7_75t_R g2247 ( 
.A(n_1962),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1881),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_1881),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_1881),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_1881),
.Y(n_2251)
);

AOI21x1_ASAP7_75t_L g2252 ( 
.A1(n_1891),
.A2(n_1430),
.B(n_1424),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_1881),
.Y(n_2253)
);

AOI21x1_ASAP7_75t_L g2254 ( 
.A1(n_1891),
.A2(n_1433),
.B(n_1432),
.Y(n_2254)
);

CKINVDCx5p33_ASAP7_75t_R g2255 ( 
.A(n_1881),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_2146),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1995),
.Y(n_2257)
);

BUFx2_ASAP7_75t_L g2258 ( 
.A(n_2177),
.Y(n_2258)
);

INVx3_ASAP7_75t_L g2259 ( 
.A(n_1985),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2172),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2131),
.B(n_1227),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2097),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2124),
.B(n_1228),
.Y(n_2263)
);

AND2x4_ASAP7_75t_L g2264 ( 
.A(n_2062),
.B(n_1222),
.Y(n_2264)
);

BUFx2_ASAP7_75t_L g2265 ( 
.A(n_2178),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2103),
.Y(n_2266)
);

AND2x6_ASAP7_75t_L g2267 ( 
.A(n_2044),
.B(n_1578),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_2125),
.B(n_1230),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2004),
.Y(n_2269)
);

NOR2x1p5_ASAP7_75t_L g2270 ( 
.A(n_2005),
.B(n_1234),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2109),
.Y(n_2271)
);

AND2x4_ASAP7_75t_L g2272 ( 
.A(n_2242),
.B(n_1224),
.Y(n_2272)
);

OR2x2_ASAP7_75t_L g2273 ( 
.A(n_2173),
.B(n_1079),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2009),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_2057),
.B(n_1237),
.Y(n_2275)
);

AOI22xp33_ASAP7_75t_L g2276 ( 
.A1(n_2019),
.A2(n_1578),
.B1(n_1589),
.B2(n_1583),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2014),
.Y(n_2277)
);

BUFx2_ASAP7_75t_L g2278 ( 
.A(n_2021),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_2225),
.B(n_1317),
.Y(n_2279)
);

INVx3_ASAP7_75t_L g2280 ( 
.A(n_1985),
.Y(n_2280)
);

INVx4_ASAP7_75t_L g2281 ( 
.A(n_2227),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2014),
.Y(n_2282)
);

INVx4_ASAP7_75t_L g2283 ( 
.A(n_2231),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_2107),
.B(n_1242),
.Y(n_2284)
);

AND2x6_ASAP7_75t_L g2285 ( 
.A(n_2113),
.B(n_1589),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2184),
.B(n_1243),
.Y(n_2286)
);

INVx5_ASAP7_75t_L g2287 ( 
.A(n_2247),
.Y(n_2287)
);

INVx4_ASAP7_75t_L g2288 ( 
.A(n_2233),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2014),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2252),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_2012),
.Y(n_2291)
);

BUFx3_ASAP7_75t_L g2292 ( 
.A(n_2201),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2110),
.B(n_1246),
.Y(n_2293)
);

OR2x6_ASAP7_75t_L g2294 ( 
.A(n_2224),
.B(n_1408),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2254),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2123),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_R g2297 ( 
.A(n_2028),
.B(n_1366),
.Y(n_2297)
);

AND2x6_ASAP7_75t_L g2298 ( 
.A(n_2128),
.B(n_1018),
.Y(n_2298)
);

BUFx3_ASAP7_75t_L g2299 ( 
.A(n_2216),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2129),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_2012),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1994),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2134),
.A2(n_2118),
.B1(n_2045),
.B2(n_2168),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_L g2304 ( 
.A(n_2029),
.B(n_1250),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2133),
.Y(n_2305)
);

AND2x6_ASAP7_75t_L g2306 ( 
.A(n_2010),
.B(n_1018),
.Y(n_2306)
);

BUFx6f_ASAP7_75t_L g2307 ( 
.A(n_1994),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1981),
.Y(n_2308)
);

BUFx6f_ASAP7_75t_L g2309 ( 
.A(n_1994),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2114),
.B(n_1254),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2230),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2230),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2013),
.B(n_1285),
.Y(n_2313)
);

BUFx3_ASAP7_75t_L g2314 ( 
.A(n_2064),
.Y(n_2314)
);

BUFx2_ASAP7_75t_L g2315 ( 
.A(n_2196),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1984),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2230),
.Y(n_2317)
);

AND2x2_ASAP7_75t_SL g2318 ( 
.A(n_2016),
.B(n_2026),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2226),
.Y(n_2319)
);

BUFx2_ASAP7_75t_L g2320 ( 
.A(n_2235),
.Y(n_2320)
);

INVx2_ASAP7_75t_SL g2321 ( 
.A(n_2244),
.Y(n_2321)
);

INVx3_ASAP7_75t_L g2322 ( 
.A(n_2200),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2229),
.Y(n_2323)
);

OAI22xp5_ASAP7_75t_L g2324 ( 
.A1(n_2188),
.A2(n_1403),
.B1(n_1411),
.B2(n_1384),
.Y(n_2324)
);

INVx3_ASAP7_75t_L g2325 ( 
.A(n_2236),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2116),
.B(n_1257),
.Y(n_2326)
);

OR2x2_ASAP7_75t_L g2327 ( 
.A(n_1998),
.B(n_1084),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_L g2328 ( 
.A(n_2104),
.B(n_1259),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_2192),
.B(n_1260),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2020),
.B(n_1285),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2232),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2024),
.B(n_1565),
.Y(n_2332)
);

OR2x2_ASAP7_75t_L g2333 ( 
.A(n_2156),
.B(n_1189),
.Y(n_2333)
);

INVx3_ASAP7_75t_L g2334 ( 
.A(n_2238),
.Y(n_2334)
);

INVx1_ASAP7_75t_SL g2335 ( 
.A(n_2189),
.Y(n_2335)
);

OR2x6_ASAP7_75t_L g2336 ( 
.A(n_2027),
.B(n_1429),
.Y(n_2336)
);

AND2x4_ASAP7_75t_L g2337 ( 
.A(n_2239),
.B(n_1493),
.Y(n_2337)
);

INVx2_ASAP7_75t_SL g2338 ( 
.A(n_2243),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_2193),
.B(n_1265),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_2195),
.B(n_2197),
.Y(n_2340)
);

INVx1_ASAP7_75t_SL g2341 ( 
.A(n_2245),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_2040),
.B(n_1266),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2144),
.B(n_1577),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_2105),
.B(n_1267),
.Y(n_2344)
);

BUFx3_ASAP7_75t_L g2345 ( 
.A(n_2246),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2120),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_L g2347 ( 
.A(n_2127),
.B(n_1289),
.Y(n_2347)
);

BUFx6f_ASAP7_75t_L g2348 ( 
.A(n_2063),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2007),
.B(n_1297),
.Y(n_2349)
);

INVx5_ASAP7_75t_L g2350 ( 
.A(n_2111),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_2198),
.B(n_1307),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_SL g2352 ( 
.A(n_2088),
.B(n_1313),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_2119),
.B(n_2121),
.Y(n_2353)
);

NAND2xp33_ASAP7_75t_R g2354 ( 
.A(n_1999),
.B(n_1314),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_2130),
.Y(n_2355)
);

NAND3x1_ASAP7_75t_L g2356 ( 
.A(n_1977),
.B(n_1581),
.C(n_1529),
.Y(n_2356)
);

AND2x4_ASAP7_75t_L g2357 ( 
.A(n_2248),
.B(n_1590),
.Y(n_2357)
);

NOR2xp33_ASAP7_75t_L g2358 ( 
.A(n_2132),
.B(n_2101),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_2143),
.B(n_1315),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_2130),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2147),
.B(n_1273),
.Y(n_2361)
);

AND2x6_ASAP7_75t_L g2362 ( 
.A(n_2023),
.B(n_1018),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2037),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2135),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2137),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2151),
.B(n_1273),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2187),
.B(n_1326),
.Y(n_2367)
);

OR2x2_ASAP7_75t_SL g2368 ( 
.A(n_1993),
.B(n_1591),
.Y(n_2368)
);

AOI22xp33_ASAP7_75t_L g2369 ( 
.A1(n_2163),
.A2(n_1488),
.B1(n_1613),
.B2(n_1107),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2161),
.B(n_1330),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2165),
.Y(n_2371)
);

INVx3_ASAP7_75t_L g2372 ( 
.A(n_2249),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2182),
.Y(n_2373)
);

AND2x6_ASAP7_75t_L g2374 ( 
.A(n_2049),
.B(n_1018),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2051),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2250),
.B(n_2251),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2185),
.Y(n_2377)
);

BUFx6f_ASAP7_75t_L g2378 ( 
.A(n_2130),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_SL g2379 ( 
.A(n_2150),
.B(n_2153),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2061),
.Y(n_2380)
);

BUFx3_ASAP7_75t_L g2381 ( 
.A(n_2253),
.Y(n_2381)
);

AOI22xp33_ASAP7_75t_L g2382 ( 
.A1(n_2148),
.A2(n_2030),
.B1(n_2174),
.B2(n_2190),
.Y(n_2382)
);

BUFx2_ASAP7_75t_L g2383 ( 
.A(n_2255),
.Y(n_2383)
);

BUFx6f_ASAP7_75t_L g2384 ( 
.A(n_2186),
.Y(n_2384)
);

NOR2x1p5_ASAP7_75t_L g2385 ( 
.A(n_2001),
.B(n_1331),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2191),
.Y(n_2386)
);

BUFx3_ASAP7_75t_L g2387 ( 
.A(n_1997),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2194),
.Y(n_2388)
);

BUFx6f_ASAP7_75t_L g2389 ( 
.A(n_2186),
.Y(n_2389)
);

INVxp67_ASAP7_75t_SL g2390 ( 
.A(n_2035),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2171),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1987),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2006),
.Y(n_2393)
);

INVx3_ASAP7_75t_L g2394 ( 
.A(n_2122),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2008),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2067),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2106),
.Y(n_2397)
);

AND2x4_ASAP7_75t_L g2398 ( 
.A(n_2031),
.B(n_1604),
.Y(n_2398)
);

BUFx6f_ASAP7_75t_L g2399 ( 
.A(n_2186),
.Y(n_2399)
);

AND3x1_ASAP7_75t_L g2400 ( 
.A(n_1989),
.B(n_1991),
.C(n_1979),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_2155),
.B(n_1332),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2157),
.B(n_1273),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2126),
.B(n_1336),
.Y(n_2403)
);

CKINVDCx20_ASAP7_75t_R g2404 ( 
.A(n_1996),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2079),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2011),
.B(n_1337),
.Y(n_2406)
);

BUFx6f_ASAP7_75t_L g2407 ( 
.A(n_2202),
.Y(n_2407)
);

CKINVDCx20_ASAP7_75t_R g2408 ( 
.A(n_2237),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2158),
.B(n_1340),
.Y(n_2409)
);

HB1xp67_ASAP7_75t_L g2410 ( 
.A(n_2075),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2079),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2169),
.B(n_1450),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2098),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2100),
.Y(n_2414)
);

INVx4_ASAP7_75t_L g2415 ( 
.A(n_2000),
.Y(n_2415)
);

AND2x2_ASAP7_75t_SL g2416 ( 
.A(n_2085),
.B(n_1518),
.Y(n_2416)
);

INVxp33_ASAP7_75t_L g2417 ( 
.A(n_2112),
.Y(n_2417)
);

INVx4_ASAP7_75t_L g2418 ( 
.A(n_2077),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2096),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2117),
.Y(n_2420)
);

INVx4_ASAP7_75t_L g2421 ( 
.A(n_2002),
.Y(n_2421)
);

INVx4_ASAP7_75t_L g2422 ( 
.A(n_2003),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2081),
.B(n_1342),
.Y(n_2423)
);

AOI22xp33_ASAP7_75t_L g2424 ( 
.A1(n_2115),
.A2(n_1107),
.B1(n_1613),
.B2(n_1488),
.Y(n_2424)
);

AND2x4_ASAP7_75t_L g2425 ( 
.A(n_2041),
.B(n_1044),
.Y(n_2425)
);

AND2x6_ASAP7_75t_L g2426 ( 
.A(n_2096),
.B(n_1039),
.Y(n_2426)
);

AND2x4_ASAP7_75t_L g2427 ( 
.A(n_2043),
.B(n_1288),
.Y(n_2427)
);

OR2x2_ASAP7_75t_L g2428 ( 
.A(n_2032),
.B(n_1596),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2138),
.Y(n_2429)
);

INVx4_ASAP7_75t_L g2430 ( 
.A(n_2086),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2160),
.B(n_1345),
.Y(n_2431)
);

AND2x6_ASAP7_75t_L g2432 ( 
.A(n_2017),
.B(n_1039),
.Y(n_2432)
);

INVx3_ASAP7_75t_L g2433 ( 
.A(n_2078),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2162),
.B(n_1350),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2164),
.B(n_1353),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2052),
.B(n_1450),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2152),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2166),
.B(n_1354),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2167),
.B(n_1356),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_L g2440 ( 
.A(n_2083),
.B(n_1363),
.Y(n_2440)
);

INVx4_ASAP7_75t_L g2441 ( 
.A(n_2087),
.Y(n_2441)
);

INVx3_ASAP7_75t_L g2442 ( 
.A(n_1986),
.Y(n_2442)
);

OR2x2_ASAP7_75t_L g2443 ( 
.A(n_1992),
.B(n_1611),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2159),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_L g2445 ( 
.A(n_2136),
.B(n_1365),
.Y(n_2445)
);

AND2x4_ASAP7_75t_L g2446 ( 
.A(n_1978),
.B(n_1512),
.Y(n_2446)
);

NOR2xp33_ASAP7_75t_L g2447 ( 
.A(n_2145),
.B(n_1374),
.Y(n_2447)
);

AND2x4_ASAP7_75t_L g2448 ( 
.A(n_1982),
.B(n_1601),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2183),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2022),
.Y(n_2450)
);

BUFx4f_ASAP7_75t_L g2451 ( 
.A(n_1986),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2025),
.Y(n_2452)
);

AOI22xp5_ASAP7_75t_L g2453 ( 
.A1(n_2149),
.A2(n_1383),
.B1(n_1385),
.B2(n_1377),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_2154),
.B(n_1391),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2141),
.B(n_1392),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2025),
.Y(n_2456)
);

INVx4_ASAP7_75t_L g2457 ( 
.A(n_2089),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2142),
.B(n_1396),
.Y(n_2458)
);

INVx3_ASAP7_75t_L g2459 ( 
.A(n_1988),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2072),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2069),
.Y(n_2461)
);

OR2x2_ASAP7_75t_L g2462 ( 
.A(n_2058),
.B(n_1397),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2074),
.Y(n_2463)
);

INVx3_ASAP7_75t_L g2464 ( 
.A(n_1988),
.Y(n_2464)
);

OR2x2_ASAP7_75t_L g2465 ( 
.A(n_2059),
.B(n_1400),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2170),
.B(n_1405),
.Y(n_2466)
);

INVx1_ASAP7_75t_SL g2467 ( 
.A(n_2199),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2076),
.Y(n_2468)
);

AND2x6_ASAP7_75t_L g2469 ( 
.A(n_2068),
.B(n_1039),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2175),
.B(n_1406),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2082),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2093),
.B(n_1585),
.Y(n_2472)
);

AND2x4_ASAP7_75t_L g2473 ( 
.A(n_1983),
.B(n_1990),
.Y(n_2473)
);

AO22x2_ASAP7_75t_L g2474 ( 
.A1(n_2240),
.A2(n_1071),
.B1(n_1085),
.B2(n_1070),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2176),
.B(n_1409),
.Y(n_2475)
);

AND2x4_ASAP7_75t_L g2476 ( 
.A(n_2015),
.B(n_1087),
.Y(n_2476)
);

BUFx3_ASAP7_75t_L g2477 ( 
.A(n_2094),
.Y(n_2477)
);

INVx4_ASAP7_75t_L g2478 ( 
.A(n_2099),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2180),
.Y(n_2479)
);

NOR3xp33_ASAP7_75t_L g2480 ( 
.A(n_2033),
.B(n_1413),
.C(n_1412),
.Y(n_2480)
);

NAND2xp33_ASAP7_75t_L g2481 ( 
.A(n_2108),
.B(n_1107),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2095),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2056),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_1980),
.B(n_1423),
.Y(n_2484)
);

BUFx3_ASAP7_75t_L g2485 ( 
.A(n_2203),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_2204),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2090),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2070),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2223),
.Y(n_2489)
);

BUFx3_ASAP7_75t_L g2490 ( 
.A(n_2208),
.Y(n_2490)
);

AND2x2_ASAP7_75t_SL g2491 ( 
.A(n_2228),
.B(n_2234),
.Y(n_2491)
);

INVx3_ASAP7_75t_L g2492 ( 
.A(n_2018),
.Y(n_2492)
);

AND2x2_ASAP7_75t_SL g2493 ( 
.A(n_2241),
.B(n_1563),
.Y(n_2493)
);

AND2x6_ASAP7_75t_L g2494 ( 
.A(n_2084),
.B(n_1039),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2091),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2092),
.Y(n_2496)
);

BUFx6f_ASAP7_75t_L g2497 ( 
.A(n_2210),
.Y(n_2497)
);

INVx1_ASAP7_75t_SL g2498 ( 
.A(n_2080),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2042),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2179),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2214),
.Y(n_2501)
);

INVx6_ASAP7_75t_L g2502 ( 
.A(n_2207),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2042),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2181),
.B(n_1427),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2212),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2102),
.B(n_1585),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2054),
.B(n_1585),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_SL g2508 ( 
.A(n_2048),
.B(n_1431),
.Y(n_2508)
);

CKINVDCx8_ASAP7_75t_R g2509 ( 
.A(n_2034),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2222),
.Y(n_2510)
);

NAND2x1p5_ASAP7_75t_L g2511 ( 
.A(n_2139),
.B(n_1441),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2222),
.Y(n_2512)
);

AND2x4_ASAP7_75t_L g2513 ( 
.A(n_2073),
.B(n_1098),
.Y(n_2513)
);

BUFx3_ASAP7_75t_L g2514 ( 
.A(n_2215),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2211),
.Y(n_2515)
);

INVx8_ASAP7_75t_L g2516 ( 
.A(n_2140),
.Y(n_2516)
);

BUFx4f_ASAP7_75t_L g2517 ( 
.A(n_2047),
.Y(n_2517)
);

INVx4_ASAP7_75t_L g2518 ( 
.A(n_2218),
.Y(n_2518)
);

AND2x4_ASAP7_75t_L g2519 ( 
.A(n_2046),
.B(n_1101),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2039),
.B(n_1435),
.Y(n_2520)
);

INVx4_ASAP7_75t_L g2521 ( 
.A(n_2219),
.Y(n_2521)
);

NOR2xp33_ASAP7_75t_L g2522 ( 
.A(n_2050),
.B(n_1443),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2220),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2213),
.Y(n_2524)
);

AND2x6_ASAP7_75t_L g2525 ( 
.A(n_2217),
.B(n_1117),
.Y(n_2525)
);

AND2x4_ASAP7_75t_L g2526 ( 
.A(n_2060),
.B(n_1109),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2221),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_SL g2528 ( 
.A(n_2038),
.B(n_1447),
.Y(n_2528)
);

INVx1_ASAP7_75t_SL g2529 ( 
.A(n_2053),
.Y(n_2529)
);

BUFx6f_ASAP7_75t_L g2530 ( 
.A(n_2036),
.Y(n_2530)
);

BUFx6f_ASAP7_75t_L g2531 ( 
.A(n_2205),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2055),
.Y(n_2532)
);

INVx4_ASAP7_75t_L g2533 ( 
.A(n_2065),
.Y(n_2533)
);

AND2x6_ASAP7_75t_L g2534 ( 
.A(n_2206),
.B(n_1117),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2066),
.Y(n_2535)
);

BUFx6f_ASAP7_75t_L g2536 ( 
.A(n_2209),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2071),
.B(n_1448),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2146),
.Y(n_2538)
);

INVx3_ASAP7_75t_L g2539 ( 
.A(n_1985),
.Y(n_2539)
);

BUFx6f_ASAP7_75t_L g2540 ( 
.A(n_1985),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2172),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2146),
.Y(n_2542)
);

NAND2xp33_ASAP7_75t_SL g2543 ( 
.A(n_2085),
.B(n_1459),
.Y(n_2543)
);

INVx4_ASAP7_75t_L g2544 ( 
.A(n_1976),
.Y(n_2544)
);

INVx3_ASAP7_75t_L g2545 ( 
.A(n_1985),
.Y(n_2545)
);

AND2x6_ASAP7_75t_L g2546 ( 
.A(n_2044),
.B(n_1117),
.Y(n_2546)
);

INVx3_ASAP7_75t_L g2547 ( 
.A(n_1985),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2057),
.B(n_1602),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2131),
.B(n_1467),
.Y(n_2549)
);

INVx1_ASAP7_75t_SL g2550 ( 
.A(n_2189),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2172),
.Y(n_2551)
);

NOR2xp33_ASAP7_75t_L g2552 ( 
.A(n_2124),
.B(n_1469),
.Y(n_2552)
);

CKINVDCx5p33_ASAP7_75t_R g2553 ( 
.A(n_2021),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2146),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2173),
.Y(n_2555)
);

INVxp67_ASAP7_75t_SL g2556 ( 
.A(n_2189),
.Y(n_2556)
);

INVx3_ASAP7_75t_L g2557 ( 
.A(n_1985),
.Y(n_2557)
);

OR2x2_ASAP7_75t_L g2558 ( 
.A(n_2173),
.B(n_1471),
.Y(n_2558)
);

AND2x4_ASAP7_75t_L g2559 ( 
.A(n_2062),
.B(n_1151),
.Y(n_2559)
);

BUFx2_ASAP7_75t_L g2560 ( 
.A(n_2177),
.Y(n_2560)
);

AND2x6_ASAP7_75t_L g2561 ( 
.A(n_2044),
.B(n_1117),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2057),
.B(n_1602),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_SL g2563 ( 
.A(n_2131),
.B(n_1475),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2172),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2131),
.B(n_1479),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2172),
.Y(n_2566)
);

BUFx10_ASAP7_75t_L g2567 ( 
.A(n_2005),
.Y(n_2567)
);

BUFx6f_ASAP7_75t_L g2568 ( 
.A(n_1985),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2146),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2172),
.Y(n_2570)
);

NAND2x1p5_ASAP7_75t_L g2571 ( 
.A(n_2027),
.B(n_1449),
.Y(n_2571)
);

INVx3_ASAP7_75t_L g2572 ( 
.A(n_1985),
.Y(n_2572)
);

AND2x2_ASAP7_75t_SL g2573 ( 
.A(n_2016),
.B(n_1563),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2172),
.Y(n_2574)
);

AO22x2_ASAP7_75t_L g2575 ( 
.A1(n_1998),
.A2(n_1182),
.B1(n_1186),
.B2(n_1153),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_SL g2576 ( 
.A(n_2131),
.B(n_1480),
.Y(n_2576)
);

BUFx3_ASAP7_75t_L g2577 ( 
.A(n_2201),
.Y(n_2577)
);

AND2x4_ASAP7_75t_L g2578 ( 
.A(n_2062),
.B(n_1201),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2131),
.B(n_1481),
.Y(n_2579)
);

CKINVDCx20_ASAP7_75t_R g2580 ( 
.A(n_2035),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2057),
.B(n_1482),
.Y(n_2581)
);

BUFx3_ASAP7_75t_L g2582 ( 
.A(n_2201),
.Y(n_2582)
);

OR2x2_ASAP7_75t_L g2583 ( 
.A(n_2173),
.B(n_1486),
.Y(n_2583)
);

INVx4_ASAP7_75t_L g2584 ( 
.A(n_1976),
.Y(n_2584)
);

NOR2xp33_ASAP7_75t_L g2585 ( 
.A(n_2124),
.B(n_1487),
.Y(n_2585)
);

INVx4_ASAP7_75t_L g2586 ( 
.A(n_1976),
.Y(n_2586)
);

INVx5_ASAP7_75t_L g2587 ( 
.A(n_2247),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2146),
.Y(n_2588)
);

AND2x6_ASAP7_75t_L g2589 ( 
.A(n_2044),
.B(n_1559),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2057),
.B(n_1490),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2131),
.B(n_1492),
.Y(n_2591)
);

BUFx3_ASAP7_75t_L g2592 ( 
.A(n_2201),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2172),
.Y(n_2593)
);

NAND3xp33_ASAP7_75t_L g2594 ( 
.A(n_2124),
.B(n_1500),
.C(n_1495),
.Y(n_2594)
);

INVx6_ASAP7_75t_L g2595 ( 
.A(n_1985),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2131),
.B(n_1501),
.Y(n_2596)
);

INVx3_ASAP7_75t_L g2597 ( 
.A(n_1985),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2146),
.Y(n_2598)
);

INVx3_ASAP7_75t_L g2599 ( 
.A(n_1985),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2146),
.Y(n_2600)
);

BUFx3_ASAP7_75t_L g2601 ( 
.A(n_2201),
.Y(n_2601)
);

OR2x6_ASAP7_75t_L g2602 ( 
.A(n_2242),
.B(n_1042),
.Y(n_2602)
);

NOR2xp33_ASAP7_75t_L g2603 ( 
.A(n_2124),
.B(n_1502),
.Y(n_2603)
);

INVxp67_ASAP7_75t_SL g2604 ( 
.A(n_2189),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_2021),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2172),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2172),
.Y(n_2607)
);

BUFx6f_ASAP7_75t_L g2608 ( 
.A(n_1985),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2262),
.B(n_1509),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2541),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2551),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2266),
.B(n_1513),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_2581),
.B(n_1516),
.Y(n_2613)
);

AND2x6_ASAP7_75t_L g2614 ( 
.A(n_2540),
.B(n_1559),
.Y(n_2614)
);

OAI22xp5_ASAP7_75t_L g2615 ( 
.A1(n_2482),
.A2(n_1524),
.B1(n_1525),
.B2(n_1519),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2564),
.Y(n_2616)
);

AND2x4_ASAP7_75t_L g2617 ( 
.A(n_2540),
.B(n_1207),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2257),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2462),
.B(n_2465),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_SL g2620 ( 
.A(n_2568),
.B(n_1532),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2271),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_2568),
.B(n_1538),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2296),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2300),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2305),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2269),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2267),
.B(n_1552),
.Y(n_2627)
);

NAND3xp33_ASAP7_75t_L g2628 ( 
.A(n_2328),
.B(n_2344),
.C(n_2552),
.Y(n_2628)
);

BUFx2_ASAP7_75t_L g2629 ( 
.A(n_2404),
.Y(n_2629)
);

BUFx3_ASAP7_75t_L g2630 ( 
.A(n_2608),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2308),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2590),
.B(n_1553),
.Y(n_2632)
);

HB1xp67_ASAP7_75t_L g2633 ( 
.A(n_2287),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2316),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2319),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2274),
.Y(n_2636)
);

NAND2x1p5_ASAP7_75t_L g2637 ( 
.A(n_2287),
.B(n_1559),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2323),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2566),
.Y(n_2639)
);

AND2x4_ASAP7_75t_L g2640 ( 
.A(n_2608),
.B(n_1208),
.Y(n_2640)
);

AND2x4_ASAP7_75t_L g2641 ( 
.A(n_2291),
.B(n_1215),
.Y(n_2641)
);

AOI22xp33_ASAP7_75t_L g2642 ( 
.A1(n_2526),
.A2(n_1557),
.B1(n_1558),
.B2(n_1556),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2570),
.Y(n_2643)
);

INVx5_ASAP7_75t_L g2644 ( 
.A(n_2595),
.Y(n_2644)
);

INVxp67_ASAP7_75t_L g2645 ( 
.A(n_2273),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2585),
.B(n_1571),
.Y(n_2646)
);

NAND2xp33_ASAP7_75t_L g2647 ( 
.A(n_2426),
.B(n_1603),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2363),
.Y(n_2648)
);

AND2x4_ASAP7_75t_L g2649 ( 
.A(n_2301),
.B(n_1219),
.Y(n_2649)
);

AO22x2_ASAP7_75t_L g2650 ( 
.A1(n_2324),
.A2(n_1470),
.B1(n_1472),
.B2(n_1453),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2375),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2380),
.Y(n_2652)
);

INVx3_ASAP7_75t_L g2653 ( 
.A(n_2355),
.Y(n_2653)
);

HB1xp67_ASAP7_75t_L g2654 ( 
.A(n_2587),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2574),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2396),
.Y(n_2656)
);

OR2x2_ASAP7_75t_L g2657 ( 
.A(n_2498),
.B(n_1586),
.Y(n_2657)
);

INVxp67_ASAP7_75t_L g2658 ( 
.A(n_2333),
.Y(n_2658)
);

BUFx6f_ASAP7_75t_L g2659 ( 
.A(n_2307),
.Y(n_2659)
);

HB1xp67_ASAP7_75t_L g2660 ( 
.A(n_2587),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2267),
.B(n_2261),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2450),
.Y(n_2662)
);

OAI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2391),
.A2(n_1595),
.B1(n_1607),
.B2(n_1587),
.Y(n_2663)
);

A2O1A1Ixp33_ASAP7_75t_L g2664 ( 
.A1(n_2369),
.A2(n_1478),
.B(n_1494),
.C(n_1477),
.Y(n_2664)
);

OA22x2_ASAP7_75t_L g2665 ( 
.A1(n_2303),
.A2(n_1608),
.B1(n_1017),
.B2(n_1019),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2593),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2549),
.B(n_1497),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2603),
.B(n_1104),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2606),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2607),
.Y(n_2670)
);

NAND2xp33_ASAP7_75t_L g2671 ( 
.A(n_2426),
.B(n_1107),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2331),
.Y(n_2672)
);

INVxp67_ASAP7_75t_L g2673 ( 
.A(n_2390),
.Y(n_2673)
);

BUFx8_ASAP7_75t_L g2674 ( 
.A(n_2320),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_L g2675 ( 
.A(n_2335),
.B(n_1026),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2364),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2327),
.B(n_1104),
.Y(n_2677)
);

AO22x2_ASAP7_75t_L g2678 ( 
.A1(n_2550),
.A2(n_1510),
.B1(n_1522),
.B2(n_1503),
.Y(n_2678)
);

AND2x4_ASAP7_75t_L g2679 ( 
.A(n_2259),
.B(n_1221),
.Y(n_2679)
);

INVxp67_ASAP7_75t_L g2680 ( 
.A(n_2555),
.Y(n_2680)
);

AO22x2_ASAP7_75t_L g2681 ( 
.A1(n_2556),
.A2(n_1539),
.B1(n_1542),
.B2(n_1523),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2365),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2371),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2373),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2565),
.B(n_1561),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2377),
.Y(n_2686)
);

NAND2x1p5_ASAP7_75t_L g2687 ( 
.A(n_2350),
.B(n_1610),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2386),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_SL g2689 ( 
.A(n_2416),
.B(n_1600),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2388),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2392),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2393),
.Y(n_2692)
);

BUFx2_ASAP7_75t_L g2693 ( 
.A(n_2604),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2522),
.B(n_1030),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2395),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2413),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2405),
.Y(n_2697)
);

HB1xp67_ASAP7_75t_L g2698 ( 
.A(n_2511),
.Y(n_2698)
);

AOI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_2445),
.A2(n_1046),
.B1(n_1048),
.B2(n_1031),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2411),
.Y(n_2700)
);

BUFx8_ASAP7_75t_L g2701 ( 
.A(n_2383),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2419),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2414),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2420),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2429),
.Y(n_2705)
);

INVx4_ASAP7_75t_L g2706 ( 
.A(n_2407),
.Y(n_2706)
);

BUFx6f_ASAP7_75t_L g2707 ( 
.A(n_2307),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2449),
.Y(n_2708)
);

NAND2x1p5_ASAP7_75t_L g2709 ( 
.A(n_2281),
.B(n_1569),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2575),
.B(n_1112),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2437),
.Y(n_2711)
);

HB1xp67_ASAP7_75t_L g2712 ( 
.A(n_2571),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2444),
.Y(n_2713)
);

BUFx3_ASAP7_75t_L g2714 ( 
.A(n_2292),
.Y(n_2714)
);

INVxp67_ASAP7_75t_L g2715 ( 
.A(n_2443),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2579),
.B(n_1575),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2346),
.Y(n_2717)
);

AOI22xp33_ASAP7_75t_L g2718 ( 
.A1(n_2519),
.A2(n_1281),
.B1(n_1290),
.B2(n_1112),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2370),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2256),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2538),
.Y(n_2721)
);

BUFx2_ASAP7_75t_L g2722 ( 
.A(n_2297),
.Y(n_2722)
);

AND2x4_ASAP7_75t_L g2723 ( 
.A(n_2280),
.B(n_1276),
.Y(n_2723)
);

AND2x4_ASAP7_75t_L g2724 ( 
.A(n_2539),
.B(n_1277),
.Y(n_2724)
);

AND2x4_ASAP7_75t_SL g2725 ( 
.A(n_2407),
.B(n_1281),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2349),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2591),
.B(n_2596),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2505),
.Y(n_2728)
);

NAND2x1p5_ASAP7_75t_L g2729 ( 
.A(n_2283),
.B(n_1588),
.Y(n_2729)
);

CKINVDCx5p33_ASAP7_75t_R g2730 ( 
.A(n_2408),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2286),
.B(n_1594),
.Y(n_2731)
);

OAI22xp5_ASAP7_75t_L g2732 ( 
.A1(n_2276),
.A2(n_1598),
.B1(n_1066),
.B2(n_1069),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2546),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2542),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2546),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2554),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2558),
.B(n_1072),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2561),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2569),
.Y(n_2739)
);

OAI221xp5_ASAP7_75t_L g2740 ( 
.A1(n_2382),
.A2(n_1076),
.B1(n_1078),
.B2(n_1074),
.C(n_1073),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2588),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2561),
.Y(n_2742)
);

OAI221xp5_ASAP7_75t_L g2743 ( 
.A1(n_2520),
.A2(n_2326),
.B1(n_2310),
.B2(n_2453),
.C(n_2293),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2598),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2561),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2589),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2575),
.B(n_2275),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2330),
.B(n_2304),
.Y(n_2748)
);

OR2x2_ASAP7_75t_L g2749 ( 
.A(n_2264),
.B(n_1086),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_2567),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2313),
.B(n_1290),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2600),
.Y(n_2752)
);

NOR2xp33_ASAP7_75t_SL g2753 ( 
.A(n_2491),
.B(n_1088),
.Y(n_2753)
);

NOR2x1p5_ASAP7_75t_L g2754 ( 
.A(n_2553),
.B(n_1090),
.Y(n_2754)
);

NOR2xp33_ASAP7_75t_L g2755 ( 
.A(n_2583),
.B(n_1092),
.Y(n_2755)
);

INVxp67_ASAP7_75t_L g2756 ( 
.A(n_2278),
.Y(n_2756)
);

BUFx3_ASAP7_75t_L g2757 ( 
.A(n_2299),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2589),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2548),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2355),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2562),
.Y(n_2761)
);

A2O1A1Ixp33_ASAP7_75t_L g2762 ( 
.A1(n_2367),
.A2(n_2403),
.B(n_2503),
.C(n_2499),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2483),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2545),
.B(n_1278),
.Y(n_2764)
);

AND2x4_ASAP7_75t_L g2765 ( 
.A(n_2547),
.B(n_1299),
.Y(n_2765)
);

NOR2xp33_ASAP7_75t_L g2766 ( 
.A(n_2379),
.B(n_1105),
.Y(n_2766)
);

INVx3_ASAP7_75t_L g2767 ( 
.A(n_2360),
.Y(n_2767)
);

AND2x4_ASAP7_75t_L g2768 ( 
.A(n_2557),
.B(n_1300),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2360),
.Y(n_2769)
);

NOR2xp33_ASAP7_75t_L g2770 ( 
.A(n_2529),
.B(n_1106),
.Y(n_2770)
);

AO22x2_ASAP7_75t_L g2771 ( 
.A1(n_2532),
.A2(n_1316),
.B1(n_1318),
.B2(n_1303),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2343),
.B(n_1121),
.Y(n_2772)
);

NAND2x1p5_ASAP7_75t_L g2773 ( 
.A(n_2288),
.B(n_1116),
.Y(n_2773)
);

BUFx2_ASAP7_75t_L g2774 ( 
.A(n_2577),
.Y(n_2774)
);

HB1xp67_ASAP7_75t_L g2775 ( 
.A(n_2582),
.Y(n_2775)
);

BUFx2_ASAP7_75t_L g2776 ( 
.A(n_2592),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2378),
.Y(n_2777)
);

AND2x4_ASAP7_75t_L g2778 ( 
.A(n_2572),
.B(n_1320),
.Y(n_2778)
);

INVxp67_ASAP7_75t_L g2779 ( 
.A(n_2315),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2479),
.Y(n_2780)
);

NAND2x1p5_ASAP7_75t_L g2781 ( 
.A(n_2544),
.B(n_1116),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2378),
.Y(n_2782)
);

OAI221xp5_ASAP7_75t_L g2783 ( 
.A1(n_2409),
.A2(n_2435),
.B1(n_2438),
.B2(n_2434),
.C(n_2431),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2397),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2460),
.Y(n_2785)
);

BUFx4f_ASAP7_75t_L g2786 ( 
.A(n_2348),
.Y(n_2786)
);

OAI21xp33_ASAP7_75t_L g2787 ( 
.A1(n_2406),
.A2(n_1127),
.B(n_1122),
.Y(n_2787)
);

BUFx6f_ASAP7_75t_L g2788 ( 
.A(n_2309),
.Y(n_2788)
);

INVxp67_ASAP7_75t_L g2789 ( 
.A(n_2602),
.Y(n_2789)
);

CKINVDCx5p33_ASAP7_75t_R g2790 ( 
.A(n_2605),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2384),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2493),
.B(n_1329),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2474),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2474),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2384),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2389),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2394),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2352),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2285),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2488),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2285),
.Y(n_2801)
);

BUFx2_ASAP7_75t_L g2802 ( 
.A(n_2601),
.Y(n_2802)
);

AO22x2_ASAP7_75t_L g2803 ( 
.A1(n_2535),
.A2(n_1328),
.B1(n_1333),
.B2(n_1322),
.Y(n_2803)
);

INVx3_ASAP7_75t_L g2804 ( 
.A(n_2389),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2399),
.Y(n_2805)
);

AOI22xp33_ASAP7_75t_L g2806 ( 
.A1(n_2480),
.A2(n_1562),
.B1(n_1329),
.B2(n_1132),
.Y(n_2806)
);

NOR2xp33_ASAP7_75t_L g2807 ( 
.A(n_2340),
.B(n_1142),
.Y(n_2807)
);

OAI22xp33_ASAP7_75t_L g2808 ( 
.A1(n_2528),
.A2(n_2354),
.B1(n_2265),
.B2(n_2258),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2285),
.B(n_1144),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2439),
.B(n_1147),
.Y(n_2810)
);

BUFx3_ASAP7_75t_L g2811 ( 
.A(n_2486),
.Y(n_2811)
);

BUFx6f_ASAP7_75t_L g2812 ( 
.A(n_2309),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2399),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2495),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2496),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2563),
.Y(n_2816)
);

NAND2x1p5_ASAP7_75t_L g2817 ( 
.A(n_2584),
.B(n_1116),
.Y(n_2817)
);

BUFx6f_ASAP7_75t_L g2818 ( 
.A(n_2426),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2332),
.B(n_1171),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2507),
.B(n_1175),
.Y(n_2820)
);

AO22x2_ASAP7_75t_L g2821 ( 
.A1(n_2467),
.A2(n_1358),
.B1(n_1367),
.B2(n_1349),
.Y(n_2821)
);

NOR2xp33_ASAP7_75t_L g2822 ( 
.A(n_2263),
.B(n_2268),
.Y(n_2822)
);

NAND2x1p5_ASAP7_75t_L g2823 ( 
.A(n_2586),
.B(n_1180),
.Y(n_2823)
);

AOI22x1_ASAP7_75t_L g2824 ( 
.A1(n_2290),
.A2(n_1043),
.B1(n_1060),
.B2(n_1042),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2576),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2461),
.Y(n_2826)
);

AOI22xp5_ASAP7_75t_L g2827 ( 
.A1(n_2447),
.A2(n_2454),
.B1(n_2358),
.B2(n_2347),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2463),
.Y(n_2828)
);

INVxp67_ASAP7_75t_L g2829 ( 
.A(n_2602),
.Y(n_2829)
);

AOI211xp5_ASAP7_75t_L g2830 ( 
.A1(n_2412),
.A2(n_2361),
.B(n_2402),
.C(n_2366),
.Y(n_2830)
);

A2O1A1Ixp33_ASAP7_75t_L g2831 ( 
.A1(n_2424),
.A2(n_1421),
.B(n_1426),
.C(n_1402),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2468),
.Y(n_2832)
);

AND2x4_ASAP7_75t_L g2833 ( 
.A(n_2597),
.B(n_1434),
.Y(n_2833)
);

INVxp67_ASAP7_75t_L g2834 ( 
.A(n_2387),
.Y(n_2834)
);

BUFx8_ASAP7_75t_L g2835 ( 
.A(n_2348),
.Y(n_2835)
);

INVxp67_ASAP7_75t_L g2836 ( 
.A(n_2410),
.Y(n_2836)
);

NAND2x1p5_ASAP7_75t_L g2837 ( 
.A(n_2599),
.B(n_1180),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2515),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2524),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2471),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2487),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2295),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2466),
.B(n_1179),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2298),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2298),
.Y(n_2845)
);

NAND2x1p5_ASAP7_75t_L g2846 ( 
.A(n_2345),
.B(n_1180),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2484),
.Y(n_2847)
);

NOR2xp33_ASAP7_75t_L g2848 ( 
.A(n_2284),
.B(n_1183),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2298),
.Y(n_2849)
);

CKINVDCx5p33_ASAP7_75t_R g2850 ( 
.A(n_2516),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2506),
.B(n_1562),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2500),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2489),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2277),
.Y(n_2854)
);

NAND2x1p5_ASAP7_75t_L g2855 ( 
.A(n_2381),
.B(n_1180),
.Y(n_2855)
);

NAND2x1p5_ASAP7_75t_L g2856 ( 
.A(n_2486),
.B(n_1232),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2470),
.B(n_1203),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2430),
.B(n_2441),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2475),
.B(n_1214),
.Y(n_2859)
);

INVx4_ASAP7_75t_L g2860 ( 
.A(n_2497),
.Y(n_2860)
);

OR2x6_ASAP7_75t_L g2861 ( 
.A(n_2516),
.B(n_1043),
.Y(n_2861)
);

NAND2x1p5_ASAP7_75t_L g2862 ( 
.A(n_2497),
.B(n_1232),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2329),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2282),
.Y(n_2864)
);

INVxp67_ASAP7_75t_L g2865 ( 
.A(n_2560),
.Y(n_2865)
);

BUFx8_ASAP7_75t_L g2866 ( 
.A(n_2376),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2436),
.B(n_2423),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2339),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_2517),
.B(n_1599),
.Y(n_2869)
);

AO22x2_ASAP7_75t_L g2870 ( 
.A1(n_2272),
.A2(n_1442),
.B1(n_1446),
.B2(n_1439),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2289),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2508),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2504),
.B(n_1238),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2510),
.Y(n_2874)
);

NOR2xp33_ASAP7_75t_L g2875 ( 
.A(n_2440),
.B(n_1240),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2442),
.Y(n_2876)
);

AND2x2_ASAP7_75t_L g2877 ( 
.A(n_2472),
.B(n_2573),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2459),
.Y(n_2878)
);

AO22x2_ASAP7_75t_L g2879 ( 
.A1(n_2533),
.A2(n_1458),
.B1(n_1461),
.B2(n_1457),
.Y(n_2879)
);

OR2x2_ASAP7_75t_L g2880 ( 
.A(n_2279),
.B(n_1251),
.Y(n_2880)
);

BUFx2_ASAP7_75t_L g2881 ( 
.A(n_2415),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2464),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2512),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2455),
.B(n_1253),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2531),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2351),
.Y(n_2886)
);

NAND2x1p5_ASAP7_75t_L g2887 ( 
.A(n_2501),
.B(n_2322),
.Y(n_2887)
);

BUFx8_ASAP7_75t_L g2888 ( 
.A(n_2338),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2433),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2359),
.Y(n_2890)
);

OAI221xp5_ASAP7_75t_L g2891 ( 
.A1(n_2458),
.A2(n_1272),
.B1(n_1280),
.B2(n_1271),
.C(n_1255),
.Y(n_2891)
);

NAND2x1p5_ASAP7_75t_L g2892 ( 
.A(n_2501),
.B(n_1232),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_2401),
.B(n_1282),
.Y(n_2893)
);

INVxp67_ASAP7_75t_L g2894 ( 
.A(n_2425),
.Y(n_2894)
);

AOI22xp5_ASAP7_75t_L g2895 ( 
.A1(n_2353),
.A2(n_1286),
.B1(n_1292),
.B2(n_1291),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2531),
.Y(n_2896)
);

BUFx8_ASAP7_75t_L g2897 ( 
.A(n_2314),
.Y(n_2897)
);

BUFx6f_ASAP7_75t_L g2898 ( 
.A(n_2432),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_L g2899 ( 
.A(n_2594),
.B(n_1298),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2536),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2536),
.Y(n_2901)
);

AO22x2_ASAP7_75t_L g2902 ( 
.A1(n_2398),
.A2(n_1465),
.B1(n_1473),
.B2(n_1464),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2523),
.Y(n_2903)
);

AND2x4_ASAP7_75t_L g2904 ( 
.A(n_2457),
.B(n_2478),
.Y(n_2904)
);

NOR2xp33_ASAP7_75t_SL g2905 ( 
.A(n_2421),
.B(n_2422),
.Y(n_2905)
);

AOI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2543),
.A2(n_2513),
.B1(n_2578),
.B2(n_2559),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2527),
.Y(n_2907)
);

AO22x2_ASAP7_75t_L g2908 ( 
.A1(n_2368),
.A2(n_1483),
.B1(n_1484),
.B2(n_1474),
.Y(n_2908)
);

OAI22xp5_ASAP7_75t_SL g2909 ( 
.A1(n_2400),
.A2(n_1568),
.B1(n_1573),
.B2(n_1566),
.Y(n_2909)
);

NAND2x1p5_ASAP7_75t_L g2910 ( 
.A(n_2485),
.B(n_1232),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2417),
.B(n_1301),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2537),
.B(n_1304),
.Y(n_2912)
);

AO22x2_ASAP7_75t_L g2913 ( 
.A1(n_2427),
.A2(n_1514),
.B1(n_1515),
.B2(n_1507),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2502),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2502),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2306),
.Y(n_2916)
);

INVxp67_ASAP7_75t_L g2917 ( 
.A(n_2321),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2451),
.Y(n_2918)
);

AND2x2_ASAP7_75t_L g2919 ( 
.A(n_2446),
.B(n_1311),
.Y(n_2919)
);

AO22x2_ASAP7_75t_L g2920 ( 
.A1(n_2337),
.A2(n_1528),
.B1(n_1536),
.B2(n_1526),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2306),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2306),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2342),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_SL g2924 ( 
.A(n_2448),
.B(n_1550),
.Y(n_2924)
);

AO22x2_ASAP7_75t_L g2925 ( 
.A1(n_2357),
.A2(n_1544),
.B1(n_1549),
.B2(n_1540),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2362),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2362),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_SL g2928 ( 
.A(n_2477),
.B(n_1576),
.Y(n_2928)
);

AND3x4_ASAP7_75t_L g2929 ( 
.A(n_2473),
.B(n_1065),
.C(n_1060),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2362),
.Y(n_2930)
);

INVx2_ASAP7_75t_SL g2931 ( 
.A(n_2490),
.Y(n_2931)
);

AOI22xp33_ASAP7_75t_L g2932 ( 
.A1(n_2476),
.A2(n_1323),
.B1(n_1324),
.B2(n_1321),
.Y(n_2932)
);

HB1xp67_ASAP7_75t_L g2933 ( 
.A(n_2341),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2374),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2374),
.Y(n_2935)
);

OAI221xp5_ASAP7_75t_L g2936 ( 
.A1(n_2336),
.A2(n_1351),
.B1(n_1352),
.B2(n_1347),
.C(n_1344),
.Y(n_2936)
);

BUFx6f_ASAP7_75t_L g2937 ( 
.A(n_2432),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_SL g2938 ( 
.A(n_2518),
.B(n_1546),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2374),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2294),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2294),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2336),
.Y(n_2942)
);

AND2x4_ASAP7_75t_L g2943 ( 
.A(n_2418),
.B(n_1564),
.Y(n_2943)
);

AND2x4_ASAP7_75t_L g2944 ( 
.A(n_2514),
.B(n_1572),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2481),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2469),
.Y(n_2946)
);

AND2x4_ASAP7_75t_L g2947 ( 
.A(n_2521),
.B(n_1582),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_SL g2948 ( 
.A(n_2318),
.B(n_1547),
.Y(n_2948)
);

BUFx10_ASAP7_75t_L g2949 ( 
.A(n_2270),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2469),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2469),
.Y(n_2951)
);

AO22x2_ASAP7_75t_L g2952 ( 
.A1(n_2325),
.A2(n_1167),
.B1(n_1192),
.B2(n_1065),
.Y(n_2952)
);

BUFx2_ASAP7_75t_L g2953 ( 
.A(n_2334),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2494),
.Y(n_2954)
);

NOR3xp33_ASAP7_75t_L g2955 ( 
.A(n_2492),
.B(n_1368),
.C(n_1357),
.Y(n_2955)
);

OAI22xp5_ASAP7_75t_SL g2956 ( 
.A1(n_2509),
.A2(n_1605),
.B1(n_1606),
.B2(n_1597),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2494),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2494),
.Y(n_2958)
);

INVxp67_ASAP7_75t_L g2959 ( 
.A(n_2372),
.Y(n_2959)
);

INVxp67_ASAP7_75t_L g2960 ( 
.A(n_2385),
.Y(n_2960)
);

BUFx6f_ASAP7_75t_L g2961 ( 
.A(n_2432),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2525),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2525),
.Y(n_2963)
);

AND2x4_ASAP7_75t_L g2964 ( 
.A(n_2530),
.B(n_1167),
.Y(n_2964)
);

AOI22xp5_ASAP7_75t_L g2965 ( 
.A1(n_2530),
.A2(n_1379),
.B1(n_1389),
.B2(n_1380),
.Y(n_2965)
);

OAI221xp5_ASAP7_75t_L g2966 ( 
.A1(n_2356),
.A2(n_1407),
.B1(n_1414),
.B2(n_1404),
.C(n_1393),
.Y(n_2966)
);

INVx2_ASAP7_75t_SL g2967 ( 
.A(n_2525),
.Y(n_2967)
);

NAND2x1p5_ASAP7_75t_L g2968 ( 
.A(n_2302),
.B(n_1296),
.Y(n_2968)
);

A2O1A1Ixp33_ASAP7_75t_L g2969 ( 
.A1(n_2311),
.A2(n_1192),
.B(n_1231),
.C(n_1204),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2534),
.Y(n_2970)
);

OAI22xp33_ASAP7_75t_L g2971 ( 
.A1(n_2312),
.A2(n_1417),
.B1(n_1420),
.B2(n_1416),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2317),
.B(n_1425),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2452),
.B(n_1428),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2456),
.B(n_1437),
.Y(n_2974)
);

NAND2x1p5_ASAP7_75t_L g2975 ( 
.A(n_2534),
.B(n_1296),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2581),
.B(n_1445),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2581),
.B(n_1454),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2257),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2257),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2262),
.B(n_1460),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2262),
.Y(n_2981)
);

NAND2x1p5_ASAP7_75t_L g2982 ( 
.A(n_2287),
.B(n_1296),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2581),
.B(n_1466),
.Y(n_2983)
);

BUFx8_ASAP7_75t_L g2984 ( 
.A(n_2540),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2257),
.Y(n_2985)
);

AO22x2_ASAP7_75t_L g2986 ( 
.A1(n_2324),
.A2(n_1231),
.B1(n_1268),
.B2(n_1204),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2262),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2262),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2257),
.Y(n_2989)
);

HB1xp67_ASAP7_75t_L g2990 ( 
.A(n_2287),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2262),
.Y(n_2991)
);

HB1xp67_ASAP7_75t_L g2992 ( 
.A(n_2287),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2257),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2262),
.B(n_1485),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2260),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2581),
.B(n_1489),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2260),
.Y(n_2997)
);

INVx2_ASAP7_75t_SL g2998 ( 
.A(n_2595),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2260),
.Y(n_2999)
);

INVxp67_ASAP7_75t_L g3000 ( 
.A(n_2428),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2260),
.Y(n_3001)
);

CKINVDCx20_ASAP7_75t_R g3002 ( 
.A(n_2580),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2262),
.B(n_1491),
.Y(n_3003)
);

NAND2x1p5_ASAP7_75t_L g3004 ( 
.A(n_2287),
.B(n_1296),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2257),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2262),
.B(n_1498),
.Y(n_3006)
);

NAND2x1p5_ASAP7_75t_L g3007 ( 
.A(n_2287),
.B(n_1268),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2260),
.Y(n_3008)
);

OR2x2_ASAP7_75t_SL g3009 ( 
.A(n_2595),
.B(n_1555),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2257),
.Y(n_3010)
);

AO22x2_ASAP7_75t_L g3011 ( 
.A1(n_2324),
.A2(n_1274),
.B1(n_1293),
.B2(n_1269),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2257),
.Y(n_3012)
);

INVxp67_ASAP7_75t_L g3013 ( 
.A(n_2428),
.Y(n_3013)
);

AND2x4_ASAP7_75t_L g3014 ( 
.A(n_2540),
.B(n_1269),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2257),
.Y(n_3015)
);

AO22x2_ASAP7_75t_L g3016 ( 
.A1(n_2324),
.A2(n_1293),
.B1(n_1339),
.B2(n_1274),
.Y(n_3016)
);

HB1xp67_ASAP7_75t_L g3017 ( 
.A(n_2287),
.Y(n_3017)
);

BUFx2_ASAP7_75t_L g3018 ( 
.A(n_2580),
.Y(n_3018)
);

INVxp67_ASAP7_75t_L g3019 ( 
.A(n_2428),
.Y(n_3019)
);

INVxp67_ASAP7_75t_L g3020 ( 
.A(n_2428),
.Y(n_3020)
);

INVxp67_ASAP7_75t_L g3021 ( 
.A(n_2428),
.Y(n_3021)
);

OR2x2_ASAP7_75t_SL g3022 ( 
.A(n_2595),
.B(n_1555),
.Y(n_3022)
);

HB1xp67_ASAP7_75t_L g3023 ( 
.A(n_2287),
.Y(n_3023)
);

NAND3xp33_ASAP7_75t_L g3024 ( 
.A(n_2328),
.B(n_1527),
.C(n_1521),
.Y(n_3024)
);

BUFx3_ASAP7_75t_L g3025 ( 
.A(n_2540),
.Y(n_3025)
);

OAI22xp5_ASAP7_75t_L g3026 ( 
.A1(n_2482),
.A2(n_1531),
.B1(n_1534),
.B2(n_1530),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_2540),
.B(n_1593),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2260),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2260),
.Y(n_3029)
);

NOR2xp33_ASAP7_75t_L g3030 ( 
.A(n_2462),
.B(n_1535),
.Y(n_3030)
);

AOI22xp5_ASAP7_75t_SL g3031 ( 
.A1(n_2580),
.A2(n_1609),
.B1(n_1545),
.B2(n_1386),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2262),
.B(n_1488),
.Y(n_3032)
);

INVx2_ASAP7_75t_SL g3033 ( 
.A(n_2595),
.Y(n_3033)
);

AND2x4_ASAP7_75t_L g3034 ( 
.A(n_2540),
.B(n_1339),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2257),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2260),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2257),
.Y(n_3037)
);

OR2x2_ASAP7_75t_L g3038 ( 
.A(n_2324),
.B(n_1386),
.Y(n_3038)
);

NOR2xp33_ASAP7_75t_L g3039 ( 
.A(n_2462),
.B(n_1468),
.Y(n_3039)
);

OAI22xp33_ASAP7_75t_L g3040 ( 
.A1(n_2303),
.A2(n_1567),
.B1(n_1468),
.B2(n_4),
.Y(n_3040)
);

BUFx3_ASAP7_75t_L g3041 ( 
.A(n_2540),
.Y(n_3041)
);

INVxp67_ASAP7_75t_L g3042 ( 
.A(n_2428),
.Y(n_3042)
);

AOI22xp5_ASAP7_75t_L g3043 ( 
.A1(n_2445),
.A2(n_1613),
.B1(n_1488),
.B2(n_1394),
.Y(n_3043)
);

INVx3_ASAP7_75t_L g3044 ( 
.A(n_2540),
.Y(n_3044)
);

NAND2x1p5_ASAP7_75t_L g3045 ( 
.A(n_2287),
.B(n_3),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2257),
.Y(n_3046)
);

OAI22xp33_ASAP7_75t_SL g3047 ( 
.A1(n_2511),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2260),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_SL g3049 ( 
.A(n_2540),
.B(n_1488),
.Y(n_3049)
);

AND2x4_ASAP7_75t_L g3050 ( 
.A(n_2540),
.B(n_5),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2581),
.B(n_1488),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2260),
.Y(n_3052)
);

AND2x4_ASAP7_75t_L g3053 ( 
.A(n_2540),
.B(n_6),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2260),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2260),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2262),
.B(n_1613),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_SL g3057 ( 
.A(n_2540),
.B(n_1613),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2581),
.B(n_1613),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2260),
.Y(n_3059)
);

BUFx2_ASAP7_75t_L g3060 ( 
.A(n_2580),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2260),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2262),
.B(n_1613),
.Y(n_3062)
);

INVx3_ASAP7_75t_L g3063 ( 
.A(n_2540),
.Y(n_3063)
);

AND2x4_ASAP7_75t_L g3064 ( 
.A(n_2540),
.B(n_6),
.Y(n_3064)
);

OAI22xp5_ASAP7_75t_SL g3065 ( 
.A1(n_2580),
.A2(n_9),
.B1(n_10),
.B2(n_8),
.Y(n_3065)
);

HB1xp67_ASAP7_75t_L g3066 ( 
.A(n_2287),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2262),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2262),
.Y(n_3068)
);

CKINVDCx5p33_ASAP7_75t_R g3069 ( 
.A(n_2580),
.Y(n_3069)
);

AO22x2_ASAP7_75t_L g3070 ( 
.A1(n_2324),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_3070)
);

AND2x4_ASAP7_75t_L g3071 ( 
.A(n_2540),
.B(n_8),
.Y(n_3071)
);

AND2x2_ASAP7_75t_L g3072 ( 
.A(n_2581),
.B(n_1154),
.Y(n_3072)
);

AO22x2_ASAP7_75t_L g3073 ( 
.A1(n_2324),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2260),
.Y(n_3074)
);

AO22x2_ASAP7_75t_L g3075 ( 
.A1(n_2324),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_3075)
);

AND2x2_ASAP7_75t_L g3076 ( 
.A(n_2581),
.B(n_1154),
.Y(n_3076)
);

NAND2x1p5_ASAP7_75t_L g3077 ( 
.A(n_2287),
.B(n_11),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2260),
.Y(n_3078)
);

BUFx4f_ASAP7_75t_L g3079 ( 
.A(n_2540),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2260),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2260),
.Y(n_3081)
);

AOI22xp33_ASAP7_75t_L g3082 ( 
.A1(n_2526),
.A2(n_1456),
.B1(n_1394),
.B2(n_14),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2257),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2257),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2260),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2260),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2260),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2260),
.Y(n_3088)
);

NAND2x1p5_ASAP7_75t_L g3089 ( 
.A(n_2287),
.B(n_12),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2260),
.Y(n_3090)
);

INVx1_ASAP7_75t_SL g3091 ( 
.A(n_2580),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2260),
.Y(n_3092)
);

INVx2_ASAP7_75t_L g3093 ( 
.A(n_2257),
.Y(n_3093)
);

A2O1A1Ixp33_ASAP7_75t_L g3094 ( 
.A1(n_2482),
.A2(n_1456),
.B(n_1394),
.C(n_14),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_2581),
.B(n_1394),
.Y(n_3095)
);

CKINVDCx16_ASAP7_75t_R g3096 ( 
.A(n_2580),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2262),
.B(n_1394),
.Y(n_3097)
);

BUFx2_ASAP7_75t_L g3098 ( 
.A(n_2580),
.Y(n_3098)
);

NAND2xp33_ASAP7_75t_L g3099 ( 
.A(n_2426),
.B(n_1394),
.Y(n_3099)
);

INVxp67_ASAP7_75t_L g3100 ( 
.A(n_2428),
.Y(n_3100)
);

NOR2x1p5_ASAP7_75t_L g3101 ( 
.A(n_2390),
.B(n_12),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_2257),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2260),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2262),
.B(n_1456),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2581),
.B(n_15),
.Y(n_3105)
);

BUFx2_ASAP7_75t_L g3106 ( 
.A(n_2580),
.Y(n_3106)
);

INVx2_ASAP7_75t_SL g3107 ( 
.A(n_2595),
.Y(n_3107)
);

AOI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_2445),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_3108)
);

AND2x2_ASAP7_75t_L g3109 ( 
.A(n_2581),
.B(n_17),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2262),
.B(n_18),
.Y(n_3110)
);

INVx3_ASAP7_75t_L g3111 ( 
.A(n_2540),
.Y(n_3111)
);

NOR2x1p5_ASAP7_75t_L g3112 ( 
.A(n_2390),
.B(n_18),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2257),
.Y(n_3113)
);

OR2x2_ASAP7_75t_L g3114 ( 
.A(n_2324),
.B(n_20),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2262),
.B(n_20),
.Y(n_3115)
);

CKINVDCx5p33_ASAP7_75t_R g3116 ( 
.A(n_2580),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2260),
.Y(n_3117)
);

CKINVDCx14_ASAP7_75t_R g3118 ( 
.A(n_2580),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2262),
.B(n_21),
.Y(n_3119)
);

INVx3_ASAP7_75t_L g3120 ( 
.A(n_2540),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2257),
.Y(n_3121)
);

CKINVDCx5p33_ASAP7_75t_R g3122 ( 
.A(n_2580),
.Y(n_3122)
);

OAI22xp33_ASAP7_75t_L g3123 ( 
.A1(n_2303),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_2257),
.Y(n_3124)
);

INVxp67_ASAP7_75t_L g3125 ( 
.A(n_2428),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2260),
.Y(n_3126)
);

HB1xp67_ASAP7_75t_L g3127 ( 
.A(n_2287),
.Y(n_3127)
);

AOI22xp5_ASAP7_75t_L g3128 ( 
.A1(n_2445),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2257),
.Y(n_3129)
);

BUFx2_ASAP7_75t_L g3130 ( 
.A(n_2580),
.Y(n_3130)
);

BUFx2_ASAP7_75t_L g3131 ( 
.A(n_2580),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2257),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2260),
.Y(n_3133)
);

NAND3xp33_ASAP7_75t_L g3134 ( 
.A(n_2328),
.B(n_23),
.C(n_24),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2260),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2262),
.B(n_25),
.Y(n_3136)
);

CKINVDCx5p33_ASAP7_75t_R g3137 ( 
.A(n_2580),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2260),
.Y(n_3138)
);

AOI22xp33_ASAP7_75t_L g3139 ( 
.A1(n_2526),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2260),
.Y(n_3140)
);

AND2x4_ASAP7_75t_L g3141 ( 
.A(n_2540),
.B(n_25),
.Y(n_3141)
);

INVx3_ASAP7_75t_L g3142 ( 
.A(n_2540),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2257),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2260),
.Y(n_3144)
);

BUFx6f_ASAP7_75t_L g3145 ( 
.A(n_2307),
.Y(n_3145)
);

AOI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_2445),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2260),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2260),
.Y(n_3148)
);

HB1xp67_ASAP7_75t_L g3149 ( 
.A(n_2287),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2257),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2262),
.B(n_26),
.Y(n_3151)
);

NOR2xp33_ASAP7_75t_L g3152 ( 
.A(n_2462),
.B(n_28),
.Y(n_3152)
);

AOI22xp5_ASAP7_75t_L g3153 ( 
.A1(n_2445),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_3153)
);

AND2x4_ASAP7_75t_L g3154 ( 
.A(n_2540),
.B(n_29),
.Y(n_3154)
);

NOR2xp33_ASAP7_75t_L g3155 ( 
.A(n_2462),
.B(n_31),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2257),
.Y(n_3156)
);

AND2x4_ASAP7_75t_L g3157 ( 
.A(n_2540),
.B(n_32),
.Y(n_3157)
);

AND2x2_ASAP7_75t_L g3158 ( 
.A(n_2581),
.B(n_33),
.Y(n_3158)
);

NAND3xp33_ASAP7_75t_L g3159 ( 
.A(n_2328),
.B(n_33),
.C(n_34),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2257),
.Y(n_3160)
);

AO22x2_ASAP7_75t_L g3161 ( 
.A1(n_2324),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2257),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2260),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2260),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_2581),
.B(n_34),
.Y(n_3165)
);

HB1xp67_ASAP7_75t_L g3166 ( 
.A(n_2287),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2257),
.Y(n_3167)
);

OAI22xp5_ASAP7_75t_L g3168 ( 
.A1(n_2482),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_SL g3169 ( 
.A(n_2540),
.B(n_39),
.Y(n_3169)
);

AND2x2_ASAP7_75t_L g3170 ( 
.A(n_2581),
.B(n_38),
.Y(n_3170)
);

AO22x2_ASAP7_75t_L g3171 ( 
.A1(n_2324),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_3171)
);

INVxp67_ASAP7_75t_L g3172 ( 
.A(n_2428),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2257),
.Y(n_3173)
);

AO22x2_ASAP7_75t_L g3174 ( 
.A1(n_2324),
.A2(n_42),
.B1(n_39),
.B2(n_40),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2262),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2262),
.B(n_40),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2262),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_L g3178 ( 
.A(n_2619),
.B(n_42),
.Y(n_3178)
);

AOI21x1_ASAP7_75t_L g3179 ( 
.A1(n_2720),
.A2(n_43),
.B(n_44),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2726),
.B(n_43),
.Y(n_3180)
);

O2A1O1Ixp33_ASAP7_75t_L g3181 ( 
.A1(n_2783),
.A2(n_2743),
.B(n_2727),
.C(n_3040),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_L g3182 ( 
.A(n_2867),
.B(n_43),
.Y(n_3182)
);

AOI22xp33_ASAP7_75t_L g3183 ( 
.A1(n_2908),
.A2(n_2794),
.B1(n_2793),
.B2(n_2929),
.Y(n_3183)
);

AOI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_2762),
.A2(n_44),
.B(n_45),
.Y(n_3184)
);

AOI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_2647),
.A2(n_44),
.B(n_45),
.Y(n_3185)
);

AOI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_2842),
.A2(n_45),
.B(n_46),
.Y(n_3186)
);

INVx2_ASAP7_75t_L g3187 ( 
.A(n_2672),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_2690),
.Y(n_3188)
);

NOR2xp33_ASAP7_75t_SL g3189 ( 
.A(n_3002),
.B(n_2984),
.Y(n_3189)
);

INVx3_ASAP7_75t_L g3190 ( 
.A(n_2984),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2610),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2611),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_SL g3193 ( 
.A(n_2808),
.B(n_724),
.Y(n_3193)
);

INVx2_ASAP7_75t_SL g3194 ( 
.A(n_3079),
.Y(n_3194)
);

INVx2_ASAP7_75t_SL g3195 ( 
.A(n_3079),
.Y(n_3195)
);

AOI21xp5_ASAP7_75t_L g3196 ( 
.A1(n_2717),
.A2(n_47),
.B(n_48),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_2678),
.B(n_49),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2616),
.Y(n_3198)
);

AOI21xp5_ASAP7_75t_L g3199 ( 
.A1(n_2721),
.A2(n_49),
.B(n_50),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2639),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2734),
.A2(n_2739),
.B(n_2736),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2618),
.Y(n_3202)
);

AOI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_2741),
.A2(n_50),
.B(n_51),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2719),
.B(n_51),
.Y(n_3204)
);

A2O1A1Ixp33_ASAP7_75t_L g3205 ( 
.A1(n_3043),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_3205)
);

AOI21xp33_ASAP7_75t_L g3206 ( 
.A1(n_2830),
.A2(n_53),
.B(n_54),
.Y(n_3206)
);

INVx4_ASAP7_75t_L g3207 ( 
.A(n_2644),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2643),
.Y(n_3208)
);

AOI22xp33_ASAP7_75t_L g3209 ( 
.A1(n_2908),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_3209)
);

OAI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_2664),
.A2(n_55),
.B(n_56),
.Y(n_3210)
);

NOR2xp67_ASAP7_75t_L g3211 ( 
.A(n_2644),
.B(n_2698),
.Y(n_3211)
);

O2A1O1Ixp33_ASAP7_75t_SL g3212 ( 
.A1(n_3094),
.A2(n_58),
.B(n_55),
.C(n_57),
.Y(n_3212)
);

O2A1O1Ixp5_ASAP7_75t_L g3213 ( 
.A1(n_2661),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_3213)
);

AOI21x1_ASAP7_75t_L g3214 ( 
.A1(n_2744),
.A2(n_2752),
.B(n_2733),
.Y(n_3214)
);

OAI321xp33_ASAP7_75t_L g3215 ( 
.A1(n_3065),
.A2(n_63),
.A3(n_65),
.B1(n_61),
.B2(n_62),
.C(n_64),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_L g3216 ( 
.A(n_2715),
.B(n_62),
.Y(n_3216)
);

AND2x4_ASAP7_75t_L g3217 ( 
.A(n_2630),
.B(n_62),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2621),
.B(n_63),
.Y(n_3218)
);

HB1xp67_ASAP7_75t_L g3219 ( 
.A(n_2709),
.Y(n_3219)
);

OR2x6_ASAP7_75t_L g3220 ( 
.A(n_2687),
.B(n_64),
.Y(n_3220)
);

AOI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_2671),
.A2(n_64),
.B(n_65),
.Y(n_3221)
);

AOI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_3032),
.A2(n_65),
.B(n_66),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2655),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_2621),
.B(n_66),
.Y(n_3224)
);

AOI21xp5_ASAP7_75t_L g3225 ( 
.A1(n_3056),
.A2(n_67),
.B(n_68),
.Y(n_3225)
);

NAND2x1p5_ASAP7_75t_L g3226 ( 
.A(n_2644),
.B(n_68),
.Y(n_3226)
);

BUFx12f_ASAP7_75t_L g3227 ( 
.A(n_2835),
.Y(n_3227)
);

NOR2xp33_ASAP7_75t_L g3228 ( 
.A(n_2906),
.B(n_68),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_2623),
.B(n_70),
.Y(n_3229)
);

NOR2xp33_ASAP7_75t_L g3230 ( 
.A(n_3000),
.B(n_70),
.Y(n_3230)
);

INVx1_ASAP7_75t_SL g3231 ( 
.A(n_2712),
.Y(n_3231)
);

OAI21xp5_ASAP7_75t_L g3232 ( 
.A1(n_2831),
.A2(n_71),
.B(n_72),
.Y(n_3232)
);

NOR2xp33_ASAP7_75t_L g3233 ( 
.A(n_3013),
.B(n_3019),
.Y(n_3233)
);

A2O1A1Ixp33_ASAP7_75t_L g3234 ( 
.A1(n_3152),
.A2(n_74),
.B(n_71),
.C(n_73),
.Y(n_3234)
);

NAND2xp33_ASAP7_75t_R g3235 ( 
.A(n_2730),
.B(n_73),
.Y(n_3235)
);

AOI21xp5_ASAP7_75t_L g3236 ( 
.A1(n_3062),
.A2(n_73),
.B(n_74),
.Y(n_3236)
);

OAI21xp33_ASAP7_75t_L g3237 ( 
.A1(n_3039),
.A2(n_75),
.B(n_76),
.Y(n_3237)
);

BUFx2_ASAP7_75t_L g3238 ( 
.A(n_2674),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_2945),
.A2(n_75),
.B(n_77),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_2623),
.B(n_77),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_2624),
.B(n_77),
.Y(n_3241)
);

AOI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_3097),
.A2(n_78),
.B(n_79),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_3020),
.B(n_78),
.Y(n_3243)
);

AO21x1_ASAP7_75t_L g3244 ( 
.A1(n_3123),
.A2(n_726),
.B(n_725),
.Y(n_3244)
);

NOR2xp33_ASAP7_75t_L g3245 ( 
.A(n_3021),
.B(n_78),
.Y(n_3245)
);

BUFx6f_ASAP7_75t_L g3246 ( 
.A(n_2659),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2624),
.B(n_2625),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_2625),
.B(n_79),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2626),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_2981),
.B(n_80),
.Y(n_3250)
);

AOI21xp5_ASAP7_75t_L g3251 ( 
.A1(n_3104),
.A2(n_80),
.B(n_81),
.Y(n_3251)
);

CKINVDCx5p33_ASAP7_75t_R g3252 ( 
.A(n_2835),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_2981),
.B(n_81),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2987),
.B(n_82),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_2987),
.B(n_82),
.Y(n_3255)
);

INVxp67_ASAP7_75t_L g3256 ( 
.A(n_2729),
.Y(n_3256)
);

OAI21xp5_ASAP7_75t_L g3257 ( 
.A1(n_2667),
.A2(n_82),
.B(n_83),
.Y(n_3257)
);

NAND2x1p5_ASAP7_75t_L g3258 ( 
.A(n_2786),
.B(n_83),
.Y(n_3258)
);

AOI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_2731),
.A2(n_83),
.B(n_84),
.Y(n_3259)
);

AOI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_3099),
.A2(n_84),
.B(n_85),
.Y(n_3260)
);

OAI21xp5_ASAP7_75t_L g3261 ( 
.A1(n_2685),
.A2(n_84),
.B(n_85),
.Y(n_3261)
);

A2O1A1Ixp33_ASAP7_75t_L g3262 ( 
.A1(n_3155),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_3262)
);

NAND3xp33_ASAP7_75t_L g3263 ( 
.A(n_3134),
.B(n_86),
.C(n_87),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2988),
.B(n_86),
.Y(n_3264)
);

OA22x2_ASAP7_75t_L g3265 ( 
.A1(n_2861),
.A2(n_90),
.B1(n_87),
.B2(n_88),
.Y(n_3265)
);

AND2x4_ASAP7_75t_L g3266 ( 
.A(n_3025),
.B(n_88),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_SL g3267 ( 
.A(n_2753),
.B(n_726),
.Y(n_3267)
);

OAI22xp5_ASAP7_75t_L g3268 ( 
.A1(n_2747),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_3268)
);

BUFx3_ASAP7_75t_L g3269 ( 
.A(n_3041),
.Y(n_3269)
);

HB1xp67_ASAP7_75t_L g3270 ( 
.A(n_2933),
.Y(n_3270)
);

OAI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_2952),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_3271)
);

INVx3_ASAP7_75t_L g3272 ( 
.A(n_2888),
.Y(n_3272)
);

O2A1O1Ixp33_ASAP7_75t_L g3273 ( 
.A1(n_2748),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_3273)
);

OAI22xp5_ASAP7_75t_L g3274 ( 
.A1(n_2952),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2666),
.Y(n_3275)
);

OAI22xp33_ASAP7_75t_L g3276 ( 
.A1(n_3114),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_3276)
);

CKINVDCx8_ASAP7_75t_R g3277 ( 
.A(n_3096),
.Y(n_3277)
);

AOI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_2662),
.A2(n_96),
.B(n_97),
.Y(n_3278)
);

NAND3xp33_ASAP7_75t_L g3279 ( 
.A(n_3159),
.B(n_96),
.C(n_97),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_2988),
.B(n_98),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2991),
.B(n_98),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_2716),
.A2(n_99),
.B(n_100),
.Y(n_3282)
);

OAI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_2969),
.A2(n_99),
.B(n_101),
.Y(n_3283)
);

AND2x4_ASAP7_75t_L g3284 ( 
.A(n_2858),
.B(n_101),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_2678),
.B(n_101),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_SL g3286 ( 
.A(n_3031),
.B(n_727),
.Y(n_3286)
);

NOR2x1_ASAP7_75t_L g3287 ( 
.A(n_2881),
.B(n_102),
.Y(n_3287)
);

AOI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_2854),
.A2(n_102),
.B(n_103),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_L g3289 ( 
.A(n_3042),
.B(n_103),
.Y(n_3289)
);

AO21x1_ASAP7_75t_L g3290 ( 
.A1(n_3168),
.A2(n_728),
.B(n_727),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_2991),
.B(n_103),
.Y(n_3291)
);

AND2x4_ASAP7_75t_L g3292 ( 
.A(n_2858),
.B(n_104),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3067),
.B(n_104),
.Y(n_3293)
);

AND2x4_ASAP7_75t_L g3294 ( 
.A(n_2904),
.B(n_105),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_2613),
.B(n_105),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2669),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_2864),
.A2(n_106),
.B(n_107),
.Y(n_3297)
);

NOR2xp33_ASAP7_75t_L g3298 ( 
.A(n_3100),
.B(n_106),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3067),
.B(n_107),
.Y(n_3299)
);

BUFx8_ASAP7_75t_L g3300 ( 
.A(n_3018),
.Y(n_3300)
);

AOI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_2871),
.A2(n_108),
.B(n_109),
.Y(n_3301)
);

AO32x2_ASAP7_75t_L g3302 ( 
.A1(n_2732),
.A2(n_2909),
.A3(n_2615),
.B1(n_2663),
.B2(n_3026),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_2972),
.A2(n_110),
.B(n_111),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3068),
.B(n_110),
.Y(n_3304)
);

AOI22x1_ASAP7_75t_L g3305 ( 
.A1(n_2637),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_3305)
);

AOI22xp5_ASAP7_75t_L g3306 ( 
.A1(n_3172),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_3306)
);

BUFx6f_ASAP7_75t_L g3307 ( 
.A(n_2659),
.Y(n_3307)
);

OAI22xp5_ASAP7_75t_L g3308 ( 
.A1(n_3125),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_3308)
);

BUFx8_ASAP7_75t_L g3309 ( 
.A(n_3060),
.Y(n_3309)
);

OAI21x1_ASAP7_75t_L g3310 ( 
.A1(n_2968),
.A2(n_115),
.B(n_116),
.Y(n_3310)
);

O2A1O1Ixp33_ASAP7_75t_L g3311 ( 
.A1(n_3047),
.A2(n_118),
.B(n_115),
.C(n_117),
.Y(n_3311)
);

AOI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_2974),
.A2(n_117),
.B(n_118),
.Y(n_3312)
);

NOR2xp33_ASAP7_75t_L g3313 ( 
.A(n_2645),
.B(n_117),
.Y(n_3313)
);

INVxp67_ASAP7_75t_L g3314 ( 
.A(n_2650),
.Y(n_3314)
);

OR2x2_ASAP7_75t_L g3315 ( 
.A(n_2658),
.B(n_118),
.Y(n_3315)
);

O2A1O1Ixp33_ASAP7_75t_L g3316 ( 
.A1(n_3169),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_3316)
);

NOR3xp33_ASAP7_75t_L g3317 ( 
.A(n_2628),
.B(n_119),
.C(n_120),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3068),
.B(n_119),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_2636),
.A2(n_120),
.B(n_122),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_2670),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_2632),
.B(n_122),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3175),
.B(n_123),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3175),
.B(n_123),
.Y(n_3323)
);

INVx2_ASAP7_75t_SL g3324 ( 
.A(n_2888),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_2648),
.A2(n_2652),
.B(n_2651),
.Y(n_3325)
);

AOI21xp5_ASAP7_75t_L g3326 ( 
.A1(n_2656),
.A2(n_123),
.B(n_124),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_2978),
.A2(n_124),
.B(n_125),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_2979),
.A2(n_124),
.B(n_125),
.Y(n_3328)
);

AOI21xp5_ASAP7_75t_L g3329 ( 
.A1(n_2985),
.A2(n_126),
.B(n_127),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_SL g3330 ( 
.A(n_2818),
.B(n_728),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3177),
.B(n_127),
.Y(n_3331)
);

AO21x1_ASAP7_75t_L g3332 ( 
.A1(n_2735),
.A2(n_732),
.B(n_731),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3177),
.B(n_128),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_2989),
.A2(n_128),
.B(n_129),
.Y(n_3334)
);

AOI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_2993),
.A2(n_129),
.B(n_130),
.Y(n_3335)
);

O2A1O1Ixp33_ASAP7_75t_L g3336 ( 
.A1(n_2710),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_3336)
);

A2O1A1Ixp33_ASAP7_75t_L g3337 ( 
.A1(n_3108),
.A2(n_3146),
.B(n_3153),
.C(n_3128),
.Y(n_3337)
);

AND2x4_ASAP7_75t_L g3338 ( 
.A(n_2904),
.B(n_131),
.Y(n_3338)
);

NOR3xp33_ASAP7_75t_L g3339 ( 
.A(n_2966),
.B(n_132),
.C(n_133),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_L g3340 ( 
.A(n_2877),
.B(n_2827),
.Y(n_3340)
);

OAI22xp5_ASAP7_75t_L g3341 ( 
.A1(n_3009),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_3341)
);

OAI22xp5_ASAP7_75t_L g3342 ( 
.A1(n_3022),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_3342)
);

NOR2xp33_ASAP7_75t_L g3343 ( 
.A(n_2673),
.B(n_134),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_3005),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3010),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_2995),
.B(n_137),
.Y(n_3346)
);

INVx2_ASAP7_75t_L g3347 ( 
.A(n_3012),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_SL g3348 ( 
.A(n_2818),
.B(n_731),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_3015),
.Y(n_3349)
);

NOR2xp33_ASAP7_75t_L g3350 ( 
.A(n_2894),
.B(n_139),
.Y(n_3350)
);

AND2x4_ASAP7_75t_L g3351 ( 
.A(n_3044),
.B(n_139),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_SL g3352 ( 
.A(n_2818),
.B(n_732),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_SL g3353 ( 
.A(n_2789),
.B(n_733),
.Y(n_3353)
);

O2A1O1Ixp5_ASAP7_75t_L g3354 ( 
.A1(n_2738),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_3354)
);

NOR3xp33_ASAP7_75t_L g3355 ( 
.A(n_2694),
.B(n_140),
.C(n_141),
.Y(n_3355)
);

INVx2_ASAP7_75t_L g3356 ( 
.A(n_3035),
.Y(n_3356)
);

INVx4_ASAP7_75t_L g3357 ( 
.A(n_2614),
.Y(n_3357)
);

O2A1O1Ixp33_ASAP7_75t_L g3358 ( 
.A1(n_2912),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_3358)
);

AOI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_3037),
.A2(n_143),
.B(n_144),
.Y(n_3359)
);

AOI21xp5_ASAP7_75t_L g3360 ( 
.A1(n_3046),
.A2(n_3084),
.B(n_3083),
.Y(n_3360)
);

NOR2x1_ASAP7_75t_L g3361 ( 
.A(n_2706),
.B(n_145),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_2997),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_SL g3363 ( 
.A(n_2829),
.B(n_2722),
.Y(n_3363)
);

AOI21xp5_ASAP7_75t_L g3364 ( 
.A1(n_3093),
.A2(n_145),
.B(n_146),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_2999),
.B(n_146),
.Y(n_3365)
);

AOI21xp5_ASAP7_75t_L g3366 ( 
.A1(n_3102),
.A2(n_147),
.B(n_148),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3001),
.B(n_148),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3008),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_2836),
.B(n_149),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_L g3370 ( 
.A(n_3091),
.B(n_149),
.Y(n_3370)
);

O2A1O1Ixp5_ASAP7_75t_L g3371 ( 
.A1(n_2742),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_2749),
.B(n_150),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3028),
.B(n_152),
.Y(n_3373)
);

NAND2x1p5_ASAP7_75t_L g3374 ( 
.A(n_2706),
.B(n_152),
.Y(n_3374)
);

AO21x2_ASAP7_75t_L g3375 ( 
.A1(n_2745),
.A2(n_153),
.B(n_154),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3029),
.Y(n_3376)
);

AOI21xp5_ASAP7_75t_L g3377 ( 
.A1(n_3113),
.A2(n_155),
.B(n_156),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3036),
.B(n_155),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3048),
.B(n_156),
.Y(n_3379)
);

AOI22xp5_ASAP7_75t_L g3380 ( 
.A1(n_3030),
.A2(n_2646),
.B1(n_2755),
.B2(n_2737),
.Y(n_3380)
);

OAI21xp5_ASAP7_75t_L g3381 ( 
.A1(n_3110),
.A2(n_3119),
.B(n_3115),
.Y(n_3381)
);

OAI22xp5_ASAP7_75t_L g3382 ( 
.A1(n_2681),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_3382)
);

NOR2xp33_ASAP7_75t_L g3383 ( 
.A(n_2680),
.B(n_157),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3052),
.Y(n_3384)
);

AOI21xp5_ASAP7_75t_L g3385 ( 
.A1(n_3121),
.A2(n_159),
.B(n_160),
.Y(n_3385)
);

OAI22xp5_ASAP7_75t_L g3386 ( 
.A1(n_2681),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_3386)
);

AOI21xp5_ASAP7_75t_L g3387 ( 
.A1(n_3124),
.A2(n_161),
.B(n_162),
.Y(n_3387)
);

NOR2xp33_ASAP7_75t_L g3388 ( 
.A(n_2880),
.B(n_164),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_3129),
.Y(n_3389)
);

INVx11_ASAP7_75t_L g3390 ( 
.A(n_2897),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_SL g3391 ( 
.A(n_2701),
.B(n_734),
.Y(n_3391)
);

BUFx2_ASAP7_75t_L g3392 ( 
.A(n_2701),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_SL g3393 ( 
.A(n_2898),
.B(n_736),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3054),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3055),
.Y(n_3395)
);

AOI21x1_ASAP7_75t_L g3396 ( 
.A1(n_2746),
.A2(n_165),
.B(n_166),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3059),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3061),
.B(n_166),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3074),
.B(n_166),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3078),
.B(n_167),
.Y(n_3400)
);

OAI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_3136),
.A2(n_168),
.B(n_169),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3132),
.A2(n_169),
.B(n_170),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_3143),
.A2(n_170),
.B(n_171),
.Y(n_3403)
);

A2O1A1Ixp33_ASAP7_75t_L g3404 ( 
.A1(n_3151),
.A2(n_174),
.B(n_172),
.C(n_173),
.Y(n_3404)
);

A2O1A1Ixp33_ASAP7_75t_L g3405 ( 
.A1(n_3176),
.A2(n_175),
.B(n_172),
.C(n_173),
.Y(n_3405)
);

AOI21xp5_ASAP7_75t_L g3406 ( 
.A1(n_3150),
.A2(n_3173),
.B(n_3167),
.Y(n_3406)
);

BUFx6f_ASAP7_75t_L g3407 ( 
.A(n_2659),
.Y(n_3407)
);

AOI21xp5_ASAP7_75t_L g3408 ( 
.A1(n_3156),
.A2(n_175),
.B(n_176),
.Y(n_3408)
);

AOI21xp5_ASAP7_75t_L g3409 ( 
.A1(n_3160),
.A2(n_176),
.B(n_177),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3080),
.B(n_177),
.Y(n_3410)
);

NOR2xp33_ASAP7_75t_L g3411 ( 
.A(n_2689),
.B(n_178),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3081),
.Y(n_3412)
);

NOR2xp33_ASAP7_75t_L g3413 ( 
.A(n_2924),
.B(n_178),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3085),
.B(n_3086),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_SL g3415 ( 
.A(n_2898),
.B(n_736),
.Y(n_3415)
);

INVx5_ASAP7_75t_L g3416 ( 
.A(n_2614),
.Y(n_3416)
);

A2O1A1Ixp33_ASAP7_75t_L g3417 ( 
.A1(n_2631),
.A2(n_182),
.B(n_179),
.C(n_181),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_SL g3418 ( 
.A(n_2898),
.B(n_737),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3087),
.B(n_181),
.Y(n_3419)
);

AOI33xp33_ASAP7_75t_L g3420 ( 
.A1(n_2718),
.A2(n_184),
.A3(n_186),
.B1(n_182),
.B2(n_183),
.B3(n_185),
.Y(n_3420)
);

BUFx6f_ASAP7_75t_L g3421 ( 
.A(n_2707),
.Y(n_3421)
);

O2A1O1Ixp5_ASAP7_75t_L g3422 ( 
.A1(n_2758),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_SL g3423 ( 
.A(n_2937),
.B(n_738),
.Y(n_3423)
);

OAI21xp5_ASAP7_75t_L g3424 ( 
.A1(n_2609),
.A2(n_184),
.B(n_185),
.Y(n_3424)
);

O2A1O1Ixp33_ASAP7_75t_L g3425 ( 
.A1(n_2772),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3088),
.B(n_186),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3090),
.Y(n_3427)
);

INVxp67_ASAP7_75t_L g3428 ( 
.A(n_2650),
.Y(n_3428)
);

AOI22xp5_ASAP7_75t_L g3429 ( 
.A1(n_2919),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_3429)
);

AOI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_3162),
.A2(n_190),
.B(n_191),
.Y(n_3430)
);

INVx1_ASAP7_75t_SL g3431 ( 
.A(n_3098),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3092),
.B(n_191),
.Y(n_3432)
);

OR2x2_ASAP7_75t_L g3433 ( 
.A(n_2657),
.B(n_191),
.Y(n_3433)
);

A2O1A1Ixp33_ASAP7_75t_L g3434 ( 
.A1(n_2634),
.A2(n_194),
.B(n_192),
.C(n_193),
.Y(n_3434)
);

OAI21xp5_ASAP7_75t_L g3435 ( 
.A1(n_2612),
.A2(n_192),
.B(n_193),
.Y(n_3435)
);

OAI22xp5_ASAP7_75t_L g3436 ( 
.A1(n_3082),
.A2(n_2821),
.B1(n_3011),
.B2(n_2986),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_2634),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3103),
.B(n_192),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_3117),
.B(n_194),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3126),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_2976),
.B(n_195),
.Y(n_3441)
);

INVx2_ASAP7_75t_SL g3442 ( 
.A(n_2866),
.Y(n_3442)
);

OAI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_3051),
.A2(n_195),
.B(n_196),
.Y(n_3443)
);

OAI22xp5_ASAP7_75t_L g3444 ( 
.A1(n_2821),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_2635),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_2693),
.B(n_197),
.Y(n_3446)
);

AOI21xp5_ASAP7_75t_L g3447 ( 
.A1(n_2697),
.A2(n_197),
.B(n_198),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3133),
.B(n_198),
.Y(n_3448)
);

AOI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_2700),
.A2(n_199),
.B(n_200),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3135),
.Y(n_3450)
);

AOI21xp5_ASAP7_75t_L g3451 ( 
.A1(n_2702),
.A2(n_199),
.B(n_200),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3138),
.B(n_201),
.Y(n_3452)
);

A2O1A1Ixp33_ASAP7_75t_L g3453 ( 
.A1(n_2635),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_2840),
.A2(n_202),
.B(n_203),
.Y(n_3454)
);

A2O1A1Ixp33_ASAP7_75t_L g3455 ( 
.A1(n_2638),
.A2(n_205),
.B(n_202),
.C(n_204),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_2638),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3140),
.B(n_204),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_2691),
.Y(n_3458)
);

AND2x2_ASAP7_75t_L g3459 ( 
.A(n_2977),
.B(n_206),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3144),
.B(n_207),
.Y(n_3460)
);

NOR2xp33_ASAP7_75t_L g3461 ( 
.A(n_2834),
.B(n_207),
.Y(n_3461)
);

INVxp67_ASAP7_75t_L g3462 ( 
.A(n_3069),
.Y(n_3462)
);

AOI21xp5_ASAP7_75t_L g3463 ( 
.A1(n_2841),
.A2(n_208),
.B(n_209),
.Y(n_3463)
);

AOI21xp5_ASAP7_75t_L g3464 ( 
.A1(n_2800),
.A2(n_208),
.B(n_209),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3147),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3148),
.B(n_208),
.Y(n_3466)
);

O2A1O1Ixp33_ASAP7_75t_L g3467 ( 
.A1(n_2891),
.A2(n_212),
.B(n_210),
.C(n_211),
.Y(n_3467)
);

OAI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_3058),
.A2(n_210),
.B(n_211),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_SL g3469 ( 
.A(n_2937),
.B(n_738),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_SL g3470 ( 
.A(n_2937),
.B(n_739),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3163),
.B(n_212),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3164),
.Y(n_3472)
);

AOI21xp5_ASAP7_75t_L g3473 ( 
.A1(n_2800),
.A2(n_2839),
.B(n_2838),
.Y(n_3473)
);

AO21x1_ASAP7_75t_L g3474 ( 
.A1(n_2846),
.A2(n_740),
.B(n_739),
.Y(n_3474)
);

NAND2x1p5_ASAP7_75t_L g3475 ( 
.A(n_2860),
.B(n_213),
.Y(n_3475)
);

AOI21xp5_ASAP7_75t_L g3476 ( 
.A1(n_2838),
.A2(n_213),
.B(n_214),
.Y(n_3476)
);

BUFx6f_ASAP7_75t_L g3477 ( 
.A(n_2707),
.Y(n_3477)
);

OAI21xp5_ASAP7_75t_L g3478 ( 
.A1(n_3072),
.A2(n_213),
.B(n_215),
.Y(n_3478)
);

NAND2x1p5_ASAP7_75t_L g3479 ( 
.A(n_2860),
.B(n_215),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_2759),
.B(n_215),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_L g3481 ( 
.A(n_2851),
.B(n_216),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_L g3482 ( 
.A1(n_2870),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_2761),
.B(n_216),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3105),
.B(n_218),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3109),
.B(n_218),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_2839),
.A2(n_219),
.B(n_220),
.Y(n_3486)
);

AOI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_2707),
.A2(n_220),
.B(n_221),
.Y(n_3487)
);

AOI21xp5_ASAP7_75t_L g3488 ( 
.A1(n_2788),
.A2(n_3145),
.B(n_2812),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_2695),
.Y(n_3489)
);

AOI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_2788),
.A2(n_220),
.B(n_221),
.Y(n_3490)
);

A2O1A1Ixp33_ASAP7_75t_L g3491 ( 
.A1(n_2787),
.A2(n_224),
.B(n_222),
.C(n_223),
.Y(n_3491)
);

NAND2xp33_ASAP7_75t_L g3492 ( 
.A(n_2614),
.B(n_223),
.Y(n_3492)
);

A2O1A1Ixp33_ASAP7_75t_L g3493 ( 
.A1(n_2822),
.A2(n_225),
.B(n_223),
.C(n_224),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3158),
.B(n_225),
.Y(n_3494)
);

AOI22xp33_ASAP7_75t_L g3495 ( 
.A1(n_2870),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_3495)
);

AO32x1_ASAP7_75t_L g3496 ( 
.A1(n_2799),
.A2(n_228),
.A3(n_226),
.B1(n_227),
.B2(n_229),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3165),
.B(n_226),
.Y(n_3497)
);

BUFx6f_ASAP7_75t_L g3498 ( 
.A(n_2788),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_2983),
.B(n_228),
.Y(n_3499)
);

BUFx3_ASAP7_75t_L g3500 ( 
.A(n_2811),
.Y(n_3500)
);

OAI21xp5_ASAP7_75t_L g3501 ( 
.A1(n_3076),
.A2(n_228),
.B(n_229),
.Y(n_3501)
);

OA22x2_ASAP7_75t_L g3502 ( 
.A1(n_3050),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3170),
.B(n_230),
.Y(n_3503)
);

AOI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_2812),
.A2(n_230),
.B(n_231),
.Y(n_3504)
);

AOI33xp33_ASAP7_75t_L g3505 ( 
.A1(n_2642),
.A2(n_233),
.A3(n_235),
.B1(n_231),
.B2(n_232),
.B3(n_234),
.Y(n_3505)
);

AOI21x1_ASAP7_75t_L g3506 ( 
.A1(n_2801),
.A2(n_232),
.B(n_233),
.Y(n_3506)
);

BUFx3_ASAP7_75t_L g3507 ( 
.A(n_2897),
.Y(n_3507)
);

OAI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_2986),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_2812),
.A2(n_235),
.B(n_236),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_2996),
.B(n_236),
.Y(n_3510)
);

A2O1A1Ixp33_ASAP7_75t_L g3511 ( 
.A1(n_2872),
.A2(n_239),
.B(n_237),
.C(n_238),
.Y(n_3511)
);

NOR2xp33_ASAP7_75t_L g3512 ( 
.A(n_3106),
.B(n_238),
.Y(n_3512)
);

NOR2xp33_ASAP7_75t_L g3513 ( 
.A(n_3130),
.B(n_238),
.Y(n_3513)
);

INVxp67_ASAP7_75t_L g3514 ( 
.A(n_3116),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_2676),
.B(n_239),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_SL g3516 ( 
.A(n_2961),
.B(n_740),
.Y(n_3516)
);

OR2x2_ASAP7_75t_L g3517 ( 
.A(n_3038),
.B(n_240),
.Y(n_3517)
);

NAND2xp33_ASAP7_75t_L g3518 ( 
.A(n_2614),
.B(n_241),
.Y(n_3518)
);

O2A1O1Ixp33_ASAP7_75t_L g3519 ( 
.A1(n_2820),
.A2(n_244),
.B(n_242),
.C(n_243),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_2682),
.B(n_2683),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_2684),
.B(n_242),
.Y(n_3521)
);

BUFx4f_ASAP7_75t_L g3522 ( 
.A(n_3045),
.Y(n_3522)
);

AOI21xp5_ASAP7_75t_L g3523 ( 
.A1(n_2708),
.A2(n_243),
.B(n_244),
.Y(n_3523)
);

INVxp67_ASAP7_75t_SL g3524 ( 
.A(n_2917),
.Y(n_3524)
);

AOI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_2826),
.A2(n_244),
.B(n_245),
.Y(n_3525)
);

AOI21xp5_ASAP7_75t_L g3526 ( 
.A1(n_2828),
.A2(n_246),
.B(n_247),
.Y(n_3526)
);

OAI22xp5_ASAP7_75t_L g3527 ( 
.A1(n_3011),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_3527)
);

BUFx8_ASAP7_75t_L g3528 ( 
.A(n_3131),
.Y(n_3528)
);

AOI21x1_ASAP7_75t_L g3529 ( 
.A1(n_2926),
.A2(n_246),
.B(n_248),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_2686),
.B(n_248),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_2832),
.A2(n_249),
.B(n_250),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_2688),
.B(n_250),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_2696),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_2852),
.B(n_250),
.Y(n_3534)
);

NOR2xp33_ASAP7_75t_L g3535 ( 
.A(n_2936),
.B(n_251),
.Y(n_3535)
);

AND2x4_ASAP7_75t_L g3536 ( 
.A(n_3044),
.B(n_251),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_2703),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_2692),
.B(n_251),
.Y(n_3538)
);

NOR2xp33_ASAP7_75t_L g3539 ( 
.A(n_2875),
.B(n_2668),
.Y(n_3539)
);

NOR3xp33_ASAP7_75t_L g3540 ( 
.A(n_2948),
.B(n_252),
.C(n_253),
.Y(n_3540)
);

NOR2xp33_ASAP7_75t_L g3541 ( 
.A(n_2792),
.B(n_252),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_2704),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_2705),
.Y(n_3543)
);

OAI22xp5_ASAP7_75t_L g3544 ( 
.A1(n_3016),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_3544)
);

BUFx3_ASAP7_75t_L g3545 ( 
.A(n_2714),
.Y(n_3545)
);

AOI21xp5_ASAP7_75t_L g3546 ( 
.A1(n_2824),
.A2(n_256),
.B(n_257),
.Y(n_3546)
);

NOR2xp33_ASAP7_75t_L g3547 ( 
.A(n_2819),
.B(n_256),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_2903),
.B(n_257),
.Y(n_3548)
);

AOI22xp33_ASAP7_75t_L g3549 ( 
.A1(n_3016),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_3549)
);

INVx3_ASAP7_75t_L g3550 ( 
.A(n_3063),
.Y(n_3550)
);

NOR2xp33_ASAP7_75t_SL g3551 ( 
.A(n_3122),
.B(n_259),
.Y(n_3551)
);

INVx2_ASAP7_75t_SL g3552 ( 
.A(n_3063),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_2711),
.Y(n_3553)
);

AOI22xp5_ASAP7_75t_L g3554 ( 
.A1(n_2770),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_2907),
.B(n_261),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_2763),
.A2(n_261),
.B(n_262),
.Y(n_3556)
);

BUFx6f_ASAP7_75t_L g3557 ( 
.A(n_2961),
.Y(n_3557)
);

BUFx6f_ASAP7_75t_L g3558 ( 
.A(n_2961),
.Y(n_3558)
);

AND2x2_ASAP7_75t_L g3559 ( 
.A(n_2677),
.B(n_262),
.Y(n_3559)
);

AOI22x1_ASAP7_75t_L g3560 ( 
.A1(n_2837),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_3560)
);

AOI22xp5_ASAP7_75t_L g3561 ( 
.A1(n_2675),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_3561)
);

O2A1O1Ixp33_ASAP7_75t_L g3562 ( 
.A1(n_2740),
.A2(n_267),
.B(n_264),
.C(n_266),
.Y(n_3562)
);

AND2x4_ASAP7_75t_L g3563 ( 
.A(n_3111),
.B(n_266),
.Y(n_3563)
);

BUFx6f_ASAP7_75t_L g3564 ( 
.A(n_3111),
.Y(n_3564)
);

NOR2x1_ASAP7_75t_L g3565 ( 
.A(n_3101),
.B(n_267),
.Y(n_3565)
);

OAI21xp5_ASAP7_75t_L g3566 ( 
.A1(n_3095),
.A2(n_2810),
.B(n_2843),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_2713),
.A2(n_267),
.B(n_268),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_2728),
.B(n_2751),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_2816),
.B(n_268),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_2825),
.B(n_269),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_SL g3571 ( 
.A(n_2617),
.B(n_741),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_2814),
.Y(n_3572)
);

AOI21xp5_ASAP7_75t_L g3573 ( 
.A1(n_2815),
.A2(n_2883),
.B(n_2874),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_2890),
.B(n_269),
.Y(n_3574)
);

NOR3xp33_ASAP7_75t_L g3575 ( 
.A(n_3024),
.B(n_270),
.C(n_271),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3070),
.Y(n_3576)
);

NOR2x1_ASAP7_75t_L g3577 ( 
.A(n_3112),
.B(n_3120),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_2798),
.B(n_270),
.Y(n_3578)
);

AND2x6_ASAP7_75t_L g3579 ( 
.A(n_3050),
.B(n_270),
.Y(n_3579)
);

BUFx3_ASAP7_75t_L g3580 ( 
.A(n_2757),
.Y(n_3580)
);

HB1xp67_ASAP7_75t_L g3581 ( 
.A(n_3137),
.Y(n_3581)
);

AOI21xp5_ASAP7_75t_L g3582 ( 
.A1(n_3049),
.A2(n_271),
.B(n_272),
.Y(n_3582)
);

AOI21x1_ASAP7_75t_L g3583 ( 
.A1(n_2927),
.A2(n_2934),
.B(n_2930),
.Y(n_3583)
);

BUFx6f_ASAP7_75t_L g3584 ( 
.A(n_3120),
.Y(n_3584)
);

NAND2xp33_ASAP7_75t_L g3585 ( 
.A(n_2850),
.B(n_273),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3070),
.Y(n_3586)
);

BUFx4f_ASAP7_75t_L g3587 ( 
.A(n_3077),
.Y(n_3587)
);

O2A1O1Ixp5_ASAP7_75t_L g3588 ( 
.A1(n_3057),
.A2(n_275),
.B(n_273),
.C(n_274),
.Y(n_3588)
);

INVx3_ASAP7_75t_L g3589 ( 
.A(n_3142),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_2863),
.B(n_274),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_2853),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_2868),
.B(n_275),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_2886),
.B(n_276),
.Y(n_3593)
);

O2A1O1Ixp33_ASAP7_75t_L g3594 ( 
.A1(n_2884),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_2847),
.A2(n_278),
.B(n_279),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_2784),
.Y(n_3596)
);

AOI21x1_ASAP7_75t_L g3597 ( 
.A1(n_2970),
.A2(n_278),
.B(n_280),
.Y(n_3597)
);

INVxp67_ASAP7_75t_L g3598 ( 
.A(n_2629),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_2760),
.A2(n_280),
.B(n_281),
.Y(n_3599)
);

AOI21xp5_ASAP7_75t_L g3600 ( 
.A1(n_2769),
.A2(n_282),
.B(n_283),
.Y(n_3600)
);

AOI21x1_ASAP7_75t_L g3601 ( 
.A1(n_2970),
.A2(n_283),
.B(n_284),
.Y(n_3601)
);

INVx3_ASAP7_75t_L g3602 ( 
.A(n_3142),
.Y(n_3602)
);

AOI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_2777),
.A2(n_283),
.B(n_284),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_2782),
.A2(n_285),
.B(n_286),
.Y(n_3604)
);

O2A1O1Ixp5_ASAP7_75t_L g3605 ( 
.A1(n_2940),
.A2(n_287),
.B(n_285),
.C(n_286),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3073),
.Y(n_3606)
);

A2O1A1Ixp33_ASAP7_75t_L g3607 ( 
.A1(n_2899),
.A2(n_288),
.B(n_286),
.C(n_287),
.Y(n_3607)
);

AND2x2_ASAP7_75t_SL g3608 ( 
.A(n_3053),
.B(n_288),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_2791),
.A2(n_289),
.B(n_290),
.Y(n_3609)
);

OAI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_2857),
.A2(n_2873),
.B(n_2859),
.Y(n_3610)
);

AOI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_2795),
.A2(n_289),
.B(n_290),
.Y(n_3611)
);

OAI22xp5_ASAP7_75t_L g3612 ( 
.A1(n_2913),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_2923),
.B(n_291),
.Y(n_3613)
);

NOR2xp67_ASAP7_75t_L g3614 ( 
.A(n_2960),
.B(n_292),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_2980),
.B(n_293),
.Y(n_3615)
);

AOI21xp5_ASAP7_75t_L g3616 ( 
.A1(n_2796),
.A2(n_293),
.B(n_294),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_2805),
.A2(n_294),
.B(n_295),
.Y(n_3617)
);

NAND3xp33_ASAP7_75t_L g3618 ( 
.A(n_3139),
.B(n_295),
.C(n_296),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_2785),
.Y(n_3619)
);

NAND2x1p5_ASAP7_75t_L g3620 ( 
.A(n_2998),
.B(n_3033),
.Y(n_3620)
);

A2O1A1Ixp33_ASAP7_75t_L g3621 ( 
.A1(n_2780),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_3621)
);

A2O1A1Ixp33_ASAP7_75t_L g3622 ( 
.A1(n_2627),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_3622)
);

AOI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_2813),
.A2(n_298),
.B(n_299),
.Y(n_3623)
);

INVx2_ASAP7_75t_L g3624 ( 
.A(n_2653),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_2617),
.B(n_742),
.Y(n_3625)
);

NOR2xp33_ASAP7_75t_L g3626 ( 
.A(n_2775),
.B(n_300),
.Y(n_3626)
);

HB1xp67_ASAP7_75t_L g3627 ( 
.A(n_3118),
.Y(n_3627)
);

AOI21xp5_ASAP7_75t_L g3628 ( 
.A1(n_2973),
.A2(n_300),
.B(n_301),
.Y(n_3628)
);

NOR2xp67_ASAP7_75t_L g3629 ( 
.A(n_2750),
.B(n_300),
.Y(n_3629)
);

OAI22xp5_ASAP7_75t_L g3630 ( 
.A1(n_2913),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_3630)
);

AOI21xp5_ASAP7_75t_L g3631 ( 
.A1(n_2994),
.A2(n_302),
.B(n_303),
.Y(n_3631)
);

INVx2_ASAP7_75t_L g3632 ( 
.A(n_2653),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3073),
.Y(n_3633)
);

NAND2x1p5_ASAP7_75t_L g3634 ( 
.A(n_3107),
.B(n_303),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3003),
.B(n_304),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_SL g3636 ( 
.A(n_2640),
.B(n_743),
.Y(n_3636)
);

AOI22xp5_ASAP7_75t_L g3637 ( 
.A1(n_2956),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_3637)
);

AOI21xp5_ASAP7_75t_L g3638 ( 
.A1(n_3006),
.A2(n_304),
.B(n_305),
.Y(n_3638)
);

INVx3_ASAP7_75t_L g3639 ( 
.A(n_2949),
.Y(n_3639)
);

O2A1O1Ixp33_ASAP7_75t_SL g3640 ( 
.A1(n_2967),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_2767),
.Y(n_3641)
);

AND2x2_ASAP7_75t_L g3642 ( 
.A(n_2771),
.B(n_307),
.Y(n_3642)
);

BUFx6f_ASAP7_75t_L g3643 ( 
.A(n_2856),
.Y(n_3643)
);

AOI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_2885),
.A2(n_2900),
.B(n_2896),
.Y(n_3644)
);

AND2x4_ASAP7_75t_L g3645 ( 
.A(n_2918),
.B(n_309),
.Y(n_3645)
);

NAND2x1_ASAP7_75t_L g3646 ( 
.A(n_2767),
.B(n_309),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_2848),
.B(n_310),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_2893),
.B(n_310),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_2804),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_2641),
.B(n_310),
.Y(n_3650)
);

AOI21x1_ASAP7_75t_L g3651 ( 
.A1(n_2946),
.A2(n_311),
.B(n_312),
.Y(n_3651)
);

OAI21x1_ASAP7_75t_L g3652 ( 
.A1(n_2804),
.A2(n_311),
.B(n_312),
.Y(n_3652)
);

OAI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3075),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_3653)
);

HB1xp67_ASAP7_75t_L g3654 ( 
.A(n_3053),
.Y(n_3654)
);

AOI21xp5_ASAP7_75t_L g3655 ( 
.A1(n_2901),
.A2(n_313),
.B(n_314),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_SL g3656 ( 
.A(n_3007),
.B(n_744),
.Y(n_3656)
);

AND2x4_ASAP7_75t_L g3657 ( 
.A(n_2953),
.B(n_313),
.Y(n_3657)
);

OAI22xp5_ASAP7_75t_L g3658 ( 
.A1(n_3075),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_3658)
);

NOR3xp33_ASAP7_75t_L g3659 ( 
.A(n_2941),
.B(n_314),
.C(n_315),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_2641),
.B(n_317),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_2975),
.Y(n_3661)
);

AOI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_2876),
.A2(n_317),
.B(n_318),
.Y(n_3662)
);

AOI21xp5_ASAP7_75t_L g3663 ( 
.A1(n_2878),
.A2(n_318),
.B(n_319),
.Y(n_3663)
);

NAND3xp33_ASAP7_75t_L g3664 ( 
.A(n_2809),
.B(n_2911),
.C(n_2943),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_2649),
.B(n_318),
.Y(n_3665)
);

INVx3_ASAP7_75t_L g3666 ( 
.A(n_2910),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_2649),
.B(n_319),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3178),
.B(n_2902),
.Y(n_3668)
);

A2O1A1Ixp33_ASAP7_75t_L g3669 ( 
.A1(n_3562),
.A2(n_3071),
.B(n_3141),
.C(n_3064),
.Y(n_3669)
);

INVx3_ASAP7_75t_L g3670 ( 
.A(n_3227),
.Y(n_3670)
);

AOI21xp5_ASAP7_75t_L g3671 ( 
.A1(n_3492),
.A2(n_3518),
.B(n_3381),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3201),
.A2(n_2845),
.B(n_2844),
.Y(n_3672)
);

AOI22xp5_ASAP7_75t_L g3673 ( 
.A1(n_3608),
.A2(n_2920),
.B1(n_2925),
.B2(n_3064),
.Y(n_3673)
);

NOR2x1_ASAP7_75t_L g3674 ( 
.A(n_3220),
.B(n_3071),
.Y(n_3674)
);

NOR2xp33_ASAP7_75t_L g3675 ( 
.A(n_3539),
.B(n_2774),
.Y(n_3675)
);

AND2x4_ASAP7_75t_SL g3676 ( 
.A(n_3272),
.B(n_2949),
.Y(n_3676)
);

BUFx6f_ASAP7_75t_L g3677 ( 
.A(n_3500),
.Y(n_3677)
);

NOR2xp33_ASAP7_75t_SL g3678 ( 
.A(n_3189),
.B(n_2905),
.Y(n_3678)
);

OAI22xp5_ASAP7_75t_L g3679 ( 
.A1(n_3436),
.A2(n_3171),
.B1(n_3174),
.B2(n_3161),
.Y(n_3679)
);

OAI22xp5_ASAP7_75t_L g3680 ( 
.A1(n_3314),
.A2(n_3171),
.B1(n_3174),
.B2(n_3161),
.Y(n_3680)
);

BUFx6f_ASAP7_75t_L g3681 ( 
.A(n_3545),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3197),
.B(n_3141),
.Y(n_3682)
);

CKINVDCx20_ASAP7_75t_R g3683 ( 
.A(n_3252),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3187),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3414),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3219),
.B(n_2920),
.Y(n_3686)
);

OR2x2_ASAP7_75t_L g3687 ( 
.A(n_3517),
.B(n_3154),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_SL g3688 ( 
.A(n_3416),
.B(n_3357),
.Y(n_3688)
);

INVx6_ASAP7_75t_L g3689 ( 
.A(n_3300),
.Y(n_3689)
);

OAI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_3428),
.A2(n_2925),
.B1(n_2771),
.B2(n_2803),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3188),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3458),
.Y(n_3692)
);

AOI21xp5_ASAP7_75t_L g3693 ( 
.A1(n_3473),
.A2(n_2849),
.B(n_2916),
.Y(n_3693)
);

HB1xp67_ASAP7_75t_L g3694 ( 
.A(n_3270),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3182),
.B(n_2803),
.Y(n_3695)
);

OAI22xp5_ASAP7_75t_L g3696 ( 
.A1(n_3337),
.A2(n_3089),
.B1(n_3157),
.B2(n_3154),
.Y(n_3696)
);

AOI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_3488),
.A2(n_2922),
.B(n_2921),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3233),
.B(n_2942),
.Y(n_3698)
);

AOI21xp5_ASAP7_75t_L g3699 ( 
.A1(n_3184),
.A2(n_2939),
.B(n_2935),
.Y(n_3699)
);

AOI21xp5_ASAP7_75t_L g3700 ( 
.A1(n_3247),
.A2(n_2954),
.B(n_2951),
.Y(n_3700)
);

INVx5_ASAP7_75t_L g3701 ( 
.A(n_3220),
.Y(n_3701)
);

OAI22xp5_ASAP7_75t_L g3702 ( 
.A1(n_3380),
.A2(n_3157),
.B1(n_2855),
.B2(n_2773),
.Y(n_3702)
);

NOR2xp33_ASAP7_75t_L g3703 ( 
.A(n_3256),
.B(n_2776),
.Y(n_3703)
);

AND2x2_ASAP7_75t_L g3704 ( 
.A(n_3285),
.B(n_3014),
.Y(n_3704)
);

NOR2xp33_ASAP7_75t_L g3705 ( 
.A(n_3431),
.B(n_2802),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3191),
.Y(n_3706)
);

INVx5_ASAP7_75t_L g3707 ( 
.A(n_3357),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3192),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_SL g3709 ( 
.A(n_3416),
.B(n_2982),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3489),
.Y(n_3710)
);

HB1xp67_ASAP7_75t_L g3711 ( 
.A(n_3231),
.Y(n_3711)
);

AOI22xp5_ASAP7_75t_L g3712 ( 
.A1(n_3340),
.A2(n_2665),
.B1(n_2879),
.B2(n_2955),
.Y(n_3712)
);

AND2x4_ASAP7_75t_L g3713 ( 
.A(n_3416),
.B(n_2882),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_3198),
.B(n_2931),
.Y(n_3714)
);

OAI21x1_ASAP7_75t_L g3715 ( 
.A1(n_3214),
.A2(n_2892),
.B(n_2862),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_SL g3716 ( 
.A(n_3577),
.B(n_3004),
.Y(n_3716)
);

OAI22xp5_ASAP7_75t_L g3717 ( 
.A1(n_3183),
.A2(n_2781),
.B1(n_2823),
.B2(n_2817),
.Y(n_3717)
);

AOI21xp5_ASAP7_75t_L g3718 ( 
.A1(n_3325),
.A2(n_2958),
.B(n_2957),
.Y(n_3718)
);

AOI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_3360),
.A2(n_2962),
.B(n_2950),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3406),
.A2(n_2963),
.B(n_2971),
.Y(n_3720)
);

NAND2x1p5_ASAP7_75t_L g3721 ( 
.A(n_3190),
.B(n_2754),
.Y(n_3721)
);

BUFx6f_ASAP7_75t_L g3722 ( 
.A(n_3580),
.Y(n_3722)
);

INVx5_ASAP7_75t_L g3723 ( 
.A(n_3190),
.Y(n_3723)
);

OAI22xp5_ASAP7_75t_L g3724 ( 
.A1(n_3549),
.A2(n_3209),
.B1(n_3495),
.B2(n_3482),
.Y(n_3724)
);

OAI21x1_ASAP7_75t_L g3725 ( 
.A1(n_3583),
.A2(n_2797),
.B(n_2889),
.Y(n_3725)
);

BUFx2_ASAP7_75t_L g3726 ( 
.A(n_3522),
.Y(n_3726)
);

INVx6_ASAP7_75t_L g3727 ( 
.A(n_3300),
.Y(n_3727)
);

AO21x1_ASAP7_75t_L g3728 ( 
.A1(n_3653),
.A2(n_3034),
.B(n_3014),
.Y(n_3728)
);

BUFx6f_ASAP7_75t_L g3729 ( 
.A(n_3269),
.Y(n_3729)
);

AOI22xp33_ASAP7_75t_L g3730 ( 
.A1(n_3339),
.A2(n_2944),
.B1(n_2964),
.B2(n_2879),
.Y(n_3730)
);

OAI22xp5_ASAP7_75t_L g3731 ( 
.A1(n_3565),
.A2(n_3034),
.B1(n_2756),
.B2(n_2779),
.Y(n_3731)
);

OAI22x1_ASAP7_75t_L g3732 ( 
.A1(n_3284),
.A2(n_2654),
.B1(n_2660),
.B2(n_2633),
.Y(n_3732)
);

O2A1O1Ixp33_ASAP7_75t_L g3733 ( 
.A1(n_3585),
.A2(n_2622),
.B(n_2620),
.C(n_2865),
.Y(n_3733)
);

INVxp67_ASAP7_75t_SL g3734 ( 
.A(n_3654),
.Y(n_3734)
);

O2A1O1Ixp5_ASAP7_75t_L g3735 ( 
.A1(n_3193),
.A2(n_2964),
.B(n_3027),
.C(n_2928),
.Y(n_3735)
);

O2A1O1Ixp33_ASAP7_75t_L g3736 ( 
.A1(n_3206),
.A2(n_2938),
.B(n_2869),
.C(n_2990),
.Y(n_3736)
);

NOR3xp33_ASAP7_75t_SL g3737 ( 
.A(n_3235),
.B(n_2790),
.C(n_2766),
.Y(n_3737)
);

NOR2x1_ASAP7_75t_L g3738 ( 
.A(n_3207),
.B(n_2947),
.Y(n_3738)
);

HB1xp67_ASAP7_75t_L g3739 ( 
.A(n_3211),
.Y(n_3739)
);

AOI21xp5_ASAP7_75t_L g3740 ( 
.A1(n_3546),
.A2(n_2723),
.B(n_2679),
.Y(n_3740)
);

OAI22xp5_ASAP7_75t_L g3741 ( 
.A1(n_3284),
.A2(n_2932),
.B1(n_2944),
.B2(n_2699),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_3644),
.A2(n_2723),
.B(n_2679),
.Y(n_3742)
);

BUFx2_ASAP7_75t_SL g3743 ( 
.A(n_3324),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3200),
.B(n_2724),
.Y(n_3744)
);

A2O1A1Ixp33_ASAP7_75t_L g3745 ( 
.A1(n_3467),
.A2(n_2807),
.B(n_2947),
.C(n_2943),
.Y(n_3745)
);

O2A1O1Ixp33_ASAP7_75t_L g3746 ( 
.A1(n_3286),
.A2(n_3017),
.B(n_3023),
.C(n_2992),
.Y(n_3746)
);

AOI22xp5_ASAP7_75t_L g3747 ( 
.A1(n_3228),
.A2(n_2764),
.B1(n_2765),
.B2(n_2724),
.Y(n_3747)
);

AND2x6_ASAP7_75t_SL g3748 ( 
.A(n_3390),
.B(n_2764),
.Y(n_3748)
);

BUFx6f_ASAP7_75t_L g3749 ( 
.A(n_3507),
.Y(n_3749)
);

AOI22xp5_ASAP7_75t_L g3750 ( 
.A1(n_3541),
.A2(n_2765),
.B1(n_2778),
.B2(n_2768),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3208),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_L g3752 ( 
.A(n_3223),
.B(n_2768),
.Y(n_3752)
);

AND2x4_ASAP7_75t_L g3753 ( 
.A(n_3437),
.B(n_2914),
.Y(n_3753)
);

AOI22xp33_ASAP7_75t_L g3754 ( 
.A1(n_3576),
.A2(n_2778),
.B1(n_2833),
.B2(n_3066),
.Y(n_3754)
);

NOR2xp33_ASAP7_75t_L g3755 ( 
.A(n_3598),
.B(n_2959),
.Y(n_3755)
);

AOI22xp5_ASAP7_75t_L g3756 ( 
.A1(n_3579),
.A2(n_2833),
.B1(n_2806),
.B2(n_2895),
.Y(n_3756)
);

AND3x1_ASAP7_75t_SL g3757 ( 
.A(n_3586),
.B(n_2915),
.C(n_2725),
.Y(n_3757)
);

NOR3xp33_ASAP7_75t_L g3758 ( 
.A(n_3664),
.B(n_3149),
.C(n_3127),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_3275),
.B(n_2887),
.Y(n_3759)
);

NOR2xp33_ASAP7_75t_L g3760 ( 
.A(n_3462),
.B(n_3166),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3642),
.B(n_3295),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_SL g3762 ( 
.A(n_3587),
.B(n_2965),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3296),
.Y(n_3763)
);

AND2x4_ASAP7_75t_L g3764 ( 
.A(n_3445),
.B(n_320),
.Y(n_3764)
);

BUFx6f_ASAP7_75t_L g3765 ( 
.A(n_3246),
.Y(n_3765)
);

NOR2xp33_ASAP7_75t_L g3766 ( 
.A(n_3514),
.B(n_321),
.Y(n_3766)
);

AND2x4_ASAP7_75t_L g3767 ( 
.A(n_3456),
.B(n_321),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3320),
.B(n_321),
.Y(n_3768)
);

INVx1_ASAP7_75t_SL g3769 ( 
.A(n_3238),
.Y(n_3769)
);

O2A1O1Ixp33_ASAP7_75t_L g3770 ( 
.A1(n_3610),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_SL g3771 ( 
.A(n_3666),
.B(n_322),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3543),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3573),
.A2(n_322),
.B(n_323),
.Y(n_3773)
);

A2O1A1Ixp33_ASAP7_75t_SL g3774 ( 
.A1(n_3317),
.A2(n_326),
.B(n_324),
.C(n_325),
.Y(n_3774)
);

OAI21xp33_ASAP7_75t_L g3775 ( 
.A1(n_3551),
.A2(n_324),
.B(n_325),
.Y(n_3775)
);

INVx2_ASAP7_75t_SL g3776 ( 
.A(n_3392),
.Y(n_3776)
);

BUFx6f_ASAP7_75t_L g3777 ( 
.A(n_3246),
.Y(n_3777)
);

CKINVDCx8_ASAP7_75t_R g3778 ( 
.A(n_3292),
.Y(n_3778)
);

INVx2_ASAP7_75t_SL g3779 ( 
.A(n_3442),
.Y(n_3779)
);

AOI22xp33_ASAP7_75t_L g3780 ( 
.A1(n_3606),
.A2(n_328),
.B1(n_325),
.B2(n_327),
.Y(n_3780)
);

OAI22xp5_ASAP7_75t_SL g3781 ( 
.A1(n_3277),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_3781)
);

INVx3_ASAP7_75t_L g3782 ( 
.A(n_3207),
.Y(n_3782)
);

OAI21x1_ASAP7_75t_L g3783 ( 
.A1(n_3179),
.A2(n_332),
.B(n_331),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3362),
.B(n_330),
.Y(n_3784)
);

NAND2x1p5_ASAP7_75t_L g3785 ( 
.A(n_3194),
.B(n_330),
.Y(n_3785)
);

INVx3_ASAP7_75t_L g3786 ( 
.A(n_3639),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3368),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3376),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3384),
.Y(n_3789)
);

OAI22xp5_ASAP7_75t_L g3790 ( 
.A1(n_3292),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3394),
.Y(n_3791)
);

AOI22xp5_ASAP7_75t_L g3792 ( 
.A1(n_3579),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_3792)
);

OAI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_3294),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_3793)
);

INVx1_ASAP7_75t_SL g3794 ( 
.A(n_3294),
.Y(n_3794)
);

CKINVDCx5p33_ASAP7_75t_R g3795 ( 
.A(n_3309),
.Y(n_3795)
);

O2A1O1Ixp33_ASAP7_75t_L g3796 ( 
.A1(n_3234),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_3796)
);

AOI22xp5_ASAP7_75t_L g3797 ( 
.A1(n_3579),
.A2(n_339),
.B1(n_336),
.B2(n_338),
.Y(n_3797)
);

AOI22xp5_ASAP7_75t_L g3798 ( 
.A1(n_3579),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_3798)
);

O2A1O1Ixp33_ASAP7_75t_L g3799 ( 
.A1(n_3262),
.A2(n_342),
.B(n_339),
.C(n_340),
.Y(n_3799)
);

AOI21xp5_ASAP7_75t_L g3800 ( 
.A1(n_3566),
.A2(n_340),
.B(n_342),
.Y(n_3800)
);

AOI21xp5_ASAP7_75t_L g3801 ( 
.A1(n_3212),
.A2(n_342),
.B(n_343),
.Y(n_3801)
);

CKINVDCx11_ASAP7_75t_R g3802 ( 
.A(n_3338),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3395),
.Y(n_3803)
);

A2O1A1Ixp33_ASAP7_75t_L g3804 ( 
.A1(n_3210),
.A2(n_345),
.B(n_343),
.C(n_344),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3553),
.Y(n_3805)
);

BUFx3_ASAP7_75t_L g3806 ( 
.A(n_3528),
.Y(n_3806)
);

NAND3xp33_ASAP7_75t_SL g3807 ( 
.A(n_3258),
.B(n_343),
.C(n_344),
.Y(n_3807)
);

A2O1A1Ixp33_ASAP7_75t_L g3808 ( 
.A1(n_3237),
.A2(n_3257),
.B(n_3261),
.C(n_3232),
.Y(n_3808)
);

O2A1O1Ixp33_ASAP7_75t_L g3809 ( 
.A1(n_3647),
.A2(n_346),
.B(n_344),
.C(n_345),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3397),
.Y(n_3810)
);

AOI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_3520),
.A2(n_346),
.B(n_347),
.Y(n_3811)
);

OA22x2_ASAP7_75t_L g3812 ( 
.A1(n_3338),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_3812)
);

O2A1O1Ixp33_ASAP7_75t_L g3813 ( 
.A1(n_3648),
.A2(n_349),
.B(n_347),
.C(n_348),
.Y(n_3813)
);

AOI22xp33_ASAP7_75t_L g3814 ( 
.A1(n_3633),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.Y(n_3814)
);

AOI22xp33_ASAP7_75t_L g3815 ( 
.A1(n_3355),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_3815)
);

O2A1O1Ixp33_ASAP7_75t_L g3816 ( 
.A1(n_3336),
.A2(n_3342),
.B(n_3341),
.C(n_3607),
.Y(n_3816)
);

AND2x2_ASAP7_75t_L g3817 ( 
.A(n_3321),
.B(n_352),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3412),
.B(n_353),
.Y(n_3818)
);

INVxp67_ASAP7_75t_L g3819 ( 
.A(n_3524),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3572),
.Y(n_3820)
);

INVx3_ASAP7_75t_SL g3821 ( 
.A(n_3217),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_3661),
.A2(n_353),
.B(n_354),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3427),
.B(n_354),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_3666),
.B(n_355),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_SL g3825 ( 
.A(n_3271),
.B(n_355),
.Y(n_3825)
);

OAI21x1_ASAP7_75t_L g3826 ( 
.A1(n_3652),
.A2(n_359),
.B(n_358),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_SL g3827 ( 
.A(n_3274),
.B(n_3657),
.Y(n_3827)
);

NOR2xp33_ASAP7_75t_R g3828 ( 
.A(n_3528),
.B(n_359),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3441),
.B(n_360),
.Y(n_3829)
);

AO32x1_ASAP7_75t_L g3830 ( 
.A1(n_3658),
.A2(n_363),
.A3(n_361),
.B1(n_362),
.B2(n_364),
.Y(n_3830)
);

BUFx12f_ASAP7_75t_L g3831 ( 
.A(n_3195),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3440),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3450),
.B(n_3465),
.Y(n_3833)
);

NOR2xp33_ASAP7_75t_L g3834 ( 
.A(n_3581),
.B(n_361),
.Y(n_3834)
);

OAI22xp5_ASAP7_75t_L g3835 ( 
.A1(n_3618),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.Y(n_3835)
);

AOI22xp33_ASAP7_75t_L g3836 ( 
.A1(n_3540),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_3836)
);

OAI22x1_ASAP7_75t_L g3837 ( 
.A1(n_3657),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3472),
.Y(n_3838)
);

NOR2xp67_ASAP7_75t_L g3839 ( 
.A(n_3627),
.B(n_367),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3591),
.Y(n_3840)
);

BUFx12f_ASAP7_75t_L g3841 ( 
.A(n_3226),
.Y(n_3841)
);

CKINVDCx20_ASAP7_75t_R g3842 ( 
.A(n_3391),
.Y(n_3842)
);

AOI221xp5_ASAP7_75t_L g3843 ( 
.A1(n_3481),
.A2(n_371),
.B1(n_369),
.B2(n_370),
.C(n_372),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3533),
.B(n_370),
.Y(n_3844)
);

BUFx6f_ASAP7_75t_L g3845 ( 
.A(n_3246),
.Y(n_3845)
);

AND2x2_ASAP7_75t_L g3846 ( 
.A(n_3459),
.B(n_373),
.Y(n_3846)
);

BUFx2_ASAP7_75t_R g3847 ( 
.A(n_3568),
.Y(n_3847)
);

AND2x2_ASAP7_75t_L g3848 ( 
.A(n_3499),
.B(n_373),
.Y(n_3848)
);

BUFx2_ASAP7_75t_L g3849 ( 
.A(n_3564),
.Y(n_3849)
);

OA22x2_ASAP7_75t_L g3850 ( 
.A1(n_3382),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_3850)
);

NOR2xp33_ASAP7_75t_L g3851 ( 
.A(n_3388),
.B(n_375),
.Y(n_3851)
);

NOR2xp33_ASAP7_75t_L g3852 ( 
.A(n_3372),
.B(n_375),
.Y(n_3852)
);

INVx2_ASAP7_75t_SL g3853 ( 
.A(n_3351),
.Y(n_3853)
);

BUFx6f_ASAP7_75t_L g3854 ( 
.A(n_3307),
.Y(n_3854)
);

A2O1A1Ixp33_ASAP7_75t_L g3855 ( 
.A1(n_3424),
.A2(n_378),
.B(n_376),
.C(n_377),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3537),
.B(n_376),
.Y(n_3856)
);

OAI22xp5_ASAP7_75t_L g3857 ( 
.A1(n_3386),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3542),
.B(n_377),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3547),
.B(n_3510),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3420),
.B(n_378),
.Y(n_3860)
);

NOR2xp33_ASAP7_75t_L g3861 ( 
.A(n_3433),
.B(n_379),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3216),
.B(n_379),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3230),
.B(n_380),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3596),
.Y(n_3864)
);

NOR2x1_ASAP7_75t_L g3865 ( 
.A(n_3287),
.B(n_380),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3619),
.Y(n_3866)
);

OR2x6_ASAP7_75t_L g3867 ( 
.A(n_3374),
.B(n_380),
.Y(n_3867)
);

BUFx2_ASAP7_75t_L g3868 ( 
.A(n_3564),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_SL g3869 ( 
.A(n_3307),
.B(n_381),
.Y(n_3869)
);

AOI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_3393),
.A2(n_381),
.B(n_382),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_3243),
.B(n_3245),
.Y(n_3871)
);

AOI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3415),
.A2(n_381),
.B(n_382),
.Y(n_3872)
);

BUFx3_ASAP7_75t_L g3873 ( 
.A(n_3620),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3289),
.B(n_382),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3298),
.B(n_383),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3346),
.Y(n_3876)
);

HB1xp67_ASAP7_75t_L g3877 ( 
.A(n_3351),
.Y(n_3877)
);

OAI22xp5_ASAP7_75t_L g3878 ( 
.A1(n_3443),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_3878)
);

AOI21xp5_ASAP7_75t_L g3879 ( 
.A1(n_3418),
.A2(n_384),
.B(n_386),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3559),
.B(n_386),
.Y(n_3880)
);

NOR2xp33_ASAP7_75t_L g3881 ( 
.A(n_3535),
.B(n_387),
.Y(n_3881)
);

AND2x4_ASAP7_75t_L g3882 ( 
.A(n_3536),
.B(n_387),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3313),
.B(n_387),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3202),
.Y(n_3884)
);

INVx2_ASAP7_75t_L g3885 ( 
.A(n_3249),
.Y(n_3885)
);

OR2x6_ASAP7_75t_L g3886 ( 
.A(n_3475),
.B(n_388),
.Y(n_3886)
);

NAND2x1p5_ASAP7_75t_L g3887 ( 
.A(n_3217),
.B(n_388),
.Y(n_3887)
);

AOI21x1_ASAP7_75t_L g3888 ( 
.A1(n_3597),
.A2(n_746),
.B(n_745),
.Y(n_3888)
);

OAI22xp5_ASAP7_75t_L g3889 ( 
.A1(n_3468),
.A2(n_3478),
.B1(n_3501),
.B2(n_3265),
.Y(n_3889)
);

HB1xp67_ASAP7_75t_L g3890 ( 
.A(n_3536),
.Y(n_3890)
);

NOR3xp33_ASAP7_75t_SL g3891 ( 
.A(n_3215),
.B(n_3630),
.C(n_3612),
.Y(n_3891)
);

O2A1O1Ixp33_ASAP7_75t_L g3892 ( 
.A1(n_3493),
.A2(n_3625),
.B(n_3636),
.C(n_3571),
.Y(n_3892)
);

INVx1_ASAP7_75t_SL g3893 ( 
.A(n_3266),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3645),
.B(n_389),
.Y(n_3894)
);

NOR2xp33_ASAP7_75t_SL g3895 ( 
.A(n_3305),
.B(n_389),
.Y(n_3895)
);

AOI21x1_ASAP7_75t_L g3896 ( 
.A1(n_3601),
.A2(n_746),
.B(n_745),
.Y(n_3896)
);

HB1xp67_ASAP7_75t_L g3897 ( 
.A(n_3563),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3344),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3365),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3367),
.Y(n_3900)
);

INVx2_ASAP7_75t_L g3901 ( 
.A(n_3345),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3505),
.B(n_389),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3180),
.B(n_390),
.Y(n_3903)
);

NOR3xp33_ASAP7_75t_L g3904 ( 
.A(n_3444),
.B(n_390),
.C(n_391),
.Y(n_3904)
);

A2O1A1Ixp33_ASAP7_75t_L g3905 ( 
.A1(n_3435),
.A2(n_393),
.B(n_391),
.C(n_392),
.Y(n_3905)
);

AOI22xp5_ASAP7_75t_L g3906 ( 
.A1(n_3446),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_3906)
);

INVx4_ASAP7_75t_L g3907 ( 
.A(n_3479),
.Y(n_3907)
);

AOI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_3423),
.A2(n_392),
.B(n_394),
.Y(n_3908)
);

AOI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_3469),
.A2(n_394),
.B(n_395),
.Y(n_3909)
);

CKINVDCx5p33_ASAP7_75t_R g3910 ( 
.A(n_3512),
.Y(n_3910)
);

AOI22xp33_ASAP7_75t_L g3911 ( 
.A1(n_3575),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_3911)
);

INVx5_ASAP7_75t_L g3912 ( 
.A(n_3307),
.Y(n_3912)
);

INVx4_ASAP7_75t_L g3913 ( 
.A(n_3584),
.Y(n_3913)
);

AOI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3413),
.A2(n_399),
.B1(n_396),
.B2(n_398),
.Y(n_3914)
);

A2O1A1Ixp33_ASAP7_75t_L g3915 ( 
.A1(n_3185),
.A2(n_401),
.B(n_399),
.C(n_400),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3347),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3470),
.A2(n_401),
.B(n_402),
.Y(n_3917)
);

NOR2xp33_ASAP7_75t_L g3918 ( 
.A(n_3363),
.B(n_402),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3349),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3369),
.B(n_403),
.Y(n_3920)
);

NOR2xp33_ASAP7_75t_L g3921 ( 
.A(n_3650),
.B(n_3660),
.Y(n_3921)
);

AOI21xp5_ASAP7_75t_L g3922 ( 
.A1(n_3516),
.A2(n_403),
.B(n_404),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3356),
.Y(n_3923)
);

AOI21xp5_ASAP7_75t_SL g3924 ( 
.A1(n_3491),
.A2(n_404),
.B(n_405),
.Y(n_3924)
);

OAI22xp5_ASAP7_75t_L g3925 ( 
.A1(n_3429),
.A2(n_3554),
.B1(n_3502),
.B2(n_3561),
.Y(n_3925)
);

OAI22x1_ASAP7_75t_L g3926 ( 
.A1(n_3634),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_3926)
);

BUFx2_ASAP7_75t_L g3927 ( 
.A(n_3584),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3383),
.B(n_406),
.Y(n_3928)
);

CKINVDCx5p33_ASAP7_75t_R g3929 ( 
.A(n_3513),
.Y(n_3929)
);

NOR2xp33_ASAP7_75t_L g3930 ( 
.A(n_3665),
.B(n_406),
.Y(n_3930)
);

AOI22xp33_ASAP7_75t_SL g3931 ( 
.A1(n_3508),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_3931)
);

OR2x6_ASAP7_75t_L g3932 ( 
.A(n_3361),
.B(n_3629),
.Y(n_3932)
);

AOI21x1_ASAP7_75t_L g3933 ( 
.A1(n_3396),
.A2(n_748),
.B(n_747),
.Y(n_3933)
);

AOI21xp5_ASAP7_75t_L g3934 ( 
.A1(n_3330),
.A2(n_408),
.B(n_409),
.Y(n_3934)
);

OAI22xp5_ASAP7_75t_L g3935 ( 
.A1(n_3527),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3373),
.Y(n_3936)
);

BUFx12f_ASAP7_75t_L g3937 ( 
.A(n_3584),
.Y(n_3937)
);

INVx3_ASAP7_75t_L g3938 ( 
.A(n_3589),
.Y(n_3938)
);

AOI21xp5_ASAP7_75t_L g3939 ( 
.A1(n_3348),
.A2(n_410),
.B(n_411),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3204),
.B(n_412),
.Y(n_3940)
);

NAND2xp33_ASAP7_75t_L g3941 ( 
.A(n_3560),
.B(n_413),
.Y(n_3941)
);

AOI21xp5_ASAP7_75t_L g3942 ( 
.A1(n_3352),
.A2(n_413),
.B(n_414),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3276),
.B(n_414),
.Y(n_3943)
);

INVx2_ASAP7_75t_SL g3944 ( 
.A(n_3550),
.Y(n_3944)
);

NOR2xp33_ASAP7_75t_L g3945 ( 
.A(n_3667),
.B(n_3315),
.Y(n_3945)
);

AOI22xp5_ASAP7_75t_L g3946 ( 
.A1(n_3659),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_3946)
);

NOR2xp33_ASAP7_75t_L g3947 ( 
.A(n_3350),
.B(n_415),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_SL g3948 ( 
.A(n_3407),
.B(n_416),
.Y(n_3948)
);

BUFx3_ASAP7_75t_L g3949 ( 
.A(n_3552),
.Y(n_3949)
);

AND2x2_ASAP7_75t_L g3950 ( 
.A(n_3343),
.B(n_417),
.Y(n_3950)
);

AOI21xp5_ASAP7_75t_L g3951 ( 
.A1(n_3283),
.A2(n_417),
.B(n_418),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3218),
.B(n_417),
.Y(n_3952)
);

BUFx12f_ASAP7_75t_L g3953 ( 
.A(n_3407),
.Y(n_3953)
);

NOR2xp33_ASAP7_75t_L g3954 ( 
.A(n_3411),
.B(n_418),
.Y(n_3954)
);

AOI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3401),
.A2(n_418),
.B(n_419),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3378),
.Y(n_3956)
);

AOI21xp5_ASAP7_75t_L g3957 ( 
.A1(n_3389),
.A2(n_419),
.B(n_420),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3224),
.B(n_420),
.Y(n_3958)
);

BUFx6f_ASAP7_75t_L g3959 ( 
.A(n_3407),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_L g3960 ( 
.A1(n_3244),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.Y(n_3960)
);

A2O1A1Ixp33_ASAP7_75t_L g3961 ( 
.A1(n_3358),
.A2(n_425),
.B(n_423),
.C(n_424),
.Y(n_3961)
);

O2A1O1Ixp33_ASAP7_75t_L g3962 ( 
.A1(n_3353),
.A2(n_429),
.B(n_427),
.C(n_428),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3379),
.Y(n_3963)
);

INVx2_ASAP7_75t_L g3964 ( 
.A(n_3310),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3398),
.Y(n_3965)
);

INVx2_ASAP7_75t_L g3966 ( 
.A(n_3421),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3421),
.Y(n_3967)
);

OAI21xp5_ASAP7_75t_L g3968 ( 
.A1(n_3588),
.A2(n_428),
.B(n_430),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3626),
.B(n_430),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3229),
.B(n_3240),
.Y(n_3970)
);

A2O1A1Ixp33_ASAP7_75t_L g3971 ( 
.A1(n_3594),
.A2(n_432),
.B(n_430),
.C(n_431),
.Y(n_3971)
);

O2A1O1Ixp5_ASAP7_75t_L g3972 ( 
.A1(n_3290),
.A2(n_433),
.B(n_431),
.C(n_432),
.Y(n_3972)
);

BUFx6f_ASAP7_75t_L g3973 ( 
.A(n_3421),
.Y(n_3973)
);

AOI221xp5_ASAP7_75t_L g3974 ( 
.A1(n_3544),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.C(n_436),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_SL g3975 ( 
.A(n_3477),
.B(n_3498),
.Y(n_3975)
);

BUFx4_ASAP7_75t_SL g3976 ( 
.A(n_3263),
.Y(n_3976)
);

AOI22xp33_ASAP7_75t_L g3977 ( 
.A1(n_3461),
.A2(n_437),
.B1(n_434),
.B2(n_435),
.Y(n_3977)
);

OAI22xp5_ASAP7_75t_L g3978 ( 
.A1(n_3637),
.A2(n_438),
.B1(n_435),
.B2(n_437),
.Y(n_3978)
);

AOI22xp5_ASAP7_75t_L g3979 ( 
.A1(n_3370),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_3979)
);

NOR2xp33_ASAP7_75t_L g3980 ( 
.A(n_3484),
.B(n_439),
.Y(n_3980)
);

A2O1A1Ixp33_ASAP7_75t_L g3981 ( 
.A1(n_3273),
.A2(n_3519),
.B(n_3311),
.C(n_3425),
.Y(n_3981)
);

HB1xp67_ASAP7_75t_L g3982 ( 
.A(n_3485),
.Y(n_3982)
);

BUFx6f_ASAP7_75t_L g3983 ( 
.A(n_3477),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3241),
.B(n_440),
.Y(n_3984)
);

BUFx6f_ASAP7_75t_L g3985 ( 
.A(n_3477),
.Y(n_3985)
);

AOI21xp5_ASAP7_75t_L g3986 ( 
.A1(n_3640),
.A2(n_3250),
.B(n_3248),
.Y(n_3986)
);

NOR2xp33_ASAP7_75t_L g3987 ( 
.A(n_3494),
.B(n_441),
.Y(n_3987)
);

AOI22x1_ASAP7_75t_L g3988 ( 
.A1(n_3282),
.A2(n_3259),
.B1(n_3260),
.B2(n_3221),
.Y(n_3988)
);

AOI21xp5_ASAP7_75t_L g3989 ( 
.A1(n_3253),
.A2(n_442),
.B(n_443),
.Y(n_3989)
);

NOR2xp33_ASAP7_75t_L g3990 ( 
.A(n_3497),
.B(n_442),
.Y(n_3990)
);

INVx2_ASAP7_75t_L g3991 ( 
.A(n_3498),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3615),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_3992)
);

NOR2xp33_ASAP7_75t_SL g3993 ( 
.A(n_3614),
.B(n_444),
.Y(n_3993)
);

O2A1O1Ixp33_ASAP7_75t_L g3994 ( 
.A1(n_3622),
.A2(n_447),
.B(n_445),
.C(n_446),
.Y(n_3994)
);

BUFx6f_ASAP7_75t_L g3995 ( 
.A(n_3498),
.Y(n_3995)
);

AOI22x1_ASAP7_75t_L g3996 ( 
.A1(n_3631),
.A2(n_447),
.B1(n_445),
.B2(n_446),
.Y(n_3996)
);

AND2x4_ASAP7_75t_L g3997 ( 
.A(n_3602),
.B(n_448),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3254),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3399),
.Y(n_3999)
);

NOR2x1_ASAP7_75t_L g4000 ( 
.A(n_3267),
.B(n_3656),
.Y(n_4000)
);

NOR2xp33_ASAP7_75t_SL g4001 ( 
.A(n_3557),
.B(n_448),
.Y(n_4001)
);

NOR2xp33_ASAP7_75t_L g4002 ( 
.A(n_3503),
.B(n_3635),
.Y(n_4002)
);

CKINVDCx5p33_ASAP7_75t_R g4003 ( 
.A(n_3308),
.Y(n_4003)
);

AOI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_3255),
.A2(n_3280),
.B(n_3264),
.Y(n_4004)
);

AND2x2_ASAP7_75t_L g4005 ( 
.A(n_3306),
.B(n_450),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_SL g4006 ( 
.A(n_3643),
.B(n_450),
.Y(n_4006)
);

BUFx6f_ASAP7_75t_L g4007 ( 
.A(n_3557),
.Y(n_4007)
);

AOI21xp5_ASAP7_75t_L g4008 ( 
.A1(n_3281),
.A2(n_451),
.B(n_452),
.Y(n_4008)
);

OAI22xp5_ASAP7_75t_L g4009 ( 
.A1(n_3205),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3480),
.B(n_451),
.Y(n_4010)
);

AOI21xp5_ASAP7_75t_L g4011 ( 
.A1(n_3291),
.A2(n_453),
.B(n_454),
.Y(n_4011)
);

NOR2xp33_ASAP7_75t_L g4012 ( 
.A(n_3483),
.B(n_3534),
.Y(n_4012)
);

AOI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_3293),
.A2(n_3304),
.B(n_3299),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3318),
.B(n_455),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_SL g4015 ( 
.A(n_3643),
.B(n_455),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3322),
.B(n_455),
.Y(n_4016)
);

AOI22xp33_ASAP7_75t_L g4017 ( 
.A1(n_3268),
.A2(n_458),
.B1(n_456),
.B2(n_457),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_SL g4018 ( 
.A(n_3474),
.B(n_456),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3323),
.B(n_456),
.Y(n_4019)
);

BUFx8_ASAP7_75t_L g4020 ( 
.A(n_3302),
.Y(n_4020)
);

OAI21x1_ASAP7_75t_L g4021 ( 
.A1(n_3529),
.A2(n_460),
.B(n_459),
.Y(n_4021)
);

AOI21xp5_ASAP7_75t_L g4022 ( 
.A1(n_3331),
.A2(n_457),
.B(n_460),
.Y(n_4022)
);

A2O1A1Ixp33_ASAP7_75t_L g4023 ( 
.A1(n_3316),
.A2(n_462),
.B(n_460),
.C(n_461),
.Y(n_4023)
);

HB1xp67_ASAP7_75t_L g4024 ( 
.A(n_3333),
.Y(n_4024)
);

AOI22xp5_ASAP7_75t_L g4025 ( 
.A1(n_3548),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.Y(n_4025)
);

AOI21xp5_ASAP7_75t_L g4026 ( 
.A1(n_3624),
.A2(n_464),
.B(n_465),
.Y(n_4026)
);

AOI21xp5_ASAP7_75t_L g4027 ( 
.A1(n_3632),
.A2(n_464),
.B(n_465),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3400),
.Y(n_4028)
);

NAND2x1p5_ASAP7_75t_L g4029 ( 
.A(n_3557),
.B(n_466),
.Y(n_4029)
);

AOI21x1_ASAP7_75t_L g4030 ( 
.A1(n_3651),
.A2(n_750),
.B(n_749),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_SL g4031 ( 
.A(n_3558),
.B(n_466),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3410),
.B(n_466),
.Y(n_4032)
);

CKINVDCx20_ASAP7_75t_R g4033 ( 
.A(n_3555),
.Y(n_4033)
);

OAI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_3404),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.Y(n_4034)
);

OR2x2_ASAP7_75t_L g4035 ( 
.A(n_3419),
.B(n_467),
.Y(n_4035)
);

INVxp67_ASAP7_75t_L g4036 ( 
.A(n_3426),
.Y(n_4036)
);

AOI21xp5_ASAP7_75t_L g4037 ( 
.A1(n_3641),
.A2(n_3649),
.B(n_3213),
.Y(n_4037)
);

INVx2_ASAP7_75t_SL g4038 ( 
.A(n_3646),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3432),
.B(n_468),
.Y(n_4039)
);

BUFx6f_ASAP7_75t_L g4040 ( 
.A(n_3558),
.Y(n_4040)
);

HB1xp67_ASAP7_75t_L g4041 ( 
.A(n_3438),
.Y(n_4041)
);

NOR2xp33_ASAP7_75t_L g4042 ( 
.A(n_3439),
.B(n_468),
.Y(n_4042)
);

AOI21xp5_ASAP7_75t_L g4043 ( 
.A1(n_3279),
.A2(n_469),
.B(n_470),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_3448),
.B(n_470),
.Y(n_4044)
);

AOI21xp5_ASAP7_75t_L g4045 ( 
.A1(n_3242),
.A2(n_470),
.B(n_471),
.Y(n_4045)
);

INVx3_ASAP7_75t_SL g4046 ( 
.A(n_3558),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3452),
.B(n_471),
.Y(n_4047)
);

NOR2xp33_ASAP7_75t_L g4048 ( 
.A(n_3457),
.B(n_471),
.Y(n_4048)
);

HB1xp67_ASAP7_75t_L g4049 ( 
.A(n_3460),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3466),
.B(n_472),
.Y(n_4050)
);

AOI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_3251),
.A2(n_472),
.B(n_474),
.Y(n_4051)
);

AOI21xp5_ASAP7_75t_L g4052 ( 
.A1(n_3222),
.A2(n_475),
.B(n_476),
.Y(n_4052)
);

O2A1O1Ixp33_ASAP7_75t_L g4053 ( 
.A1(n_3405),
.A2(n_478),
.B(n_475),
.C(n_477),
.Y(n_4053)
);

INVx3_ASAP7_75t_L g4054 ( 
.A(n_3375),
.Y(n_4054)
);

OAI22xp5_ASAP7_75t_L g4055 ( 
.A1(n_3417),
.A2(n_479),
.B1(n_477),
.B2(n_478),
.Y(n_4055)
);

NAND2x1p5_ASAP7_75t_L g4056 ( 
.A(n_3628),
.B(n_477),
.Y(n_4056)
);

AO21x2_ASAP7_75t_L g4057 ( 
.A1(n_3332),
.A2(n_478),
.B(n_480),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3471),
.Y(n_4058)
);

A2O1A1Ixp33_ASAP7_75t_L g4059 ( 
.A1(n_3638),
.A2(n_3312),
.B(n_3303),
.C(n_3236),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3515),
.B(n_480),
.Y(n_4060)
);

AOI21xp5_ASAP7_75t_L g4061 ( 
.A1(n_3225),
.A2(n_481),
.B(n_482),
.Y(n_4061)
);

AOI21xp5_ASAP7_75t_L g4062 ( 
.A1(n_3496),
.A2(n_481),
.B(n_482),
.Y(n_4062)
);

HB1xp67_ASAP7_75t_L g4063 ( 
.A(n_3521),
.Y(n_4063)
);

BUFx12f_ASAP7_75t_L g4064 ( 
.A(n_3302),
.Y(n_4064)
);

NOR2xp33_ASAP7_75t_L g4065 ( 
.A(n_3530),
.B(n_3532),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_3302),
.B(n_3538),
.Y(n_4066)
);

INVx2_ASAP7_75t_L g4067 ( 
.A(n_3506),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_3578),
.B(n_483),
.Y(n_4068)
);

NOR2xp33_ASAP7_75t_L g4069 ( 
.A(n_3574),
.B(n_483),
.Y(n_4069)
);

NOR2xp33_ASAP7_75t_L g4070 ( 
.A(n_3590),
.B(n_483),
.Y(n_4070)
);

INVx4_ASAP7_75t_L g4071 ( 
.A(n_3621),
.Y(n_4071)
);

CKINVDCx14_ASAP7_75t_R g4072 ( 
.A(n_3592),
.Y(n_4072)
);

BUFx2_ASAP7_75t_L g4073 ( 
.A(n_3593),
.Y(n_4073)
);

OAI221xp5_ASAP7_75t_L g4074 ( 
.A1(n_3511),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.C(n_487),
.Y(n_4074)
);

OA21x2_ASAP7_75t_L g4075 ( 
.A1(n_3354),
.A2(n_484),
.B(n_485),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3613),
.Y(n_4076)
);

AND2x2_ASAP7_75t_L g4077 ( 
.A(n_3569),
.B(n_486),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3371),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_SL g4079 ( 
.A(n_3422),
.B(n_486),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_SL g4080 ( 
.A(n_3605),
.B(n_487),
.Y(n_4080)
);

AO21x1_ASAP7_75t_L g4081 ( 
.A1(n_3239),
.A2(n_3196),
.B(n_3186),
.Y(n_4081)
);

O2A1O1Ixp33_ASAP7_75t_L g4082 ( 
.A1(n_3434),
.A2(n_490),
.B(n_488),
.C(n_489),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3570),
.Y(n_4083)
);

NOR2xp33_ASAP7_75t_L g4084 ( 
.A(n_3662),
.B(n_488),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3556),
.B(n_488),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3567),
.B(n_489),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_3453),
.B(n_489),
.Y(n_4087)
);

INVx2_ASAP7_75t_SL g4088 ( 
.A(n_3487),
.Y(n_4088)
);

INVx4_ASAP7_75t_L g4089 ( 
.A(n_3455),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_SL g4090 ( 
.A(n_3199),
.B(n_490),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3496),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_3278),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3663),
.B(n_3595),
.Y(n_4093)
);

BUFx2_ASAP7_75t_SL g4094 ( 
.A(n_3490),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3464),
.B(n_491),
.Y(n_4095)
);

AOI21xp5_ASAP7_75t_L g4096 ( 
.A1(n_3203),
.A2(n_492),
.B(n_493),
.Y(n_4096)
);

NOR3xp33_ASAP7_75t_L g4097 ( 
.A(n_3476),
.B(n_492),
.C(n_493),
.Y(n_4097)
);

A2O1A1Ixp33_ASAP7_75t_L g4098 ( 
.A1(n_3486),
.A2(n_495),
.B(n_492),
.C(n_494),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3454),
.B(n_494),
.Y(n_4099)
);

AOI21xp5_ASAP7_75t_L g4100 ( 
.A1(n_3288),
.A2(n_495),
.B(n_496),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3319),
.Y(n_4101)
);

HB1xp67_ASAP7_75t_L g4102 ( 
.A(n_3582),
.Y(n_4102)
);

O2A1O1Ixp33_ASAP7_75t_L g4103 ( 
.A1(n_3463),
.A2(n_499),
.B(n_497),
.C(n_498),
.Y(n_4103)
);

O2A1O1Ixp33_ASAP7_75t_L g4104 ( 
.A1(n_3504),
.A2(n_499),
.B(n_497),
.C(n_498),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_3447),
.B(n_3449),
.Y(n_4105)
);

OAI22xp5_ASAP7_75t_L g4106 ( 
.A1(n_3326),
.A2(n_500),
.B1(n_498),
.B2(n_499),
.Y(n_4106)
);

OR2x2_ASAP7_75t_L g4107 ( 
.A(n_3451),
.B(n_500),
.Y(n_4107)
);

AOI21xp5_ASAP7_75t_L g4108 ( 
.A1(n_3297),
.A2(n_501),
.B(n_502),
.Y(n_4108)
);

O2A1O1Ixp33_ASAP7_75t_L g4109 ( 
.A1(n_3509),
.A2(n_503),
.B(n_501),
.C(n_502),
.Y(n_4109)
);

INVx2_ASAP7_75t_L g4110 ( 
.A(n_3301),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_3327),
.Y(n_4111)
);

AOI22xp5_ASAP7_75t_L g4112 ( 
.A1(n_3328),
.A2(n_3334),
.B1(n_3335),
.B2(n_3329),
.Y(n_4112)
);

AOI21xp5_ASAP7_75t_L g4113 ( 
.A1(n_3359),
.A2(n_503),
.B(n_504),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_3364),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3366),
.B(n_503),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3377),
.Y(n_4116)
);

BUFx6f_ASAP7_75t_L g4117 ( 
.A(n_3599),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_3385),
.Y(n_4118)
);

AND2x4_ASAP7_75t_L g4119 ( 
.A(n_3387),
.B(n_504),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_3402),
.B(n_506),
.Y(n_4120)
);

AO32x2_ASAP7_75t_L g4121 ( 
.A1(n_3403),
.A2(n_509),
.A3(n_507),
.B1(n_508),
.B2(n_510),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_SL g4122 ( 
.A(n_3408),
.B(n_508),
.Y(n_4122)
);

AND2x6_ASAP7_75t_L g4123 ( 
.A(n_3409),
.B(n_509),
.Y(n_4123)
);

INVx3_ASAP7_75t_L g4124 ( 
.A(n_3430),
.Y(n_4124)
);

A2O1A1Ixp33_ASAP7_75t_L g4125 ( 
.A1(n_3523),
.A2(n_511),
.B(n_509),
.C(n_510),
.Y(n_4125)
);

AOI21xp5_ASAP7_75t_L g4126 ( 
.A1(n_3525),
.A2(n_510),
.B(n_511),
.Y(n_4126)
);

INVx1_ASAP7_75t_SL g4127 ( 
.A(n_3600),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3526),
.Y(n_4128)
);

AOI21xp5_ASAP7_75t_L g4129 ( 
.A1(n_3531),
.A2(n_511),
.B(n_512),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_3603),
.Y(n_4130)
);

AOI22xp33_ASAP7_75t_L g4131 ( 
.A1(n_3655),
.A2(n_514),
.B1(n_512),
.B2(n_513),
.Y(n_4131)
);

OAI22xp5_ASAP7_75t_L g4132 ( 
.A1(n_3604),
.A2(n_514),
.B1(n_512),
.B2(n_513),
.Y(n_4132)
);

OAI21xp5_ASAP7_75t_L g4133 ( 
.A1(n_3609),
.A2(n_515),
.B(n_516),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3611),
.B(n_515),
.Y(n_4134)
);

OAI22xp5_ASAP7_75t_L g4135 ( 
.A1(n_3623),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_4135)
);

AOI21xp5_ASAP7_75t_L g4136 ( 
.A1(n_3616),
.A2(n_516),
.B(n_517),
.Y(n_4136)
);

AOI21xp5_ASAP7_75t_L g4137 ( 
.A1(n_3617),
.A2(n_518),
.B(n_519),
.Y(n_4137)
);

O2A1O1Ixp5_ASAP7_75t_L g4138 ( 
.A1(n_3193),
.A2(n_520),
.B(n_518),
.C(n_519),
.Y(n_4138)
);

BUFx2_ASAP7_75t_L g4139 ( 
.A(n_3219),
.Y(n_4139)
);

INVx5_ASAP7_75t_L g4140 ( 
.A(n_3227),
.Y(n_4140)
);

NOR3xp33_ASAP7_75t_L g4141 ( 
.A(n_3181),
.B(n_520),
.C(n_521),
.Y(n_4141)
);

NOR2xp33_ASAP7_75t_SL g4142 ( 
.A(n_3189),
.B(n_520),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_3178),
.B(n_521),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_3187),
.Y(n_4144)
);

O2A1O1Ixp33_ASAP7_75t_L g4145 ( 
.A1(n_3181),
.A2(n_524),
.B(n_522),
.C(n_523),
.Y(n_4145)
);

BUFx6f_ASAP7_75t_L g4146 ( 
.A(n_3227),
.Y(n_4146)
);

NOR2xp33_ASAP7_75t_L g4147 ( 
.A(n_3539),
.B(n_522),
.Y(n_4147)
);

NAND2xp33_ASAP7_75t_SL g4148 ( 
.A(n_3357),
.B(n_523),
.Y(n_4148)
);

INVx2_ASAP7_75t_SL g4149 ( 
.A(n_4140),
.Y(n_4149)
);

BUFx6f_ASAP7_75t_L g4150 ( 
.A(n_3681),
.Y(n_4150)
);

INVx2_ASAP7_75t_SL g4151 ( 
.A(n_4140),
.Y(n_4151)
);

BUFx6f_ASAP7_75t_L g4152 ( 
.A(n_3681),
.Y(n_4152)
);

BUFx6f_ASAP7_75t_L g4153 ( 
.A(n_3722),
.Y(n_4153)
);

BUFx6f_ASAP7_75t_L g4154 ( 
.A(n_3722),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3706),
.Y(n_4155)
);

INVx3_ASAP7_75t_L g4156 ( 
.A(n_3726),
.Y(n_4156)
);

CKINVDCx11_ASAP7_75t_R g4157 ( 
.A(n_3683),
.Y(n_4157)
);

BUFx6f_ASAP7_75t_L g4158 ( 
.A(n_3677),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3708),
.Y(n_4159)
);

INVxp67_ASAP7_75t_SL g4160 ( 
.A(n_3694),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3751),
.Y(n_4161)
);

BUFx3_ASAP7_75t_L g4162 ( 
.A(n_4140),
.Y(n_4162)
);

AND2x4_ASAP7_75t_L g4163 ( 
.A(n_3701),
.B(n_526),
.Y(n_4163)
);

BUFx2_ASAP7_75t_L g4164 ( 
.A(n_3953),
.Y(n_4164)
);

BUFx3_ASAP7_75t_L g4165 ( 
.A(n_3677),
.Y(n_4165)
);

BUFx2_ASAP7_75t_L g4166 ( 
.A(n_3765),
.Y(n_4166)
);

INVx2_ASAP7_75t_SL g4167 ( 
.A(n_3689),
.Y(n_4167)
);

CKINVDCx16_ASAP7_75t_R g4168 ( 
.A(n_3828),
.Y(n_4168)
);

INVx2_ASAP7_75t_L g4169 ( 
.A(n_3684),
.Y(n_4169)
);

BUFx2_ASAP7_75t_SL g4170 ( 
.A(n_3701),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3763),
.Y(n_4171)
);

BUFx12f_ASAP7_75t_L g4172 ( 
.A(n_4146),
.Y(n_4172)
);

BUFx3_ASAP7_75t_L g4173 ( 
.A(n_3729),
.Y(n_4173)
);

BUFx2_ASAP7_75t_SL g4174 ( 
.A(n_3701),
.Y(n_4174)
);

INVx2_ASAP7_75t_L g4175 ( 
.A(n_3691),
.Y(n_4175)
);

BUFx3_ASAP7_75t_L g4176 ( 
.A(n_3729),
.Y(n_4176)
);

INVx1_ASAP7_75t_SL g4177 ( 
.A(n_3802),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_3787),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_3685),
.B(n_525),
.Y(n_4179)
);

BUFx3_ASAP7_75t_L g4180 ( 
.A(n_3749),
.Y(n_4180)
);

BUFx6f_ASAP7_75t_SL g4181 ( 
.A(n_4146),
.Y(n_4181)
);

BUFx6f_ASAP7_75t_L g4182 ( 
.A(n_3937),
.Y(n_4182)
);

INVx3_ASAP7_75t_L g4183 ( 
.A(n_3841),
.Y(n_4183)
);

BUFx2_ASAP7_75t_L g4184 ( 
.A(n_4139),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_3692),
.Y(n_4185)
);

BUFx3_ASAP7_75t_L g4186 ( 
.A(n_3749),
.Y(n_4186)
);

INVx1_ASAP7_75t_SL g4187 ( 
.A(n_3743),
.Y(n_4187)
);

BUFx2_ASAP7_75t_L g4188 ( 
.A(n_3821),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_3788),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_4066),
.B(n_526),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_SL g4191 ( 
.A(n_3707),
.B(n_526),
.Y(n_4191)
);

INVx3_ASAP7_75t_L g4192 ( 
.A(n_3778),
.Y(n_4192)
);

BUFx4f_ASAP7_75t_SL g4193 ( 
.A(n_3806),
.Y(n_4193)
);

AOI22xp33_ASAP7_75t_SL g4194 ( 
.A1(n_4020),
.A2(n_529),
.B1(n_527),
.B2(n_528),
.Y(n_4194)
);

INVx5_ASAP7_75t_SL g4195 ( 
.A(n_3867),
.Y(n_4195)
);

INVx3_ASAP7_75t_L g4196 ( 
.A(n_3748),
.Y(n_4196)
);

INVx6_ASAP7_75t_L g4197 ( 
.A(n_3723),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_3789),
.Y(n_4198)
);

BUFx10_ASAP7_75t_L g4199 ( 
.A(n_3727),
.Y(n_4199)
);

INVx2_ASAP7_75t_L g4200 ( 
.A(n_3710),
.Y(n_4200)
);

INVx2_ASAP7_75t_SL g4201 ( 
.A(n_3727),
.Y(n_4201)
);

CKINVDCx6p67_ASAP7_75t_R g4202 ( 
.A(n_3723),
.Y(n_4202)
);

BUFx3_ASAP7_75t_L g4203 ( 
.A(n_3831),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_3791),
.Y(n_4204)
);

INVxp67_ASAP7_75t_SL g4205 ( 
.A(n_3877),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_3803),
.Y(n_4206)
);

OR2x6_ASAP7_75t_L g4207 ( 
.A(n_3867),
.B(n_527),
.Y(n_4207)
);

BUFx6f_ASAP7_75t_L g4208 ( 
.A(n_3873),
.Y(n_4208)
);

BUFx3_ASAP7_75t_L g4209 ( 
.A(n_3670),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_3810),
.Y(n_4210)
);

INVx8_ASAP7_75t_L g4211 ( 
.A(n_3723),
.Y(n_4211)
);

INVxp67_ASAP7_75t_SL g4212 ( 
.A(n_3890),
.Y(n_4212)
);

INVx3_ASAP7_75t_L g4213 ( 
.A(n_3907),
.Y(n_4213)
);

INVx5_ASAP7_75t_L g4214 ( 
.A(n_3886),
.Y(n_4214)
);

BUFx3_ASAP7_75t_L g4215 ( 
.A(n_3676),
.Y(n_4215)
);

BUFx6f_ASAP7_75t_L g4216 ( 
.A(n_4046),
.Y(n_4216)
);

BUFx4f_ASAP7_75t_L g4217 ( 
.A(n_3721),
.Y(n_4217)
);

AND2x2_ASAP7_75t_L g4218 ( 
.A(n_3761),
.B(n_529),
.Y(n_4218)
);

OR2x6_ASAP7_75t_L g4219 ( 
.A(n_3886),
.B(n_529),
.Y(n_4219)
);

BUFx3_ASAP7_75t_L g4220 ( 
.A(n_3776),
.Y(n_4220)
);

INVxp67_ASAP7_75t_SL g4221 ( 
.A(n_3897),
.Y(n_4221)
);

INVx3_ASAP7_75t_SL g4222 ( 
.A(n_3795),
.Y(n_4222)
);

BUFx6f_ASAP7_75t_L g4223 ( 
.A(n_3912),
.Y(n_4223)
);

BUFx3_ASAP7_75t_L g4224 ( 
.A(n_3779),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_3690),
.B(n_530),
.Y(n_4225)
);

BUFx2_ASAP7_75t_L g4226 ( 
.A(n_3711),
.Y(n_4226)
);

AND2x4_ASAP7_75t_L g4227 ( 
.A(n_3674),
.B(n_531),
.Y(n_4227)
);

BUFx2_ASAP7_75t_SL g4228 ( 
.A(n_3707),
.Y(n_4228)
);

INVx1_ASAP7_75t_SL g4229 ( 
.A(n_3769),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3832),
.Y(n_4230)
);

BUFx3_ASAP7_75t_L g4231 ( 
.A(n_3786),
.Y(n_4231)
);

NAND2x1p5_ASAP7_75t_L g4232 ( 
.A(n_3738),
.B(n_530),
.Y(n_4232)
);

INVx3_ASAP7_75t_L g4233 ( 
.A(n_3782),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_3838),
.Y(n_4234)
);

BUFx3_ASAP7_75t_L g4235 ( 
.A(n_3949),
.Y(n_4235)
);

OAI22xp5_ASAP7_75t_L g4236 ( 
.A1(n_3673),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_4236)
);

OR2x6_ASAP7_75t_L g4237 ( 
.A(n_3887),
.B(n_532),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_3668),
.B(n_532),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_3840),
.Y(n_4239)
);

INVx5_ASAP7_75t_L g4240 ( 
.A(n_3912),
.Y(n_4240)
);

INVx3_ASAP7_75t_SL g4241 ( 
.A(n_3842),
.Y(n_4241)
);

BUFx3_ASAP7_75t_L g4242 ( 
.A(n_3739),
.Y(n_4242)
);

INVx2_ASAP7_75t_SL g4243 ( 
.A(n_3732),
.Y(n_4243)
);

BUFx6f_ASAP7_75t_L g4244 ( 
.A(n_3777),
.Y(n_4244)
);

BUFx2_ASAP7_75t_L g4245 ( 
.A(n_3819),
.Y(n_4245)
);

INVx5_ASAP7_75t_L g4246 ( 
.A(n_3932),
.Y(n_4246)
);

BUFx6f_ASAP7_75t_L g4247 ( 
.A(n_3777),
.Y(n_4247)
);

BUFx2_ASAP7_75t_SL g4248 ( 
.A(n_3882),
.Y(n_4248)
);

INVx3_ASAP7_75t_L g4249 ( 
.A(n_3997),
.Y(n_4249)
);

BUFx3_ASAP7_75t_L g4250 ( 
.A(n_3703),
.Y(n_4250)
);

INVxp67_ASAP7_75t_SL g4251 ( 
.A(n_3764),
.Y(n_4251)
);

INVx5_ASAP7_75t_L g4252 ( 
.A(n_3932),
.Y(n_4252)
);

BUFx12f_ASAP7_75t_L g4253 ( 
.A(n_3882),
.Y(n_4253)
);

INVx1_ASAP7_75t_SL g4254 ( 
.A(n_3847),
.Y(n_4254)
);

BUFx12f_ASAP7_75t_L g4255 ( 
.A(n_3785),
.Y(n_4255)
);

INVx5_ASAP7_75t_SL g4256 ( 
.A(n_3764),
.Y(n_4256)
);

BUFx2_ASAP7_75t_L g4257 ( 
.A(n_3765),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_3820),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_3833),
.Y(n_4259)
);

INVx5_ASAP7_75t_L g4260 ( 
.A(n_3845),
.Y(n_4260)
);

INVx4_ASAP7_75t_L g4261 ( 
.A(n_3913),
.Y(n_4261)
);

BUFx3_ASAP7_75t_L g4262 ( 
.A(n_3705),
.Y(n_4262)
);

CKINVDCx5p33_ASAP7_75t_R g4263 ( 
.A(n_3737),
.Y(n_4263)
);

NOR2xp67_ASAP7_75t_SL g4264 ( 
.A(n_3709),
.B(n_3678),
.Y(n_4264)
);

BUFx3_ASAP7_75t_L g4265 ( 
.A(n_3760),
.Y(n_4265)
);

BUFx3_ASAP7_75t_L g4266 ( 
.A(n_3849),
.Y(n_4266)
);

INVx5_ASAP7_75t_L g4267 ( 
.A(n_3845),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_3864),
.Y(n_4268)
);

BUFx12f_ASAP7_75t_L g4269 ( 
.A(n_3910),
.Y(n_4269)
);

BUFx3_ASAP7_75t_L g4270 ( 
.A(n_3868),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_3695),
.B(n_534),
.Y(n_4271)
);

CKINVDCx5p33_ASAP7_75t_R g4272 ( 
.A(n_3929),
.Y(n_4272)
);

BUFx24_ASAP7_75t_L g4273 ( 
.A(n_3767),
.Y(n_4273)
);

INVx2_ASAP7_75t_SL g4274 ( 
.A(n_3853),
.Y(n_4274)
);

AND2x2_ASAP7_75t_L g4275 ( 
.A(n_3772),
.B(n_535),
.Y(n_4275)
);

BUFx3_ASAP7_75t_L g4276 ( 
.A(n_3927),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_3866),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_3805),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_3982),
.B(n_535),
.Y(n_4279)
);

BUFx3_ASAP7_75t_L g4280 ( 
.A(n_3944),
.Y(n_4280)
);

AND2x4_ASAP7_75t_L g4281 ( 
.A(n_3794),
.B(n_536),
.Y(n_4281)
);

BUFx6f_ASAP7_75t_L g4282 ( 
.A(n_3854),
.Y(n_4282)
);

BUFx6f_ASAP7_75t_L g4283 ( 
.A(n_3854),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_4144),
.B(n_535),
.Y(n_4284)
);

INVx5_ASAP7_75t_SL g4285 ( 
.A(n_3767),
.Y(n_4285)
);

INVx5_ASAP7_75t_L g4286 ( 
.A(n_3959),
.Y(n_4286)
);

BUFx6f_ASAP7_75t_L g4287 ( 
.A(n_3959),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_3884),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_3885),
.Y(n_4289)
);

NOR2xp33_ASAP7_75t_L g4290 ( 
.A(n_4072),
.B(n_3762),
.Y(n_4290)
);

INVx1_ASAP7_75t_SL g4291 ( 
.A(n_3893),
.Y(n_4291)
);

BUFx3_ASAP7_75t_L g4292 ( 
.A(n_3753),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_3898),
.Y(n_4293)
);

CKINVDCx5p33_ASAP7_75t_R g4294 ( 
.A(n_3834),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_3901),
.Y(n_4295)
);

BUFx8_ASAP7_75t_L g4296 ( 
.A(n_3894),
.Y(n_4296)
);

INVx2_ASAP7_75t_L g4297 ( 
.A(n_3916),
.Y(n_4297)
);

OR2x2_ASAP7_75t_L g4298 ( 
.A(n_3679),
.B(n_536),
.Y(n_4298)
);

INVx2_ASAP7_75t_SL g4299 ( 
.A(n_3714),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_3919),
.Y(n_4300)
);

BUFx3_ASAP7_75t_L g4301 ( 
.A(n_3753),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_3876),
.B(n_537),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_3923),
.Y(n_4303)
);

BUFx3_ASAP7_75t_L g4304 ( 
.A(n_4033),
.Y(n_4304)
);

INVx8_ASAP7_75t_L g4305 ( 
.A(n_3713),
.Y(n_4305)
);

BUFx3_ASAP7_75t_L g4306 ( 
.A(n_3755),
.Y(n_4306)
);

INVx1_ASAP7_75t_SL g4307 ( 
.A(n_3817),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_3826),
.Y(n_4308)
);

BUFx2_ASAP7_75t_L g4309 ( 
.A(n_3734),
.Y(n_4309)
);

INVx3_ASAP7_75t_SL g4310 ( 
.A(n_3716),
.Y(n_4310)
);

INVx3_ASAP7_75t_L g4311 ( 
.A(n_3938),
.Y(n_4311)
);

BUFx3_ASAP7_75t_L g4312 ( 
.A(n_3829),
.Y(n_4312)
);

BUFx10_ASAP7_75t_L g4313 ( 
.A(n_3766),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_3899),
.B(n_537),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_3759),
.Y(n_4315)
);

BUFx4_ASAP7_75t_SL g4316 ( 
.A(n_3687),
.Y(n_4316)
);

BUFx3_ASAP7_75t_L g4317 ( 
.A(n_3846),
.Y(n_4317)
);

CKINVDCx20_ASAP7_75t_R g4318 ( 
.A(n_3757),
.Y(n_4318)
);

NAND2x1p5_ASAP7_75t_L g4319 ( 
.A(n_3688),
.B(n_537),
.Y(n_4319)
);

BUFx6f_ASAP7_75t_L g4320 ( 
.A(n_3973),
.Y(n_4320)
);

INVx3_ASAP7_75t_SL g4321 ( 
.A(n_3812),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_3998),
.Y(n_4322)
);

CKINVDCx11_ASAP7_75t_R g4323 ( 
.A(n_3983),
.Y(n_4323)
);

BUFx2_ASAP7_75t_L g4324 ( 
.A(n_3983),
.Y(n_4324)
);

INVx1_ASAP7_75t_SL g4325 ( 
.A(n_3848),
.Y(n_4325)
);

INVx4_ASAP7_75t_L g4326 ( 
.A(n_3985),
.Y(n_4326)
);

INVx3_ASAP7_75t_SL g4327 ( 
.A(n_3985),
.Y(n_4327)
);

BUFx6f_ASAP7_75t_L g4328 ( 
.A(n_3995),
.Y(n_4328)
);

INVxp67_ASAP7_75t_SL g4329 ( 
.A(n_3671),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_3744),
.Y(n_4330)
);

INVx3_ASAP7_75t_L g4331 ( 
.A(n_4038),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_3900),
.B(n_538),
.Y(n_4332)
);

INVx2_ASAP7_75t_SL g4333 ( 
.A(n_3995),
.Y(n_4333)
);

BUFx2_ASAP7_75t_L g4334 ( 
.A(n_3765),
.Y(n_4334)
);

BUFx3_ASAP7_75t_L g4335 ( 
.A(n_4040),
.Y(n_4335)
);

INVx3_ASAP7_75t_SL g4336 ( 
.A(n_4003),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_3752),
.Y(n_4337)
);

NAND2x1p5_ASAP7_75t_L g4338 ( 
.A(n_3792),
.B(n_538),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_3768),
.Y(n_4339)
);

CKINVDCx11_ASAP7_75t_R g4340 ( 
.A(n_4064),
.Y(n_4340)
);

INVx3_ASAP7_75t_L g4341 ( 
.A(n_4029),
.Y(n_4341)
);

BUFx4f_ASAP7_75t_SL g4342 ( 
.A(n_3827),
.Y(n_4342)
);

INVx1_ASAP7_75t_SL g4343 ( 
.A(n_3698),
.Y(n_4343)
);

INVxp67_ASAP7_75t_SL g4344 ( 
.A(n_4024),
.Y(n_4344)
);

INVx8_ASAP7_75t_L g4345 ( 
.A(n_4142),
.Y(n_4345)
);

BUFx2_ASAP7_75t_SL g4346 ( 
.A(n_3839),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_3783),
.Y(n_4347)
);

BUFx2_ASAP7_75t_SL g4348 ( 
.A(n_3702),
.Y(n_4348)
);

INVx6_ASAP7_75t_L g4349 ( 
.A(n_3704),
.Y(n_4349)
);

BUFx6f_ASAP7_75t_SL g4350 ( 
.A(n_3936),
.Y(n_4350)
);

BUFx12f_ASAP7_75t_L g4351 ( 
.A(n_4073),
.Y(n_4351)
);

NAND2x1p5_ASAP7_75t_L g4352 ( 
.A(n_3797),
.B(n_538),
.Y(n_4352)
);

BUFx4f_ASAP7_75t_SL g4353 ( 
.A(n_3682),
.Y(n_4353)
);

BUFx4f_ASAP7_75t_L g4354 ( 
.A(n_4056),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_3956),
.B(n_539),
.Y(n_4355)
);

BUFx4f_ASAP7_75t_L g4356 ( 
.A(n_4005),
.Y(n_4356)
);

INVx6_ASAP7_75t_L g4357 ( 
.A(n_4007),
.Y(n_4357)
);

BUFx3_ASAP7_75t_L g4358 ( 
.A(n_3675),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_3784),
.Y(n_4359)
);

CKINVDCx20_ASAP7_75t_R g4360 ( 
.A(n_3781),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_3818),
.Y(n_4361)
);

CKINVDCx6p67_ASAP7_75t_R g4362 ( 
.A(n_3837),
.Y(n_4362)
);

INVx1_ASAP7_75t_SL g4363 ( 
.A(n_3686),
.Y(n_4363)
);

INVx2_ASAP7_75t_L g4364 ( 
.A(n_4021),
.Y(n_4364)
);

BUFx12f_ASAP7_75t_L g4365 ( 
.A(n_4119),
.Y(n_4365)
);

INVx3_ASAP7_75t_L g4366 ( 
.A(n_4007),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4091),
.Y(n_4367)
);

NOR2xp33_ASAP7_75t_L g4368 ( 
.A(n_3712),
.B(n_539),
.Y(n_4368)
);

BUFx6f_ASAP7_75t_L g4369 ( 
.A(n_4007),
.Y(n_4369)
);

BUFx3_ASAP7_75t_L g4370 ( 
.A(n_3966),
.Y(n_4370)
);

BUFx2_ASAP7_75t_L g4371 ( 
.A(n_3964),
.Y(n_4371)
);

NAND2x1p5_ASAP7_75t_L g4372 ( 
.A(n_3798),
.B(n_539),
.Y(n_4372)
);

INVx3_ASAP7_75t_L g4373 ( 
.A(n_3967),
.Y(n_4373)
);

INVxp67_ASAP7_75t_SL g4374 ( 
.A(n_4041),
.Y(n_4374)
);

INVx5_ASAP7_75t_L g4375 ( 
.A(n_4123),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_3963),
.B(n_540),
.Y(n_4376)
);

INVx5_ASAP7_75t_L g4377 ( 
.A(n_4123),
.Y(n_4377)
);

INVxp67_ASAP7_75t_SL g4378 ( 
.A(n_4049),
.Y(n_4378)
);

CKINVDCx16_ASAP7_75t_R g4379 ( 
.A(n_4001),
.Y(n_4379)
);

BUFx8_ASAP7_75t_L g4380 ( 
.A(n_3969),
.Y(n_4380)
);

AOI22xp33_ASAP7_75t_L g4381 ( 
.A1(n_4141),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_4381)
);

BUFx3_ASAP7_75t_L g4382 ( 
.A(n_3991),
.Y(n_4382)
);

INVxp67_ASAP7_75t_SL g4383 ( 
.A(n_4063),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4076),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_3965),
.B(n_541),
.Y(n_4385)
);

INVx6_ASAP7_75t_L g4386 ( 
.A(n_4089),
.Y(n_4386)
);

INVx1_ASAP7_75t_SL g4387 ( 
.A(n_3880),
.Y(n_4387)
);

CKINVDCx20_ASAP7_75t_R g4388 ( 
.A(n_3750),
.Y(n_4388)
);

BUFx12f_ASAP7_75t_L g4389 ( 
.A(n_4035),
.Y(n_4389)
);

INVx1_ASAP7_75t_SL g4390 ( 
.A(n_3975),
.Y(n_4390)
);

BUFx2_ASAP7_75t_SL g4391 ( 
.A(n_3717),
.Y(n_4391)
);

BUFx12f_ASAP7_75t_L g4392 ( 
.A(n_4123),
.Y(n_4392)
);

INVx1_ASAP7_75t_SL g4393 ( 
.A(n_3920),
.Y(n_4393)
);

CKINVDCx20_ASAP7_75t_R g4394 ( 
.A(n_3731),
.Y(n_4394)
);

INVx4_ASAP7_75t_L g4395 ( 
.A(n_3950),
.Y(n_4395)
);

BUFx3_ASAP7_75t_L g4396 ( 
.A(n_3928),
.Y(n_4396)
);

NAND2xp5_ASAP7_75t_L g4397 ( 
.A(n_3999),
.B(n_541),
.Y(n_4397)
);

AND2x2_ASAP7_75t_L g4398 ( 
.A(n_4028),
.B(n_542),
.Y(n_4398)
);

BUFx3_ASAP7_75t_L g4399 ( 
.A(n_3861),
.Y(n_4399)
);

BUFx3_ASAP7_75t_L g4400 ( 
.A(n_3926),
.Y(n_4400)
);

NAND2x1p5_ASAP7_75t_L g4401 ( 
.A(n_3771),
.B(n_542),
.Y(n_4401)
);

INVx3_ASAP7_75t_L g4402 ( 
.A(n_4071),
.Y(n_4402)
);

INVx6_ASAP7_75t_SL g4403 ( 
.A(n_3976),
.Y(n_4403)
);

AOI22xp5_ASAP7_75t_L g4404 ( 
.A1(n_3696),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_4404)
);

CKINVDCx16_ASAP7_75t_R g4405 ( 
.A(n_3993),
.Y(n_4405)
);

BUFx4_ASAP7_75t_SL g4406 ( 
.A(n_4058),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_3823),
.Y(n_4407)
);

BUFx4_ASAP7_75t_SL g4408 ( 
.A(n_4083),
.Y(n_4408)
);

INVx5_ASAP7_75t_L g4409 ( 
.A(n_4010),
.Y(n_4409)
);

INVx1_ASAP7_75t_SL g4410 ( 
.A(n_4148),
.Y(n_4410)
);

INVx5_ASAP7_75t_L g4411 ( 
.A(n_4117),
.Y(n_4411)
);

BUFx6f_ASAP7_75t_L g4412 ( 
.A(n_4117),
.Y(n_4412)
);

INVx3_ASAP7_75t_L g4413 ( 
.A(n_3725),
.Y(n_4413)
);

NAND2x1p5_ASAP7_75t_L g4414 ( 
.A(n_3824),
.B(n_544),
.Y(n_4414)
);

AND2x2_ASAP7_75t_L g4415 ( 
.A(n_4054),
.B(n_546),
.Y(n_4415)
);

BUFx6f_ASAP7_75t_L g4416 ( 
.A(n_3715),
.Y(n_4416)
);

BUFx6f_ASAP7_75t_L g4417 ( 
.A(n_4088),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_3844),
.Y(n_4418)
);

INVx2_ASAP7_75t_SL g4419 ( 
.A(n_3865),
.Y(n_4419)
);

BUFx6f_ASAP7_75t_L g4420 ( 
.A(n_3860),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_3856),
.Y(n_4421)
);

INVx4_ASAP7_75t_L g4422 ( 
.A(n_3850),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_3858),
.Y(n_4423)
);

BUFx3_ASAP7_75t_L g4424 ( 
.A(n_3859),
.Y(n_4424)
);

BUFx2_ASAP7_75t_SL g4425 ( 
.A(n_3728),
.Y(n_4425)
);

NAND2x1p5_ASAP7_75t_L g4426 ( 
.A(n_3756),
.B(n_547),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_3680),
.Y(n_4427)
);

INVx5_ASAP7_75t_L g4428 ( 
.A(n_4077),
.Y(n_4428)
);

BUFx3_ASAP7_75t_L g4429 ( 
.A(n_4147),
.Y(n_4429)
);

BUFx6f_ASAP7_75t_L g4430 ( 
.A(n_4107),
.Y(n_4430)
);

BUFx12f_ASAP7_75t_L g4431 ( 
.A(n_3758),
.Y(n_4431)
);

INVx3_ASAP7_75t_L g4432 ( 
.A(n_4075),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_3888),
.Y(n_4433)
);

INVx2_ASAP7_75t_L g4434 ( 
.A(n_3896),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_3902),
.Y(n_4435)
);

BUFx3_ASAP7_75t_L g4436 ( 
.A(n_3747),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4121),
.Y(n_4437)
);

INVx6_ASAP7_75t_L g4438 ( 
.A(n_3746),
.Y(n_4438)
);

INVx2_ASAP7_75t_L g4439 ( 
.A(n_4121),
.Y(n_4439)
);

BUFx12f_ASAP7_75t_L g4440 ( 
.A(n_3775),
.Y(n_4440)
);

INVx3_ASAP7_75t_SL g4441 ( 
.A(n_4006),
.Y(n_4441)
);

BUFx6f_ASAP7_75t_L g4442 ( 
.A(n_3869),
.Y(n_4442)
);

INVx4_ASAP7_75t_L g4443 ( 
.A(n_4124),
.Y(n_4443)
);

BUFx3_ASAP7_75t_L g4444 ( 
.A(n_3945),
.Y(n_4444)
);

INVx3_ASAP7_75t_SL g4445 ( 
.A(n_4015),
.Y(n_4445)
);

CKINVDCx16_ASAP7_75t_R g4446 ( 
.A(n_3807),
.Y(n_4446)
);

BUFx6f_ASAP7_75t_L g4447 ( 
.A(n_3948),
.Y(n_4447)
);

AOI22xp33_ASAP7_75t_L g4448 ( 
.A1(n_3889),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.Y(n_4448)
);

NAND2x1p5_ASAP7_75t_L g4449 ( 
.A(n_4031),
.B(n_548),
.Y(n_4449)
);

OR2x2_ASAP7_75t_L g4450 ( 
.A(n_4036),
.B(n_548),
.Y(n_4450)
);

AND2x2_ASAP7_75t_L g4451 ( 
.A(n_4067),
.B(n_549),
.Y(n_4451)
);

BUFx3_ASAP7_75t_L g4452 ( 
.A(n_3918),
.Y(n_4452)
);

INVx2_ASAP7_75t_SL g4453 ( 
.A(n_3790),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_3921),
.B(n_549),
.Y(n_4454)
);

HB1xp67_ASAP7_75t_L g4455 ( 
.A(n_4102),
.Y(n_4455)
);

BUFx3_ASAP7_75t_L g4456 ( 
.A(n_3980),
.Y(n_4456)
);

AOI22xp33_ASAP7_75t_L g4457 ( 
.A1(n_3904),
.A2(n_3925),
.B1(n_3724),
.B2(n_3730),
.Y(n_4457)
);

INVx2_ASAP7_75t_SL g4458 ( 
.A(n_3793),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4092),
.B(n_550),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_L g4460 ( 
.A(n_4002),
.B(n_550),
.Y(n_4460)
);

AND2x4_ASAP7_75t_L g4461 ( 
.A(n_3754),
.B(n_552),
.Y(n_4461)
);

BUFx2_ASAP7_75t_L g4462 ( 
.A(n_3669),
.Y(n_4462)
);

BUFx2_ASAP7_75t_SL g4463 ( 
.A(n_3741),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_3933),
.Y(n_4464)
);

INVx5_ASAP7_75t_L g4465 ( 
.A(n_4130),
.Y(n_4465)
);

INVx2_ASAP7_75t_L g4466 ( 
.A(n_4030),
.Y(n_4466)
);

AO21x1_ASAP7_75t_L g4467 ( 
.A1(n_4018),
.A2(n_3895),
.B(n_3941),
.Y(n_4467)
);

AOI22xp33_ASAP7_75t_L g4468 ( 
.A1(n_4097),
.A2(n_553),
.B1(n_551),
.B2(n_552),
.Y(n_4468)
);

CKINVDCx20_ASAP7_75t_R g4469 ( 
.A(n_3979),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_4065),
.B(n_4012),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_3952),
.Y(n_4471)
);

INVx4_ASAP7_75t_L g4472 ( 
.A(n_4057),
.Y(n_4472)
);

BUFx8_ASAP7_75t_L g4473 ( 
.A(n_4078),
.Y(n_4473)
);

BUFx2_ASAP7_75t_L g4474 ( 
.A(n_4000),
.Y(n_4474)
);

INVx3_ASAP7_75t_L g4475 ( 
.A(n_4143),
.Y(n_4475)
);

BUFx3_ASAP7_75t_L g4476 ( 
.A(n_3987),
.Y(n_4476)
);

OR2x2_ASAP7_75t_L g4477 ( 
.A(n_3970),
.B(n_551),
.Y(n_4477)
);

CKINVDCx8_ASAP7_75t_R g4478 ( 
.A(n_4094),
.Y(n_4478)
);

BUFx6f_ASAP7_75t_L g4479 ( 
.A(n_4134),
.Y(n_4479)
);

INVx1_ASAP7_75t_SL g4480 ( 
.A(n_3742),
.Y(n_4480)
);

BUFx3_ASAP7_75t_L g4481 ( 
.A(n_3990),
.Y(n_4481)
);

BUFx3_ASAP7_75t_L g4482 ( 
.A(n_3851),
.Y(n_4482)
);

CKINVDCx14_ASAP7_75t_R g4483 ( 
.A(n_3878),
.Y(n_4483)
);

AND2x2_ASAP7_75t_L g4484 ( 
.A(n_4101),
.B(n_551),
.Y(n_4484)
);

OR2x2_ASAP7_75t_L g4485 ( 
.A(n_3958),
.B(n_552),
.Y(n_4485)
);

CKINVDCx20_ASAP7_75t_R g4486 ( 
.A(n_3914),
.Y(n_4486)
);

BUFx3_ASAP7_75t_L g4487 ( 
.A(n_3852),
.Y(n_4487)
);

BUFx6f_ASAP7_75t_SL g4488 ( 
.A(n_4111),
.Y(n_4488)
);

INVx4_ASAP7_75t_L g4489 ( 
.A(n_4110),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_3984),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4014),
.Y(n_4491)
);

INVx1_ASAP7_75t_SL g4492 ( 
.A(n_3862),
.Y(n_4492)
);

AOI22xp5_ASAP7_75t_L g4493 ( 
.A1(n_3881),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.Y(n_4493)
);

BUFx6f_ASAP7_75t_L g4494 ( 
.A(n_4115),
.Y(n_4494)
);

NAND2x1p5_ASAP7_75t_L g4495 ( 
.A(n_3946),
.B(n_555),
.Y(n_4495)
);

BUFx2_ASAP7_75t_L g4496 ( 
.A(n_4133),
.Y(n_4496)
);

BUFx2_ASAP7_75t_L g4497 ( 
.A(n_3943),
.Y(n_4497)
);

INVx3_ASAP7_75t_L g4498 ( 
.A(n_3863),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_3871),
.B(n_556),
.Y(n_4499)
);

NAND2x1p5_ASAP7_75t_L g4500 ( 
.A(n_3996),
.B(n_556),
.Y(n_4500)
);

BUFx5_ASAP7_75t_L g4501 ( 
.A(n_4114),
.Y(n_4501)
);

BUFx2_ASAP7_75t_L g4502 ( 
.A(n_3874),
.Y(n_4502)
);

BUFx3_ASAP7_75t_L g4503 ( 
.A(n_3875),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_3930),
.B(n_4042),
.Y(n_4504)
);

BUFx3_ASAP7_75t_L g4505 ( 
.A(n_3883),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4016),
.Y(n_4506)
);

BUFx3_ASAP7_75t_L g4507 ( 
.A(n_3947),
.Y(n_4507)
);

BUFx3_ASAP7_75t_L g4508 ( 
.A(n_3954),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4019),
.Y(n_4509)
);

INVx3_ASAP7_75t_SL g4510 ( 
.A(n_3825),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_4118),
.Y(n_4511)
);

AND2x2_ASAP7_75t_L g4512 ( 
.A(n_4116),
.B(n_556),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4032),
.Y(n_4513)
);

INVx4_ASAP7_75t_L g4514 ( 
.A(n_4128),
.Y(n_4514)
);

NAND2x1p5_ASAP7_75t_L g4515 ( 
.A(n_3740),
.B(n_557),
.Y(n_4515)
);

BUFx6f_ASAP7_75t_L g4516 ( 
.A(n_4120),
.Y(n_4516)
);

INVx2_ASAP7_75t_SL g4517 ( 
.A(n_3903),
.Y(n_4517)
);

INVx3_ASAP7_75t_L g4518 ( 
.A(n_4085),
.Y(n_4518)
);

CKINVDCx5p33_ASAP7_75t_R g4519 ( 
.A(n_3906),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4048),
.B(n_557),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4039),
.Y(n_4521)
);

BUFx12f_ASAP7_75t_L g4522 ( 
.A(n_3733),
.Y(n_4522)
);

INVx3_ASAP7_75t_L g4523 ( 
.A(n_4086),
.Y(n_4523)
);

INVx5_ASAP7_75t_L g4524 ( 
.A(n_3736),
.Y(n_4524)
);

HB1xp67_ASAP7_75t_L g4525 ( 
.A(n_3940),
.Y(n_4525)
);

INVx1_ASAP7_75t_SL g4526 ( 
.A(n_4044),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_4069),
.B(n_557),
.Y(n_4527)
);

INVx2_ASAP7_75t_L g4528 ( 
.A(n_3972),
.Y(n_4528)
);

AND2x2_ASAP7_75t_L g4529 ( 
.A(n_3891),
.B(n_558),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4047),
.Y(n_4530)
);

BUFx6f_ASAP7_75t_L g4531 ( 
.A(n_4095),
.Y(n_4531)
);

AND2x4_ASAP7_75t_L g4532 ( 
.A(n_3745),
.B(n_559),
.Y(n_4532)
);

CKINVDCx5p33_ASAP7_75t_R g4533 ( 
.A(n_3978),
.Y(n_4533)
);

BUFx6f_ASAP7_75t_L g4534 ( 
.A(n_4099),
.Y(n_4534)
);

BUFx6f_ASAP7_75t_L g4535 ( 
.A(n_4050),
.Y(n_4535)
);

AND2x2_ASAP7_75t_L g4536 ( 
.A(n_4004),
.B(n_558),
.Y(n_4536)
);

CKINVDCx20_ASAP7_75t_R g4537 ( 
.A(n_4025),
.Y(n_4537)
);

BUFx2_ASAP7_75t_SL g4538 ( 
.A(n_3800),
.Y(n_4538)
);

CKINVDCx20_ASAP7_75t_R g4539 ( 
.A(n_3857),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4060),
.Y(n_4540)
);

BUFx2_ASAP7_75t_R g4541 ( 
.A(n_4068),
.Y(n_4541)
);

BUFx3_ASAP7_75t_L g4542 ( 
.A(n_4070),
.Y(n_4542)
);

INVx3_ASAP7_75t_SL g4543 ( 
.A(n_4090),
.Y(n_4543)
);

INVx2_ASAP7_75t_SL g4544 ( 
.A(n_4087),
.Y(n_4544)
);

INVx2_ASAP7_75t_SL g4545 ( 
.A(n_4122),
.Y(n_4545)
);

BUFx6f_ASAP7_75t_L g4546 ( 
.A(n_4105),
.Y(n_4546)
);

INVx5_ASAP7_75t_L g4547 ( 
.A(n_3830),
.Y(n_4547)
);

BUFx3_ASAP7_75t_L g4548 ( 
.A(n_4084),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_3830),
.Y(n_4549)
);

BUFx3_ASAP7_75t_L g4550 ( 
.A(n_4081),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_L g4551 ( 
.A(n_4013),
.B(n_559),
.Y(n_4551)
);

INVx2_ASAP7_75t_L g4552 ( 
.A(n_4127),
.Y(n_4552)
);

BUFx6f_ASAP7_75t_L g4553 ( 
.A(n_4093),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_3935),
.Y(n_4554)
);

INVx2_ASAP7_75t_SL g4555 ( 
.A(n_3835),
.Y(n_4555)
);

BUFx6f_ASAP7_75t_L g4556 ( 
.A(n_4080),
.Y(n_4556)
);

AND2x4_ASAP7_75t_L g4557 ( 
.A(n_3811),
.B(n_561),
.Y(n_4557)
);

OAI22xp33_ASAP7_75t_L g4558 ( 
.A1(n_4342),
.A2(n_4405),
.B1(n_4219),
.B2(n_4207),
.Y(n_4558)
);

HB1xp67_ASAP7_75t_L g4559 ( 
.A(n_4309),
.Y(n_4559)
);

OAI22xp5_ASAP7_75t_L g4560 ( 
.A1(n_4483),
.A2(n_3804),
.B1(n_3931),
.B2(n_3960),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4427),
.B(n_3700),
.Y(n_4561)
);

INVx1_ASAP7_75t_SL g4562 ( 
.A(n_4406),
.Y(n_4562)
);

OAI22x1_ASAP7_75t_L g4563 ( 
.A1(n_4321),
.A2(n_3988),
.B1(n_4112),
.B2(n_4079),
.Y(n_4563)
);

INVx2_ASAP7_75t_L g4564 ( 
.A(n_4169),
.Y(n_4564)
);

OAI21x1_ASAP7_75t_L g4565 ( 
.A1(n_4433),
.A2(n_3718),
.B(n_3697),
.Y(n_4565)
);

OAI21x1_ASAP7_75t_L g4566 ( 
.A1(n_4434),
.A2(n_3719),
.B(n_3693),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_4330),
.B(n_3808),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_4337),
.B(n_3780),
.Y(n_4568)
);

AND2x4_ASAP7_75t_L g4569 ( 
.A(n_4214),
.B(n_4037),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4155),
.Y(n_4570)
);

AND2x2_ASAP7_75t_L g4571 ( 
.A(n_4367),
.B(n_4062),
.Y(n_4571)
);

OAI21x1_ASAP7_75t_L g4572 ( 
.A1(n_4466),
.A2(n_3672),
.B(n_3699),
.Y(n_4572)
);

AO21x2_ASAP7_75t_L g4573 ( 
.A1(n_4464),
.A2(n_3774),
.B(n_3801),
.Y(n_4573)
);

OAI21x1_ASAP7_75t_L g4574 ( 
.A1(n_4432),
.A2(n_3720),
.B(n_3986),
.Y(n_4574)
);

INVx2_ASAP7_75t_L g4575 ( 
.A(n_4175),
.Y(n_4575)
);

AO21x2_ASAP7_75t_L g4576 ( 
.A1(n_4415),
.A2(n_3968),
.B(n_3951),
.Y(n_4576)
);

BUFx6f_ASAP7_75t_L g4577 ( 
.A(n_4215),
.Y(n_4577)
);

INVx1_ASAP7_75t_SL g4578 ( 
.A(n_4408),
.Y(n_4578)
);

AND2x4_ASAP7_75t_L g4579 ( 
.A(n_4214),
.B(n_3855),
.Y(n_4579)
);

OAI22xp33_ASAP7_75t_L g4580 ( 
.A1(n_4219),
.A2(n_4074),
.B1(n_3955),
.B2(n_4034),
.Y(n_4580)
);

AND2x4_ASAP7_75t_L g4581 ( 
.A(n_4292),
.B(n_4301),
.Y(n_4581)
);

AOI221xp5_ASAP7_75t_L g4582 ( 
.A1(n_4457),
.A2(n_3843),
.B1(n_3813),
.B2(n_3809),
.C(n_3977),
.Y(n_4582)
);

BUFx3_ASAP7_75t_L g4583 ( 
.A(n_4172),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4159),
.Y(n_4584)
);

INVx3_ASAP7_75t_L g4585 ( 
.A(n_4217),
.Y(n_4585)
);

INVxp67_ASAP7_75t_L g4586 ( 
.A(n_4312),
.Y(n_4586)
);

OAI21xp5_ASAP7_75t_L g4587 ( 
.A1(n_4354),
.A2(n_3735),
.B(n_3905),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4161),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4546),
.B(n_4059),
.Y(n_4589)
);

OA21x2_ASAP7_75t_L g4590 ( 
.A1(n_4439),
.A2(n_4043),
.B(n_4138),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_4185),
.Y(n_4591)
);

BUFx12f_ASAP7_75t_L g4592 ( 
.A(n_4157),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4546),
.B(n_4552),
.Y(n_4593)
);

INVx2_ASAP7_75t_SL g4594 ( 
.A(n_4182),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_L g4595 ( 
.A(n_4259),
.B(n_3814),
.Y(n_4595)
);

OAI21x1_ASAP7_75t_L g4596 ( 
.A1(n_4413),
.A2(n_3872),
.B(n_3870),
.Y(n_4596)
);

OAI22xp5_ASAP7_75t_L g4597 ( 
.A1(n_4394),
.A2(n_3815),
.B1(n_3911),
.B2(n_4017),
.Y(n_4597)
);

OR2x6_ASAP7_75t_L g4598 ( 
.A(n_4345),
.B(n_3924),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4171),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_4200),
.Y(n_4600)
);

AOI22xp33_ASAP7_75t_SL g4601 ( 
.A1(n_4463),
.A2(n_4009),
.B1(n_4055),
.B2(n_4106),
.Y(n_4601)
);

AND2x4_ASAP7_75t_L g4602 ( 
.A(n_4184),
.B(n_4026),
.Y(n_4602)
);

NOR2xp67_ASAP7_75t_L g4603 ( 
.A(n_4149),
.B(n_560),
.Y(n_4603)
);

AOI222xp33_ASAP7_75t_L g4604 ( 
.A1(n_4356),
.A2(n_3974),
.B1(n_3992),
.B2(n_3836),
.C1(n_4135),
.C2(n_4132),
.Y(n_4604)
);

OAI21x1_ASAP7_75t_L g4605 ( 
.A1(n_4364),
.A2(n_3908),
.B(n_3879),
.Y(n_4605)
);

NOR2x1_ASAP7_75t_SL g4606 ( 
.A(n_4170),
.B(n_3770),
.Y(n_4606)
);

A2O1A1Ixp33_ASAP7_75t_L g4607 ( 
.A1(n_4345),
.A2(n_4145),
.B(n_3796),
.C(n_3799),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4178),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4189),
.Y(n_4609)
);

INVx4_ASAP7_75t_L g4610 ( 
.A(n_4211),
.Y(n_4610)
);

OA21x2_ASAP7_75t_L g4611 ( 
.A1(n_4329),
.A2(n_3981),
.B(n_3773),
.Y(n_4611)
);

OAI21x1_ASAP7_75t_L g4612 ( 
.A1(n_4347),
.A2(n_3917),
.B(n_3909),
.Y(n_4612)
);

NOR2xp33_ASAP7_75t_L g4613 ( 
.A(n_4336),
.B(n_562),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_L g4614 ( 
.A(n_4343),
.B(n_3989),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4198),
.Y(n_4615)
);

OAI21x1_ASAP7_75t_L g4616 ( 
.A1(n_4308),
.A2(n_3934),
.B(n_3922),
.Y(n_4616)
);

OAI21x1_ASAP7_75t_L g4617 ( 
.A1(n_4511),
.A2(n_3942),
.B(n_3939),
.Y(n_4617)
);

BUFx3_ASAP7_75t_L g4618 ( 
.A(n_4193),
.Y(n_4618)
);

NAND2x1p5_ASAP7_75t_L g4619 ( 
.A(n_4162),
.B(n_3822),
.Y(n_4619)
);

INVxp67_ASAP7_75t_L g4620 ( 
.A(n_4317),
.Y(n_4620)
);

OAI21x1_ASAP7_75t_SL g4621 ( 
.A1(n_4243),
.A2(n_3892),
.B(n_3962),
.Y(n_4621)
);

HB1xp67_ASAP7_75t_L g4622 ( 
.A(n_4245),
.Y(n_4622)
);

AOI221xp5_ASAP7_75t_L g4623 ( 
.A1(n_4368),
.A2(n_4109),
.B1(n_4104),
.B2(n_3816),
.C(n_4008),
.Y(n_4623)
);

NOR2xp67_ASAP7_75t_L g4624 ( 
.A(n_4151),
.B(n_4246),
.Y(n_4624)
);

INVx2_ASAP7_75t_L g4625 ( 
.A(n_4239),
.Y(n_4625)
);

OAI21x1_ASAP7_75t_L g4626 ( 
.A1(n_4515),
.A2(n_4027),
.B(n_3957),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4204),
.Y(n_4627)
);

OA21x2_ASAP7_75t_L g4628 ( 
.A1(n_4437),
.A2(n_4474),
.B(n_4496),
.Y(n_4628)
);

INVx3_ASAP7_75t_L g4629 ( 
.A(n_4183),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4455),
.B(n_563),
.Y(n_4630)
);

AND2x6_ASAP7_75t_L g4631 ( 
.A(n_4256),
.B(n_3915),
.Y(n_4631)
);

OAI21x1_ASAP7_75t_L g4632 ( 
.A1(n_4331),
.A2(n_4100),
.B(n_4096),
.Y(n_4632)
);

OAI21x1_ASAP7_75t_L g4633 ( 
.A1(n_4402),
.A2(n_4113),
.B(n_4108),
.Y(n_4633)
);

OA21x2_ASAP7_75t_L g4634 ( 
.A1(n_4467),
.A2(n_4022),
.B(n_4011),
.Y(n_4634)
);

NOR2xp33_ASAP7_75t_L g4635 ( 
.A(n_4290),
.B(n_563),
.Y(n_4635)
);

OAI21x1_ASAP7_75t_L g4636 ( 
.A1(n_4366),
.A2(n_4129),
.B(n_4126),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_4363),
.B(n_4190),
.Y(n_4637)
);

INVx2_ASAP7_75t_L g4638 ( 
.A(n_4293),
.Y(n_4638)
);

OR2x2_ASAP7_75t_L g4639 ( 
.A(n_4307),
.B(n_564),
.Y(n_4639)
);

OAI21x1_ASAP7_75t_L g4640 ( 
.A1(n_4467),
.A2(n_4137),
.B(n_4136),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4206),
.Y(n_4641)
);

NOR2xp67_ASAP7_75t_L g4642 ( 
.A(n_4246),
.B(n_564),
.Y(n_4642)
);

OAI21x1_ASAP7_75t_L g4643 ( 
.A1(n_4500),
.A2(n_4051),
.B(n_4045),
.Y(n_4643)
);

OAI21x1_ASAP7_75t_L g4644 ( 
.A1(n_4528),
.A2(n_4061),
.B(n_4052),
.Y(n_4644)
);

AND2x2_ASAP7_75t_L g4645 ( 
.A(n_4190),
.B(n_565),
.Y(n_4645)
);

AO21x2_ASAP7_75t_L g4646 ( 
.A1(n_4551),
.A2(n_3971),
.B(n_3961),
.Y(n_4646)
);

OA21x2_ASAP7_75t_L g4647 ( 
.A1(n_4549),
.A2(n_4023),
.B(n_4125),
.Y(n_4647)
);

NAND2x1p5_ASAP7_75t_L g4648 ( 
.A(n_4240),
.B(n_565),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4210),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4384),
.B(n_4098),
.Y(n_4650)
);

AOI21xp5_ASAP7_75t_L g4651 ( 
.A1(n_4480),
.A2(n_3994),
.B(n_4053),
.Y(n_4651)
);

OAI21x1_ASAP7_75t_L g4652 ( 
.A1(n_4233),
.A2(n_4082),
.B(n_4103),
.Y(n_4652)
);

OA21x2_ASAP7_75t_L g4653 ( 
.A1(n_4462),
.A2(n_4131),
.B(n_565),
.Y(n_4653)
);

OAI21xp5_ASAP7_75t_L g4654 ( 
.A1(n_4194),
.A2(n_566),
.B(n_567),
.Y(n_4654)
);

AND2x2_ASAP7_75t_L g4655 ( 
.A(n_4550),
.B(n_567),
.Y(n_4655)
);

AOI21xp5_ASAP7_75t_L g4656 ( 
.A1(n_4375),
.A2(n_568),
.B(n_569),
.Y(n_4656)
);

AOI21x1_ASAP7_75t_L g4657 ( 
.A1(n_4264),
.A2(n_4191),
.B(n_4462),
.Y(n_4657)
);

INVx3_ASAP7_75t_L g4658 ( 
.A(n_4211),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_L g4659 ( 
.A(n_4322),
.B(n_570),
.Y(n_4659)
);

INVx2_ASAP7_75t_L g4660 ( 
.A(n_4297),
.Y(n_4660)
);

INVx2_ASAP7_75t_L g4661 ( 
.A(n_4300),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4230),
.Y(n_4662)
);

OAI21x1_ASAP7_75t_L g4663 ( 
.A1(n_4373),
.A2(n_752),
.B(n_751),
.Y(n_4663)
);

CKINVDCx6p67_ASAP7_75t_R g4664 ( 
.A(n_4181),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4234),
.Y(n_4665)
);

INVx3_ASAP7_75t_L g4666 ( 
.A(n_4305),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_4258),
.Y(n_4667)
);

OAI21x1_ASAP7_75t_L g4668 ( 
.A1(n_4518),
.A2(n_754),
.B(n_753),
.Y(n_4668)
);

OAI222xp33_ASAP7_75t_L g4669 ( 
.A1(n_4237),
.A2(n_572),
.B1(n_574),
.B2(n_570),
.C1(n_571),
.C2(n_573),
.Y(n_4669)
);

OR2x6_ASAP7_75t_L g4670 ( 
.A(n_4174),
.B(n_571),
.Y(n_4670)
);

OAI21x1_ASAP7_75t_L g4671 ( 
.A1(n_4523),
.A2(n_756),
.B(n_755),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4278),
.Y(n_4672)
);

OR2x6_ASAP7_75t_SL g4673 ( 
.A(n_4272),
.B(n_4403),
.Y(n_4673)
);

NAND2x1p5_ASAP7_75t_L g4674 ( 
.A(n_4203),
.B(n_572),
.Y(n_4674)
);

INVx2_ASAP7_75t_SL g4675 ( 
.A(n_4182),
.Y(n_4675)
);

BUFx6f_ASAP7_75t_L g4676 ( 
.A(n_4323),
.Y(n_4676)
);

NOR2xp67_ASAP7_75t_L g4677 ( 
.A(n_4252),
.B(n_572),
.Y(n_4677)
);

AO31x2_ASAP7_75t_L g4678 ( 
.A1(n_4472),
.A2(n_575),
.A3(n_573),
.B(n_574),
.Y(n_4678)
);

O2A1O1Ixp33_ASAP7_75t_L g4679 ( 
.A1(n_4237),
.A2(n_577),
.B(n_575),
.C(n_576),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4288),
.Y(n_4680)
);

NAND2x1p5_ASAP7_75t_L g4681 ( 
.A(n_4187),
.B(n_577),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4268),
.Y(n_4682)
);

AND2x4_ASAP7_75t_L g4683 ( 
.A(n_4375),
.B(n_577),
.Y(n_4683)
);

OAI22xp5_ASAP7_75t_L g4684 ( 
.A1(n_4539),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_4684)
);

OAI21x1_ASAP7_75t_L g4685 ( 
.A1(n_4249),
.A2(n_759),
.B(n_758),
.Y(n_4685)
);

INVx2_ASAP7_75t_L g4686 ( 
.A(n_4289),
.Y(n_4686)
);

AO21x2_ASAP7_75t_L g4687 ( 
.A1(n_4225),
.A2(n_4271),
.B(n_4238),
.Y(n_4687)
);

OAI21x1_ASAP7_75t_L g4688 ( 
.A1(n_4435),
.A2(n_761),
.B(n_760),
.Y(n_4688)
);

INVx1_ASAP7_75t_SL g4689 ( 
.A(n_4316),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_SL g4690 ( 
.A(n_4377),
.B(n_4379),
.Y(n_4690)
);

HB1xp67_ASAP7_75t_L g4691 ( 
.A(n_4344),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4277),
.Y(n_4692)
);

NAND2x1p5_ASAP7_75t_L g4693 ( 
.A(n_4164),
.B(n_578),
.Y(n_4693)
);

OAI22xp33_ASAP7_75t_L g4694 ( 
.A1(n_4392),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_4694)
);

AO31x2_ASAP7_75t_L g4695 ( 
.A1(n_4443),
.A2(n_582),
.A3(n_579),
.B(n_581),
.Y(n_4695)
);

BUFx6f_ASAP7_75t_L g4696 ( 
.A(n_4216),
.Y(n_4696)
);

NAND2xp5_ASAP7_75t_L g4697 ( 
.A(n_4315),
.B(n_581),
.Y(n_4697)
);

INVx4_ASAP7_75t_L g4698 ( 
.A(n_4202),
.Y(n_4698)
);

AOI221xp5_ASAP7_75t_L g4699 ( 
.A1(n_4236),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.C(n_584),
.Y(n_4699)
);

OR2x2_ASAP7_75t_L g4700 ( 
.A(n_4325),
.B(n_582),
.Y(n_4700)
);

OAI21xp5_ASAP7_75t_L g4701 ( 
.A1(n_4532),
.A2(n_4426),
.B(n_4536),
.Y(n_4701)
);

OAI21x1_ASAP7_75t_L g4702 ( 
.A1(n_4319),
.A2(n_4451),
.B(n_4459),
.Y(n_4702)
);

AND2x4_ASAP7_75t_L g4703 ( 
.A(n_4377),
.B(n_583),
.Y(n_4703)
);

NAND2xp5_ASAP7_75t_SL g4704 ( 
.A(n_4524),
.B(n_583),
.Y(n_4704)
);

BUFx2_ASAP7_75t_L g4705 ( 
.A(n_4365),
.Y(n_4705)
);

OAI21x1_ASAP7_75t_L g4706 ( 
.A1(n_4451),
.A2(n_762),
.B(n_761),
.Y(n_4706)
);

AO31x2_ASAP7_75t_L g4707 ( 
.A1(n_4489),
.A2(n_587),
.A3(n_585),
.B(n_586),
.Y(n_4707)
);

INVx1_ASAP7_75t_SL g4708 ( 
.A(n_4188),
.Y(n_4708)
);

INVx2_ASAP7_75t_L g4709 ( 
.A(n_4295),
.Y(n_4709)
);

OA21x2_ASAP7_75t_L g4710 ( 
.A1(n_4371),
.A2(n_585),
.B(n_587),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4374),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4378),
.B(n_4383),
.Y(n_4712)
);

BUFx2_ASAP7_75t_L g4713 ( 
.A(n_4242),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4160),
.Y(n_4714)
);

INVx2_ASAP7_75t_L g4715 ( 
.A(n_4303),
.Y(n_4715)
);

NOR2xp67_ASAP7_75t_L g4716 ( 
.A(n_4252),
.B(n_588),
.Y(n_4716)
);

AO32x2_ASAP7_75t_L g4717 ( 
.A1(n_4299),
.A2(n_591),
.A3(n_589),
.B1(n_590),
.B2(n_592),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4355),
.B(n_589),
.Y(n_4718)
);

AND2x6_ASAP7_75t_L g4719 ( 
.A(n_4256),
.B(n_590),
.Y(n_4719)
);

OAI21x1_ASAP7_75t_L g4720 ( 
.A1(n_4459),
.A2(n_765),
.B(n_762),
.Y(n_4720)
);

OAI222xp33_ASAP7_75t_L g4721 ( 
.A1(n_4422),
.A2(n_595),
.B1(n_597),
.B2(n_591),
.C1(n_594),
.C2(n_596),
.Y(n_4721)
);

AND2x4_ASAP7_75t_L g4722 ( 
.A(n_4266),
.B(n_594),
.Y(n_4722)
);

OAI22xp5_ASAP7_75t_L g4723 ( 
.A1(n_4195),
.A2(n_597),
.B1(n_594),
.B2(n_596),
.Y(n_4723)
);

INVx4_ASAP7_75t_L g4724 ( 
.A(n_4208),
.Y(n_4724)
);

INVx2_ASAP7_75t_L g4725 ( 
.A(n_4370),
.Y(n_4725)
);

INVx2_ASAP7_75t_L g4726 ( 
.A(n_4382),
.Y(n_4726)
);

OAI21x1_ASAP7_75t_L g4727 ( 
.A1(n_4484),
.A2(n_766),
.B(n_765),
.Y(n_4727)
);

OAI22xp33_ASAP7_75t_L g4728 ( 
.A1(n_4510),
.A2(n_598),
.B1(n_596),
.B2(n_597),
.Y(n_4728)
);

INVx2_ASAP7_75t_L g4729 ( 
.A(n_4284),
.Y(n_4729)
);

OR2x2_ASAP7_75t_L g4730 ( 
.A(n_4393),
.B(n_598),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_4226),
.Y(n_4731)
);

INVx6_ASAP7_75t_L g4732 ( 
.A(n_4199),
.Y(n_4732)
);

INVx1_ASAP7_75t_L g4733 ( 
.A(n_4205),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_4212),
.Y(n_4734)
);

INVx2_ASAP7_75t_SL g4735 ( 
.A(n_4216),
.Y(n_4735)
);

O2A1O1Ixp33_ASAP7_75t_SL g4736 ( 
.A1(n_4254),
.A2(n_600),
.B(n_598),
.C(n_599),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4221),
.Y(n_4737)
);

OA21x2_ASAP7_75t_L g4738 ( 
.A1(n_4166),
.A2(n_599),
.B(n_601),
.Y(n_4738)
);

HB1xp67_ASAP7_75t_L g4739 ( 
.A(n_4430),
.Y(n_4739)
);

AO21x2_ASAP7_75t_L g4740 ( 
.A1(n_4536),
.A2(n_599),
.B(n_601),
.Y(n_4740)
);

NOR2x1_ASAP7_75t_SL g4741 ( 
.A(n_4228),
.B(n_601),
.Y(n_4741)
);

OAI22xp5_ASAP7_75t_L g4742 ( 
.A1(n_4195),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.Y(n_4742)
);

OAI21x1_ASAP7_75t_L g4743 ( 
.A1(n_4512),
.A2(n_768),
.B(n_767),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4450),
.Y(n_4744)
);

OAI21x1_ASAP7_75t_L g4745 ( 
.A1(n_4311),
.A2(n_770),
.B(n_769),
.Y(n_4745)
);

INVx2_ASAP7_75t_L g4746 ( 
.A(n_4275),
.Y(n_4746)
);

INVx2_ASAP7_75t_SL g4747 ( 
.A(n_4150),
.Y(n_4747)
);

OAI21x1_ASAP7_75t_L g4748 ( 
.A1(n_4449),
.A2(n_771),
.B(n_769),
.Y(n_4748)
);

INVx6_ASAP7_75t_L g4749 ( 
.A(n_4150),
.Y(n_4749)
);

OAI22xp5_ASAP7_75t_L g4750 ( 
.A1(n_4362),
.A2(n_4446),
.B1(n_4388),
.B2(n_4285),
.Y(n_4750)
);

OA21x2_ASAP7_75t_L g4751 ( 
.A1(n_4166),
.A2(n_602),
.B(n_603),
.Y(n_4751)
);

INVx2_ASAP7_75t_L g4752 ( 
.A(n_4275),
.Y(n_4752)
);

BUFx6f_ASAP7_75t_L g4753 ( 
.A(n_4223),
.Y(n_4753)
);

BUFx2_ASAP7_75t_L g4754 ( 
.A(n_4351),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4450),
.Y(n_4755)
);

NOR2xp67_ASAP7_75t_L g4756 ( 
.A(n_4196),
.B(n_603),
.Y(n_4756)
);

INVx2_ASAP7_75t_L g4757 ( 
.A(n_4553),
.Y(n_4757)
);

AO31x2_ASAP7_75t_L g4758 ( 
.A1(n_4514),
.A2(n_606),
.A3(n_604),
.B(n_605),
.Y(n_4758)
);

AOI221x1_ASAP7_75t_L g4759 ( 
.A1(n_4163),
.A2(n_775),
.B1(n_776),
.B2(n_773),
.C(n_771),
.Y(n_4759)
);

AOI22xp5_ASAP7_75t_L g4760 ( 
.A1(n_4537),
.A2(n_607),
.B1(n_605),
.B2(n_606),
.Y(n_4760)
);

O2A1O1Ixp33_ASAP7_75t_SL g4761 ( 
.A1(n_4177),
.A2(n_609),
.B(n_607),
.C(n_608),
.Y(n_4761)
);

NOR2xp33_ASAP7_75t_L g4762 ( 
.A(n_4353),
.B(n_608),
.Y(n_4762)
);

OR2x6_ASAP7_75t_L g4763 ( 
.A(n_4248),
.B(n_609),
.Y(n_4763)
);

INVx2_ASAP7_75t_L g4764 ( 
.A(n_4553),
.Y(n_4764)
);

AND2x4_ASAP7_75t_L g4765 ( 
.A(n_4270),
.B(n_610),
.Y(n_4765)
);

INVx1_ASAP7_75t_SL g4766 ( 
.A(n_4165),
.Y(n_4766)
);

AOI221xp5_ASAP7_75t_L g4767 ( 
.A1(n_4420),
.A2(n_614),
.B1(n_611),
.B2(n_612),
.C(n_615),
.Y(n_4767)
);

BUFx2_ASAP7_75t_L g4768 ( 
.A(n_4276),
.Y(n_4768)
);

NOR2xp33_ASAP7_75t_L g4769 ( 
.A(n_4470),
.B(n_611),
.Y(n_4769)
);

OAI21x1_ASAP7_75t_L g4770 ( 
.A1(n_4341),
.A2(n_777),
.B(n_775),
.Y(n_4770)
);

AOI22xp33_ASAP7_75t_SL g4771 ( 
.A1(n_4348),
.A2(n_615),
.B1(n_612),
.B2(n_614),
.Y(n_4771)
);

OAI21xp5_ASAP7_75t_L g4772 ( 
.A1(n_4493),
.A2(n_4404),
.B(n_4529),
.Y(n_4772)
);

AOI22x1_ASAP7_75t_L g4773 ( 
.A1(n_4168),
.A2(n_616),
.B1(n_612),
.B2(n_615),
.Y(n_4773)
);

O2A1O1Ixp33_ASAP7_75t_L g4774 ( 
.A1(n_4419),
.A2(n_618),
.B(n_616),
.C(n_617),
.Y(n_4774)
);

INVx2_ASAP7_75t_L g4775 ( 
.A(n_4257),
.Y(n_4775)
);

AO21x2_ASAP7_75t_L g4776 ( 
.A1(n_4529),
.A2(n_618),
.B(n_619),
.Y(n_4776)
);

AO21x2_ASAP7_75t_L g4777 ( 
.A1(n_4279),
.A2(n_620),
.B(n_621),
.Y(n_4777)
);

OA21x2_ASAP7_75t_L g4778 ( 
.A1(n_4251),
.A2(n_620),
.B(n_621),
.Y(n_4778)
);

INVx2_ASAP7_75t_L g4779 ( 
.A(n_4334),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4298),
.Y(n_4780)
);

HB1xp67_ASAP7_75t_L g4781 ( 
.A(n_4291),
.Y(n_4781)
);

OR2x2_ASAP7_75t_L g4782 ( 
.A(n_4424),
.B(n_622),
.Y(n_4782)
);

BUFx2_ASAP7_75t_SL g4783 ( 
.A(n_4213),
.Y(n_4783)
);

NOR2x1_ASAP7_75t_SL g4784 ( 
.A(n_4253),
.B(n_622),
.Y(n_4784)
);

OAI21x1_ASAP7_75t_L g4785 ( 
.A1(n_4232),
.A2(n_779),
.B(n_778),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4298),
.Y(n_4786)
);

NOR2xp67_ASAP7_75t_L g4787 ( 
.A(n_4409),
.B(n_623),
.Y(n_4787)
);

AO31x2_ASAP7_75t_L g4788 ( 
.A1(n_4324),
.A2(n_625),
.A3(n_623),
.B(n_624),
.Y(n_4788)
);

INVx2_ASAP7_75t_L g4789 ( 
.A(n_4479),
.Y(n_4789)
);

AOI21xp5_ASAP7_75t_L g4790 ( 
.A1(n_4410),
.A2(n_626),
.B(n_627),
.Y(n_4790)
);

OAI22xp5_ASAP7_75t_L g4791 ( 
.A1(n_4338),
.A2(n_628),
.B1(n_626),
.B2(n_627),
.Y(n_4791)
);

AOI221xp5_ASAP7_75t_L g4792 ( 
.A1(n_4420),
.A2(n_630),
.B1(n_628),
.B2(n_629),
.C(n_631),
.Y(n_4792)
);

AND2x4_ASAP7_75t_L g4793 ( 
.A(n_4235),
.B(n_628),
.Y(n_4793)
);

BUFx3_ASAP7_75t_L g4794 ( 
.A(n_4180),
.Y(n_4794)
);

OAI21xp5_ASAP7_75t_L g4795 ( 
.A1(n_4352),
.A2(n_629),
.B(n_631),
.Y(n_4795)
);

OA21x2_ASAP7_75t_L g4796 ( 
.A1(n_4390),
.A2(n_629),
.B(n_632),
.Y(n_4796)
);

INVx1_ASAP7_75t_SL g4797 ( 
.A(n_4173),
.Y(n_4797)
);

AOI21xp5_ASAP7_75t_L g4798 ( 
.A1(n_4465),
.A2(n_632),
.B(n_633),
.Y(n_4798)
);

AOI21x1_ASAP7_75t_L g4799 ( 
.A1(n_4497),
.A2(n_632),
.B(n_634),
.Y(n_4799)
);

OAI21x1_ASAP7_75t_L g4800 ( 
.A1(n_4372),
.A2(n_783),
.B(n_782),
.Y(n_4800)
);

OAI21x1_ASAP7_75t_L g4801 ( 
.A1(n_4401),
.A2(n_784),
.B(n_782),
.Y(n_4801)
);

NOR4xp25_ASAP7_75t_L g4802 ( 
.A(n_4492),
.B(n_4526),
.C(n_4387),
.D(n_4229),
.Y(n_4802)
);

AO21x2_ASAP7_75t_L g4803 ( 
.A1(n_4179),
.A2(n_634),
.B(n_635),
.Y(n_4803)
);

NOR2x1_ASAP7_75t_SL g4804 ( 
.A(n_4255),
.B(n_635),
.Y(n_4804)
);

OR2x6_ASAP7_75t_L g4805 ( 
.A(n_4346),
.B(n_635),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4525),
.Y(n_4806)
);

HB1xp67_ASAP7_75t_L g4807 ( 
.A(n_4396),
.Y(n_4807)
);

NOR2x1_ASAP7_75t_L g4808 ( 
.A(n_4220),
.B(n_636),
.Y(n_4808)
);

OAI21x1_ASAP7_75t_L g4809 ( 
.A1(n_4414),
.A2(n_4554),
.B(n_4495),
.Y(n_4809)
);

AO31x2_ASAP7_75t_L g4810 ( 
.A1(n_4339),
.A2(n_4359),
.A3(n_4407),
.B(n_4361),
.Y(n_4810)
);

OAI21x1_ASAP7_75t_L g4811 ( 
.A1(n_4418),
.A2(n_787),
.B(n_786),
.Y(n_4811)
);

OA21x2_ASAP7_75t_L g4812 ( 
.A1(n_4421),
.A2(n_636),
.B(n_637),
.Y(n_4812)
);

OAI22xp5_ASAP7_75t_SL g4813 ( 
.A1(n_4241),
.A2(n_638),
.B1(n_636),
.B2(n_637),
.Y(n_4813)
);

OAI21x1_ASAP7_75t_L g4814 ( 
.A1(n_4423),
.A2(n_790),
.B(n_789),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4355),
.Y(n_4815)
);

OA21x2_ASAP7_75t_L g4816 ( 
.A1(n_4471),
.A2(n_637),
.B(n_638),
.Y(n_4816)
);

O2A1O1Ixp33_ASAP7_75t_L g4817 ( 
.A1(n_4504),
.A2(n_640),
.B(n_638),
.C(n_639),
.Y(n_4817)
);

OAI21xp5_ASAP7_75t_L g4818 ( 
.A1(n_4381),
.A2(n_639),
.B(n_640),
.Y(n_4818)
);

AND2x4_ASAP7_75t_L g4819 ( 
.A(n_4176),
.B(n_4409),
.Y(n_4819)
);

INVx2_ASAP7_75t_L g4820 ( 
.A(n_4564),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4810),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4810),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4806),
.Y(n_4823)
);

INVx2_ASAP7_75t_L g4824 ( 
.A(n_4575),
.Y(n_4824)
);

INVx3_ASAP7_75t_L g4825 ( 
.A(n_4610),
.Y(n_4825)
);

INVx2_ASAP7_75t_L g4826 ( 
.A(n_4591),
.Y(n_4826)
);

BUFx2_ASAP7_75t_R g4827 ( 
.A(n_4673),
.Y(n_4827)
);

INVx3_ASAP7_75t_L g4828 ( 
.A(n_4577),
.Y(n_4828)
);

BUFx2_ASAP7_75t_L g4829 ( 
.A(n_4559),
.Y(n_4829)
);

AO21x2_ASAP7_75t_L g4830 ( 
.A1(n_4558),
.A2(n_4314),
.B(n_4302),
.Y(n_4830)
);

AO21x2_ASAP7_75t_L g4831 ( 
.A1(n_4621),
.A2(n_4376),
.B(n_4332),
.Y(n_4831)
);

BUFx3_ASAP7_75t_L g4832 ( 
.A(n_4583),
.Y(n_4832)
);

OAI21x1_ASAP7_75t_SL g4833 ( 
.A1(n_4804),
.A2(n_4741),
.B(n_4784),
.Y(n_4833)
);

NOR2xp67_ASAP7_75t_SL g4834 ( 
.A(n_4783),
.B(n_4197),
.Y(n_4834)
);

AOI22xp33_ASAP7_75t_SL g4835 ( 
.A1(n_4807),
.A2(n_4391),
.B1(n_4713),
.B2(n_4425),
.Y(n_4835)
);

AND2x2_ASAP7_75t_L g4836 ( 
.A(n_4637),
.B(n_4395),
.Y(n_4836)
);

OAI22xp33_ASAP7_75t_L g4837 ( 
.A1(n_4763),
.A2(n_4440),
.B1(n_4400),
.B2(n_4428),
.Y(n_4837)
);

AO21x2_ASAP7_75t_L g4838 ( 
.A1(n_4704),
.A2(n_4397),
.B(n_4385),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4570),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4584),
.Y(n_4840)
);

AOI22xp33_ASAP7_75t_L g4841 ( 
.A1(n_4631),
.A2(n_4436),
.B1(n_4508),
.B2(n_4548),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4588),
.Y(n_4842)
);

INVx2_ASAP7_75t_L g4843 ( 
.A(n_4600),
.Y(n_4843)
);

OAI21x1_ASAP7_75t_L g4844 ( 
.A1(n_4574),
.A2(n_4156),
.B(n_4192),
.Y(n_4844)
);

AOI22xp33_ASAP7_75t_L g4845 ( 
.A1(n_4631),
.A2(n_4429),
.B1(n_4487),
.B2(n_4482),
.Y(n_4845)
);

AND2x2_ASAP7_75t_L g4846 ( 
.A(n_4637),
.B(n_4358),
.Y(n_4846)
);

AOI22xp5_ASAP7_75t_L g4847 ( 
.A1(n_4560),
.A2(n_4486),
.B1(n_4360),
.B2(n_4533),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4599),
.Y(n_4848)
);

AND2x4_ASAP7_75t_L g4849 ( 
.A(n_4768),
.B(n_4428),
.Y(n_4849)
);

HB1xp67_ASAP7_75t_L g4850 ( 
.A(n_4691),
.Y(n_4850)
);

HB1xp67_ASAP7_75t_L g4851 ( 
.A(n_4622),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4608),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4609),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4615),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4627),
.Y(n_4855)
);

CKINVDCx11_ASAP7_75t_R g4856 ( 
.A(n_4592),
.Y(n_4856)
);

AOI21x1_ASAP7_75t_L g4857 ( 
.A1(n_4657),
.A2(n_4281),
.B(n_4398),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4641),
.Y(n_4858)
);

OA21x2_ASAP7_75t_L g4859 ( 
.A1(n_4567),
.A2(n_4491),
.B(n_4490),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4649),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4662),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4665),
.Y(n_4862)
);

AOI22xp5_ASAP7_75t_L g4863 ( 
.A1(n_4631),
.A2(n_4469),
.B1(n_4519),
.B2(n_4522),
.Y(n_4863)
);

OAI21x1_ASAP7_75t_L g4864 ( 
.A1(n_4572),
.A2(n_4398),
.B(n_4273),
.Y(n_4864)
);

AOI22xp33_ASAP7_75t_L g4865 ( 
.A1(n_4601),
.A2(n_4507),
.B1(n_4542),
.B2(n_4476),
.Y(n_4865)
);

AOI21x1_ASAP7_75t_L g4866 ( 
.A1(n_4799),
.A2(n_4502),
.B(n_4218),
.Y(n_4866)
);

HB1xp67_ASAP7_75t_L g4867 ( 
.A(n_4712),
.Y(n_4867)
);

OA21x2_ASAP7_75t_L g4868 ( 
.A1(n_4565),
.A2(n_4509),
.B(n_4506),
.Y(n_4868)
);

OR2x6_ASAP7_75t_L g4869 ( 
.A(n_4763),
.B(n_4386),
.Y(n_4869)
);

INVx2_ASAP7_75t_L g4870 ( 
.A(n_4625),
.Y(n_4870)
);

BUFx2_ASAP7_75t_L g4871 ( 
.A(n_4581),
.Y(n_4871)
);

HB1xp67_ASAP7_75t_L g4872 ( 
.A(n_4781),
.Y(n_4872)
);

OAI21x1_ASAP7_75t_SL g4873 ( 
.A1(n_4750),
.A2(n_4201),
.B(n_4167),
.Y(n_4873)
);

INVx2_ASAP7_75t_L g4874 ( 
.A(n_4638),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4682),
.Y(n_4875)
);

CKINVDCx20_ASAP7_75t_R g4876 ( 
.A(n_4664),
.Y(n_4876)
);

INVx2_ASAP7_75t_L g4877 ( 
.A(n_4660),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4692),
.Y(n_4878)
);

AND2x2_ASAP7_75t_L g4879 ( 
.A(n_4739),
.B(n_4262),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4711),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4714),
.Y(n_4881)
);

INVx2_ASAP7_75t_L g4882 ( 
.A(n_4661),
.Y(n_4882)
);

INVx2_ASAP7_75t_SL g4883 ( 
.A(n_4696),
.Y(n_4883)
);

OR2x6_ASAP7_75t_L g4884 ( 
.A(n_4624),
.B(n_4386),
.Y(n_4884)
);

INVx6_ASAP7_75t_L g4885 ( 
.A(n_4698),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4667),
.Y(n_4886)
);

AO21x1_ASAP7_75t_SL g4887 ( 
.A1(n_4701),
.A2(n_4478),
.B(n_4197),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4733),
.Y(n_4888)
);

HB1xp67_ASAP7_75t_L g4889 ( 
.A(n_4734),
.Y(n_4889)
);

OAI22xp5_ASAP7_75t_L g4890 ( 
.A1(n_4598),
.A2(n_4318),
.B1(n_4438),
.B2(n_4543),
.Y(n_4890)
);

INVx2_ASAP7_75t_L g4891 ( 
.A(n_4672),
.Y(n_4891)
);

CKINVDCx5p33_ASAP7_75t_R g4892 ( 
.A(n_4562),
.Y(n_4892)
);

AOI22xp33_ASAP7_75t_L g4893 ( 
.A1(n_4623),
.A2(n_4456),
.B1(n_4481),
.B2(n_4452),
.Y(n_4893)
);

AOI22xp33_ASAP7_75t_SL g4894 ( 
.A1(n_4719),
.A2(n_4431),
.B1(n_4438),
.B2(n_4350),
.Y(n_4894)
);

HB1xp67_ASAP7_75t_L g4895 ( 
.A(n_4737),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4680),
.Y(n_4896)
);

AOI22xp33_ASAP7_75t_L g4897 ( 
.A1(n_4598),
.A2(n_4399),
.B1(n_4555),
.B2(n_4389),
.Y(n_4897)
);

INVx2_ASAP7_75t_SL g4898 ( 
.A(n_4696),
.Y(n_4898)
);

BUFx6f_ASAP7_75t_L g4899 ( 
.A(n_4753),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4686),
.Y(n_4900)
);

OAI22xp5_ASAP7_75t_L g4901 ( 
.A1(n_4670),
.A2(n_4445),
.B1(n_4441),
.B2(n_4453),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4709),
.Y(n_4902)
);

CKINVDCx5p33_ASAP7_75t_R g4903 ( 
.A(n_4578),
.Y(n_4903)
);

AOI22xp33_ASAP7_75t_SL g4904 ( 
.A1(n_4719),
.A2(n_4488),
.B1(n_4473),
.B2(n_4458),
.Y(n_4904)
);

INVx2_ASAP7_75t_L g4905 ( 
.A(n_4715),
.Y(n_4905)
);

AOI22xp5_ASAP7_75t_L g4906 ( 
.A1(n_4813),
.A2(n_4534),
.B1(n_4531),
.B2(n_4544),
.Y(n_4906)
);

AND2x2_ASAP7_75t_L g4907 ( 
.A(n_4731),
.B(n_4444),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4744),
.Y(n_4908)
);

INVx2_ASAP7_75t_L g4909 ( 
.A(n_4593),
.Y(n_4909)
);

AND2x2_ASAP7_75t_L g4910 ( 
.A(n_4593),
.B(n_4349),
.Y(n_4910)
);

OAI22xp33_ASAP7_75t_L g4911 ( 
.A1(n_4670),
.A2(n_4310),
.B1(n_4265),
.B2(n_4250),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4755),
.Y(n_4912)
);

OAI21x1_ASAP7_75t_L g4913 ( 
.A1(n_4566),
.A2(n_4498),
.B(n_4475),
.Y(n_4913)
);

OAI21x1_ASAP7_75t_L g4914 ( 
.A1(n_4809),
.A2(n_4521),
.B(n_4513),
.Y(n_4914)
);

AND2x2_ASAP7_75t_L g4915 ( 
.A(n_4789),
.B(n_4349),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4630),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4630),
.Y(n_4917)
);

AND2x2_ASAP7_75t_L g4918 ( 
.A(n_4725),
.B(n_4218),
.Y(n_4918)
);

BUFx2_ASAP7_75t_L g4919 ( 
.A(n_4775),
.Y(n_4919)
);

INVx2_ASAP7_75t_L g4920 ( 
.A(n_4779),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_4729),
.Y(n_4921)
);

AND2x2_ASAP7_75t_L g4922 ( 
.A(n_4726),
.B(n_4503),
.Y(n_4922)
);

OAI21x1_ASAP7_75t_L g4923 ( 
.A1(n_4605),
.A2(n_4540),
.B(n_4530),
.Y(n_4923)
);

OAI21x1_ASAP7_75t_L g4924 ( 
.A1(n_4612),
.A2(n_4616),
.B(n_4596),
.Y(n_4924)
);

INVx2_ASAP7_75t_L g4925 ( 
.A(n_4746),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4752),
.Y(n_4926)
);

INVx2_ASAP7_75t_L g4927 ( 
.A(n_4757),
.Y(n_4927)
);

AOI22xp33_ASAP7_75t_SL g4928 ( 
.A1(n_4606),
.A2(n_4780),
.B1(n_4786),
.B2(n_4689),
.Y(n_4928)
);

BUFx6f_ASAP7_75t_L g4929 ( 
.A(n_4753),
.Y(n_4929)
);

INVx2_ASAP7_75t_L g4930 ( 
.A(n_4764),
.Y(n_4930)
);

BUFx2_ASAP7_75t_L g4931 ( 
.A(n_4586),
.Y(n_4931)
);

HB1xp67_ASAP7_75t_L g4932 ( 
.A(n_4620),
.Y(n_4932)
);

NOR2xp33_ASAP7_75t_L g4933 ( 
.A(n_4735),
.B(n_4541),
.Y(n_4933)
);

AND2x2_ASAP7_75t_L g4934 ( 
.A(n_4815),
.B(n_4505),
.Y(n_4934)
);

INVx2_ASAP7_75t_L g4935 ( 
.A(n_4589),
.Y(n_4935)
);

BUFx2_ASAP7_75t_L g4936 ( 
.A(n_4819),
.Y(n_4936)
);

INVx2_ASAP7_75t_SL g4937 ( 
.A(n_4732),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4561),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4561),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4655),
.Y(n_4940)
);

CKINVDCx5p33_ASAP7_75t_R g4941 ( 
.A(n_4618),
.Y(n_4941)
);

INVx2_ASAP7_75t_L g4942 ( 
.A(n_4589),
.Y(n_4942)
);

OAI21x1_ASAP7_75t_L g4943 ( 
.A1(n_4640),
.A2(n_4477),
.B(n_4448),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4655),
.Y(n_4944)
);

HB1xp67_ASAP7_75t_L g4945 ( 
.A(n_4802),
.Y(n_4945)
);

AND2x4_ASAP7_75t_L g4946 ( 
.A(n_4708),
.B(n_4794),
.Y(n_4946)
);

BUFx12f_ASAP7_75t_L g4947 ( 
.A(n_4676),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_4571),
.Y(n_4948)
);

AOI21xp33_ASAP7_75t_SL g4949 ( 
.A1(n_4690),
.A2(n_4222),
.B(n_4294),
.Y(n_4949)
);

INVx2_ASAP7_75t_L g4950 ( 
.A(n_4571),
.Y(n_4950)
);

OA21x2_ASAP7_75t_L g4951 ( 
.A1(n_4614),
.A2(n_4545),
.B(n_4333),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4730),
.Y(n_4952)
);

INVx6_ASAP7_75t_L g4953 ( 
.A(n_4724),
.Y(n_4953)
);

INVx2_ASAP7_75t_L g4954 ( 
.A(n_4628),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4639),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4700),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4645),
.B(n_4517),
.Y(n_4957)
);

AND2x2_ASAP7_75t_L g4958 ( 
.A(n_4645),
.B(n_4766),
.Y(n_4958)
);

INVx2_ASAP7_75t_L g4959 ( 
.A(n_4710),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4782),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4889),
.Y(n_4961)
);

NOR2xp33_ASAP7_75t_R g4962 ( 
.A(n_4876),
.B(n_4585),
.Y(n_4962)
);

OR2x2_ASAP7_75t_SL g4963 ( 
.A(n_4885),
.B(n_4732),
.Y(n_4963)
);

INVx2_ASAP7_75t_L g4964 ( 
.A(n_4829),
.Y(n_4964)
);

OR2x2_ASAP7_75t_L g4965 ( 
.A(n_4850),
.B(n_4829),
.Y(n_4965)
);

AND2x2_ASAP7_75t_L g4966 ( 
.A(n_4867),
.B(n_4797),
.Y(n_4966)
);

CKINVDCx20_ASAP7_75t_R g4967 ( 
.A(n_4856),
.Y(n_4967)
);

INVxp33_ASAP7_75t_SL g4968 ( 
.A(n_4834),
.Y(n_4968)
);

INVx1_ASAP7_75t_SL g4969 ( 
.A(n_4832),
.Y(n_4969)
);

INVx2_ASAP7_75t_L g4970 ( 
.A(n_4919),
.Y(n_4970)
);

AND2x2_ASAP7_75t_L g4971 ( 
.A(n_4871),
.B(n_4705),
.Y(n_4971)
);

NAND2xp5_ASAP7_75t_L g4972 ( 
.A(n_4938),
.B(n_4687),
.Y(n_4972)
);

AO32x2_ASAP7_75t_L g4973 ( 
.A1(n_4890),
.A2(n_4684),
.A3(n_4594),
.B1(n_4675),
.B2(n_4723),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4895),
.Y(n_4974)
);

AOI22xp33_ASAP7_75t_L g4975 ( 
.A1(n_4830),
.A2(n_4579),
.B1(n_4772),
.B2(n_4597),
.Y(n_4975)
);

INVx2_ASAP7_75t_L g4976 ( 
.A(n_4859),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4939),
.B(n_4740),
.Y(n_4977)
);

OAI22xp5_ASAP7_75t_L g4978 ( 
.A1(n_4928),
.A2(n_4787),
.B1(n_4805),
.B2(n_4603),
.Y(n_4978)
);

OAI22xp33_ASAP7_75t_L g4979 ( 
.A1(n_4869),
.A2(n_4805),
.B1(n_4677),
.B2(n_4716),
.Y(n_4979)
);

OR2x6_ASAP7_75t_L g4980 ( 
.A(n_4869),
.B(n_4658),
.Y(n_4980)
);

CKINVDCx5p33_ASAP7_75t_R g4981 ( 
.A(n_4892),
.Y(n_4981)
);

INVx2_ASAP7_75t_L g4982 ( 
.A(n_4859),
.Y(n_4982)
);

HB1xp67_ASAP7_75t_L g4983 ( 
.A(n_4851),
.Y(n_4983)
);

AND2x2_ASAP7_75t_L g4984 ( 
.A(n_4871),
.B(n_4306),
.Y(n_4984)
);

INVx2_ASAP7_75t_L g4985 ( 
.A(n_4935),
.Y(n_4985)
);

NAND2xp5_ASAP7_75t_L g4986 ( 
.A(n_4916),
.B(n_4576),
.Y(n_4986)
);

OA21x2_ASAP7_75t_L g4987 ( 
.A1(n_4873),
.A2(n_4702),
.B(n_4569),
.Y(n_4987)
);

OR2x6_ASAP7_75t_L g4988 ( 
.A(n_4884),
.B(n_4666),
.Y(n_4988)
);

AND2x2_ASAP7_75t_L g4989 ( 
.A(n_4942),
.B(n_4754),
.Y(n_4989)
);

NOR2xp33_ASAP7_75t_R g4990 ( 
.A(n_4903),
.B(n_4263),
.Y(n_4990)
);

CKINVDCx5p33_ASAP7_75t_R g4991 ( 
.A(n_4947),
.Y(n_4991)
);

CKINVDCx5p33_ASAP7_75t_R g4992 ( 
.A(n_4941),
.Y(n_4992)
);

CKINVDCx5p33_ASAP7_75t_R g4993 ( 
.A(n_4827),
.Y(n_4993)
);

AND2x2_ASAP7_75t_L g4994 ( 
.A(n_4846),
.B(n_4340),
.Y(n_4994)
);

OAI21xp5_ASAP7_75t_L g4995 ( 
.A1(n_4866),
.A2(n_4808),
.B(n_4857),
.Y(n_4995)
);

AOI22xp33_ASAP7_75t_L g4996 ( 
.A1(n_4865),
.A2(n_4534),
.B1(n_4531),
.B2(n_4479),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4917),
.B(n_4602),
.Y(n_4997)
);

INVx2_ASAP7_75t_SL g4998 ( 
.A(n_4885),
.Y(n_4998)
);

CKINVDCx16_ASAP7_75t_R g4999 ( 
.A(n_4946),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4839),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4840),
.Y(n_5001)
);

AOI222xp33_ASAP7_75t_L g5002 ( 
.A1(n_4901),
.A2(n_4613),
.B1(n_4756),
.B2(n_4669),
.C1(n_4635),
.C2(n_4582),
.Y(n_5002)
);

NOR2x1_ASAP7_75t_L g5003 ( 
.A(n_4884),
.B(n_4629),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4836),
.B(n_4304),
.Y(n_5004)
);

INVx1_ASAP7_75t_L g5005 ( 
.A(n_4842),
.Y(n_5005)
);

AND2x2_ASAP7_75t_L g5006 ( 
.A(n_4909),
.B(n_4747),
.Y(n_5006)
);

INVxp67_ASAP7_75t_L g5007 ( 
.A(n_4931),
.Y(n_5007)
);

NOR2x1_ASAP7_75t_L g5008 ( 
.A(n_4911),
.B(n_4642),
.Y(n_5008)
);

A2O1A1Ixp33_ASAP7_75t_L g5009 ( 
.A1(n_4904),
.A2(n_4762),
.B(n_4679),
.C(n_4587),
.Y(n_5009)
);

AO21x1_ASAP7_75t_L g5010 ( 
.A1(n_4945),
.A2(n_4681),
.B(n_4683),
.Y(n_5010)
);

OR2x6_ASAP7_75t_L g5011 ( 
.A(n_4953),
.B(n_4703),
.Y(n_5011)
);

BUFx2_ASAP7_75t_L g5012 ( 
.A(n_4936),
.Y(n_5012)
);

OAI21xp5_ASAP7_75t_L g5013 ( 
.A1(n_4847),
.A2(n_4863),
.B(n_4773),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4848),
.Y(n_5014)
);

NOR2xp33_ASAP7_75t_R g5015 ( 
.A(n_4825),
.B(n_4209),
.Y(n_5015)
);

OR2x6_ASAP7_75t_L g5016 ( 
.A(n_4953),
.B(n_4674),
.Y(n_5016)
);

INVxp67_ASAP7_75t_L g5017 ( 
.A(n_4872),
.Y(n_5017)
);

NOR2xp33_ASAP7_75t_R g5018 ( 
.A(n_4937),
.B(n_4269),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4852),
.Y(n_5019)
);

OR2x2_ASAP7_75t_L g5020 ( 
.A(n_4948),
.B(n_4417),
.Y(n_5020)
);

INVx2_ASAP7_75t_L g5021 ( 
.A(n_4950),
.Y(n_5021)
);

INVx1_ASAP7_75t_SL g5022 ( 
.A(n_4879),
.Y(n_5022)
);

BUFx3_ASAP7_75t_L g5023 ( 
.A(n_4828),
.Y(n_5023)
);

O2A1O1Ixp33_ASAP7_75t_SL g5024 ( 
.A1(n_4837),
.A2(n_4694),
.B(n_4721),
.C(n_4728),
.Y(n_5024)
);

XOR2x2_ASAP7_75t_SL g5025 ( 
.A(n_4894),
.B(n_4693),
.Y(n_5025)
);

AND2x4_ASAP7_75t_SL g5026 ( 
.A(n_4849),
.B(n_4152),
.Y(n_5026)
);

BUFx3_ASAP7_75t_L g5027 ( 
.A(n_4922),
.Y(n_5027)
);

BUFx6f_ASAP7_75t_L g5028 ( 
.A(n_4899),
.Y(n_5028)
);

NAND2xp33_ASAP7_75t_R g5029 ( 
.A(n_4936),
.B(n_4793),
.Y(n_5029)
);

BUFx3_ASAP7_75t_L g5030 ( 
.A(n_4899),
.Y(n_5030)
);

INVx2_ASAP7_75t_L g5031 ( 
.A(n_4820),
.Y(n_5031)
);

AND2x4_ASAP7_75t_L g5032 ( 
.A(n_4910),
.B(n_4958),
.Y(n_5032)
);

NAND2xp5_ASAP7_75t_L g5033 ( 
.A(n_4921),
.B(n_4769),
.Y(n_5033)
);

AND2x4_ASAP7_75t_L g5034 ( 
.A(n_4915),
.B(n_4940),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4853),
.Y(n_5035)
);

INVx2_ASAP7_75t_SL g5036 ( 
.A(n_4929),
.Y(n_5036)
);

INVx2_ASAP7_75t_L g5037 ( 
.A(n_4824),
.Y(n_5037)
);

HB1xp67_ASAP7_75t_L g5038 ( 
.A(n_4918),
.Y(n_5038)
);

OAI21xp5_ASAP7_75t_L g5039 ( 
.A1(n_4835),
.A2(n_4771),
.B(n_4817),
.Y(n_5039)
);

AND2x2_ASAP7_75t_L g5040 ( 
.A(n_4907),
.B(n_4224),
.Y(n_5040)
);

NAND2xp33_ASAP7_75t_R g5041 ( 
.A(n_4949),
.B(n_4796),
.Y(n_5041)
);

INVx2_ASAP7_75t_L g5042 ( 
.A(n_4826),
.Y(n_5042)
);

CKINVDCx16_ASAP7_75t_R g5043 ( 
.A(n_4933),
.Y(n_5043)
);

AO31x2_ASAP7_75t_L g5044 ( 
.A1(n_4821),
.A2(n_4563),
.A3(n_4759),
.B(n_4607),
.Y(n_5044)
);

AO31x2_ASAP7_75t_L g5045 ( 
.A1(n_4822),
.A2(n_4651),
.A3(n_4697),
.B(n_4742),
.Y(n_5045)
);

OR2x6_ASAP7_75t_L g5046 ( 
.A(n_4833),
.B(n_4648),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_4854),
.Y(n_5047)
);

AOI22xp33_ASAP7_75t_L g5048 ( 
.A1(n_4831),
.A2(n_4494),
.B1(n_4516),
.B2(n_4538),
.Y(n_5048)
);

AND2x2_ASAP7_75t_L g5049 ( 
.A(n_4932),
.B(n_4934),
.Y(n_5049)
);

OR2x6_ASAP7_75t_L g5050 ( 
.A(n_4864),
.B(n_4722),
.Y(n_5050)
);

NOR2xp33_ASAP7_75t_L g5051 ( 
.A(n_4952),
.B(n_4153),
.Y(n_5051)
);

INVxp67_ASAP7_75t_L g5052 ( 
.A(n_4957),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4855),
.Y(n_5053)
);

OAI21xp5_ASAP7_75t_SL g5054 ( 
.A1(n_4906),
.A2(n_4654),
.B(n_4760),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_4858),
.Y(n_5055)
);

AND2x2_ASAP7_75t_L g5056 ( 
.A(n_4944),
.B(n_4412),
.Y(n_5056)
);

AOI22xp33_ASAP7_75t_L g5057 ( 
.A1(n_4893),
.A2(n_4646),
.B1(n_4580),
.B2(n_4653),
.Y(n_5057)
);

NAND2xp5_ASAP7_75t_L g5058 ( 
.A(n_4926),
.B(n_4611),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_4860),
.Y(n_5059)
);

AND2x2_ASAP7_75t_L g5060 ( 
.A(n_4920),
.B(n_4412),
.Y(n_5060)
);

AND2x4_ASAP7_75t_L g5061 ( 
.A(n_4883),
.B(n_4186),
.Y(n_5061)
);

NOR2xp67_ASAP7_75t_L g5062 ( 
.A(n_4954),
.B(n_4765),
.Y(n_5062)
);

AND2x4_ASAP7_75t_L g5063 ( 
.A(n_4898),
.B(n_4280),
.Y(n_5063)
);

AND2x2_ASAP7_75t_L g5064 ( 
.A(n_4823),
.B(n_4535),
.Y(n_5064)
);

NAND5xp2_ASAP7_75t_L g5065 ( 
.A(n_5002),
.B(n_4897),
.C(n_4841),
.D(n_4604),
.E(n_4845),
.Y(n_5065)
);

AND2x2_ASAP7_75t_L g5066 ( 
.A(n_5012),
.B(n_4955),
.Y(n_5066)
);

HB1xp67_ASAP7_75t_L g5067 ( 
.A(n_4983),
.Y(n_5067)
);

AO22x1_ASAP7_75t_L g5068 ( 
.A1(n_5003),
.A2(n_4380),
.B1(n_4959),
.B2(n_4296),
.Y(n_5068)
);

INVx2_ASAP7_75t_L g5069 ( 
.A(n_4965),
.Y(n_5069)
);

AND2x2_ASAP7_75t_L g5070 ( 
.A(n_5049),
.B(n_4956),
.Y(n_5070)
);

AND2x2_ASAP7_75t_L g5071 ( 
.A(n_4966),
.B(n_4951),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4976),
.Y(n_5072)
);

AND2x2_ASAP7_75t_L g5073 ( 
.A(n_5032),
.B(n_4951),
.Y(n_5073)
);

INVx2_ASAP7_75t_L g5074 ( 
.A(n_4982),
.Y(n_5074)
);

INVxp67_ASAP7_75t_L g5075 ( 
.A(n_5029),
.Y(n_5075)
);

INVx3_ASAP7_75t_L g5076 ( 
.A(n_4999),
.Y(n_5076)
);

AND2x2_ASAP7_75t_L g5077 ( 
.A(n_5038),
.B(n_4908),
.Y(n_5077)
);

INVx2_ASAP7_75t_L g5078 ( 
.A(n_4970),
.Y(n_5078)
);

NAND2xp5_ASAP7_75t_L g5079 ( 
.A(n_4986),
.B(n_4960),
.Y(n_5079)
);

BUFx3_ASAP7_75t_L g5080 ( 
.A(n_4969),
.Y(n_5080)
);

AND2x4_ASAP7_75t_L g5081 ( 
.A(n_5062),
.B(n_4923),
.Y(n_5081)
);

OR2x2_ASAP7_75t_L g5082 ( 
.A(n_4972),
.B(n_4925),
.Y(n_5082)
);

INVx2_ASAP7_75t_L g5083 ( 
.A(n_4964),
.Y(n_5083)
);

OAI22xp5_ASAP7_75t_L g5084 ( 
.A1(n_4963),
.A2(n_4980),
.B1(n_4988),
.B2(n_4975),
.Y(n_5084)
);

INVxp67_ASAP7_75t_SL g5085 ( 
.A(n_5025),
.Y(n_5085)
);

BUFx6f_ASAP7_75t_SL g5086 ( 
.A(n_5016),
.Y(n_5086)
);

AND2x2_ASAP7_75t_L g5087 ( 
.A(n_5022),
.B(n_4912),
.Y(n_5087)
);

AND2x4_ASAP7_75t_L g5088 ( 
.A(n_5050),
.B(n_4844),
.Y(n_5088)
);

BUFx2_ASAP7_75t_L g5089 ( 
.A(n_5015),
.Y(n_5089)
);

AND2x2_ASAP7_75t_L g5090 ( 
.A(n_4984),
.B(n_4880),
.Y(n_5090)
);

NAND2xp5_ASAP7_75t_L g5091 ( 
.A(n_4977),
.B(n_4881),
.Y(n_5091)
);

AND2x2_ASAP7_75t_L g5092 ( 
.A(n_5027),
.B(n_4888),
.Y(n_5092)
);

OR2x2_ASAP7_75t_L g5093 ( 
.A(n_4985),
.B(n_4891),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_5031),
.Y(n_5094)
);

INVx2_ASAP7_75t_L g5095 ( 
.A(n_5037),
.Y(n_5095)
);

AND2x4_ASAP7_75t_L g5096 ( 
.A(n_5050),
.B(n_4914),
.Y(n_5096)
);

AND2x2_ASAP7_75t_L g5097 ( 
.A(n_4971),
.B(n_5034),
.Y(n_5097)
);

INVx3_ASAP7_75t_L g5098 ( 
.A(n_4987),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_4961),
.Y(n_5099)
);

INVx2_ASAP7_75t_L g5100 ( 
.A(n_5042),
.Y(n_5100)
);

INVx2_ASAP7_75t_L g5101 ( 
.A(n_5021),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_4974),
.Y(n_5102)
);

CKINVDCx20_ASAP7_75t_R g5103 ( 
.A(n_4967),
.Y(n_5103)
);

NOR2x1_ASAP7_75t_SL g5104 ( 
.A(n_4988),
.B(n_4887),
.Y(n_5104)
);

AND2x2_ASAP7_75t_L g5105 ( 
.A(n_4989),
.B(n_4927),
.Y(n_5105)
);

AND2x2_ASAP7_75t_L g5106 ( 
.A(n_5007),
.B(n_4930),
.Y(n_5106)
);

BUFx3_ASAP7_75t_L g5107 ( 
.A(n_4991),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_5000),
.Y(n_5108)
);

OR2x2_ASAP7_75t_L g5109 ( 
.A(n_5017),
.B(n_4997),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_5001),
.Y(n_5110)
);

BUFx3_ASAP7_75t_L g5111 ( 
.A(n_4998),
.Y(n_5111)
);

INVx2_ASAP7_75t_L g5112 ( 
.A(n_5005),
.Y(n_5112)
);

AND2x2_ASAP7_75t_L g5113 ( 
.A(n_5006),
.B(n_4905),
.Y(n_5113)
);

INVx2_ASAP7_75t_L g5114 ( 
.A(n_5014),
.Y(n_5114)
);

BUFx3_ASAP7_75t_L g5115 ( 
.A(n_4992),
.Y(n_5115)
);

AND2x2_ASAP7_75t_L g5116 ( 
.A(n_5052),
.B(n_4875),
.Y(n_5116)
);

AND2x4_ASAP7_75t_L g5117 ( 
.A(n_4980),
.B(n_4913),
.Y(n_5117)
);

AND2x4_ASAP7_75t_L g5118 ( 
.A(n_5056),
.B(n_4886),
.Y(n_5118)
);

BUFx3_ASAP7_75t_L g5119 ( 
.A(n_5040),
.Y(n_5119)
);

NAND2xp5_ASAP7_75t_L g5120 ( 
.A(n_5019),
.B(n_4896),
.Y(n_5120)
);

AND2x2_ASAP7_75t_L g5121 ( 
.A(n_5064),
.B(n_4878),
.Y(n_5121)
);

OR2x2_ASAP7_75t_L g5122 ( 
.A(n_5058),
.B(n_4900),
.Y(n_5122)
);

INVx2_ASAP7_75t_L g5123 ( 
.A(n_5035),
.Y(n_5123)
);

BUFx3_ASAP7_75t_L g5124 ( 
.A(n_4981),
.Y(n_5124)
);

INVx3_ASAP7_75t_L g5125 ( 
.A(n_5011),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_5047),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_5053),
.Y(n_5127)
);

INVx3_ASAP7_75t_L g5128 ( 
.A(n_5011),
.Y(n_5128)
);

BUFx3_ASAP7_75t_L g5129 ( 
.A(n_5004),
.Y(n_5129)
);

INVxp67_ASAP7_75t_SL g5130 ( 
.A(n_5008),
.Y(n_5130)
);

AOI221x1_ASAP7_75t_SL g5131 ( 
.A1(n_4979),
.A2(n_4718),
.B1(n_4791),
.B2(n_4227),
.C(n_4454),
.Y(n_5131)
);

INVx2_ASAP7_75t_L g5132 ( 
.A(n_5055),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_5059),
.Y(n_5133)
);

INVx2_ASAP7_75t_L g5134 ( 
.A(n_5020),
.Y(n_5134)
);

AND2x4_ASAP7_75t_L g5135 ( 
.A(n_5048),
.B(n_5036),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_5033),
.Y(n_5136)
);

INVx2_ASAP7_75t_L g5137 ( 
.A(n_5060),
.Y(n_5137)
);

HB1xp67_ASAP7_75t_L g5138 ( 
.A(n_5023),
.Y(n_5138)
);

INVx2_ASAP7_75t_L g5139 ( 
.A(n_5063),
.Y(n_5139)
);

NOR2xp33_ASAP7_75t_L g5140 ( 
.A(n_4993),
.B(n_4153),
.Y(n_5140)
);

HB1xp67_ASAP7_75t_L g5141 ( 
.A(n_4994),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_5051),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_5044),
.Y(n_5143)
);

BUFx2_ASAP7_75t_L g5144 ( 
.A(n_5018),
.Y(n_5144)
);

AND2x2_ASAP7_75t_L g5145 ( 
.A(n_5030),
.B(n_4861),
.Y(n_5145)
);

INVx2_ASAP7_75t_L g5146 ( 
.A(n_5061),
.Y(n_5146)
);

NAND2xp5_ASAP7_75t_L g5147 ( 
.A(n_5045),
.B(n_4902),
.Y(n_5147)
);

INVx2_ASAP7_75t_SL g5148 ( 
.A(n_4962),
.Y(n_5148)
);

AOI22xp5_ASAP7_75t_L g5149 ( 
.A1(n_5085),
.A2(n_5041),
.B1(n_4968),
.B2(n_5013),
.Y(n_5149)
);

BUFx3_ASAP7_75t_L g5150 ( 
.A(n_5080),
.Y(n_5150)
);

NAND2xp5_ASAP7_75t_L g5151 ( 
.A(n_5079),
.B(n_5045),
.Y(n_5151)
);

INVx3_ASAP7_75t_L g5152 ( 
.A(n_5076),
.Y(n_5152)
);

OAI21x1_ASAP7_75t_L g5153 ( 
.A1(n_5098),
.A2(n_4995),
.B(n_4978),
.Y(n_5153)
);

INVx2_ASAP7_75t_L g5154 ( 
.A(n_5067),
.Y(n_5154)
);

AOI211xp5_ASAP7_75t_L g5155 ( 
.A1(n_5084),
.A2(n_5024),
.B(n_5010),
.C(n_5009),
.Y(n_5155)
);

INVx2_ASAP7_75t_L g5156 ( 
.A(n_5074),
.Y(n_5156)
);

BUFx6f_ASAP7_75t_L g5157 ( 
.A(n_5107),
.Y(n_5157)
);

AND2x2_ASAP7_75t_L g5158 ( 
.A(n_5125),
.B(n_5043),
.Y(n_5158)
);

AND2x2_ASAP7_75t_L g5159 ( 
.A(n_5125),
.B(n_5026),
.Y(n_5159)
);

NAND2xp5_ASAP7_75t_SL g5160 ( 
.A(n_5075),
.B(n_5088),
.Y(n_5160)
);

NAND4xp25_ASAP7_75t_L g5161 ( 
.A(n_5065),
.B(n_5039),
.C(n_5057),
.D(n_5054),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_5122),
.Y(n_5162)
);

AOI211xp5_ASAP7_75t_L g5163 ( 
.A1(n_5068),
.A2(n_4973),
.B(n_4736),
.C(n_4761),
.Y(n_5163)
);

OAI21x1_ASAP7_75t_L g5164 ( 
.A1(n_5098),
.A2(n_5128),
.B(n_5130),
.Y(n_5164)
);

INVx2_ASAP7_75t_L g5165 ( 
.A(n_5072),
.Y(n_5165)
);

AOI22xp33_ASAP7_75t_L g5166 ( 
.A1(n_5086),
.A2(n_5046),
.B1(n_4996),
.B2(n_5016),
.Y(n_5166)
);

NAND2xp5_ASAP7_75t_L g5167 ( 
.A(n_5091),
.B(n_5044),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_5110),
.Y(n_5168)
);

OAI221xp5_ASAP7_75t_L g5169 ( 
.A1(n_5131),
.A2(n_5128),
.B1(n_5089),
.B2(n_5148),
.C(n_5144),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_L g5170 ( 
.A(n_5143),
.B(n_4862),
.Y(n_5170)
);

INVx2_ASAP7_75t_L g5171 ( 
.A(n_5072),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_5110),
.Y(n_5172)
);

NAND2x1_ASAP7_75t_L g5173 ( 
.A(n_5088),
.B(n_4868),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_5127),
.Y(n_5174)
);

OAI22xp33_ASAP7_75t_L g5175 ( 
.A1(n_5138),
.A2(n_5141),
.B1(n_5129),
.B2(n_5119),
.Y(n_5175)
);

OR2x2_ASAP7_75t_L g5176 ( 
.A(n_5082),
.B(n_4843),
.Y(n_5176)
);

HB1xp67_ASAP7_75t_L g5177 ( 
.A(n_5093),
.Y(n_5177)
);

INVx1_ASAP7_75t_L g5178 ( 
.A(n_5127),
.Y(n_5178)
);

AND2x4_ASAP7_75t_L g5179 ( 
.A(n_5104),
.B(n_5028),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_5112),
.Y(n_5180)
);

AOI21xp5_ASAP7_75t_L g5181 ( 
.A1(n_5096),
.A2(n_4751),
.B(n_4738),
.Y(n_5181)
);

OA21x2_ASAP7_75t_L g5182 ( 
.A1(n_5143),
.A2(n_4924),
.B(n_4943),
.Y(n_5182)
);

A2O1A1Ixp33_ASAP7_75t_L g5183 ( 
.A1(n_5096),
.A2(n_4795),
.B(n_4656),
.C(n_4790),
.Y(n_5183)
);

HB1xp67_ASAP7_75t_L g5184 ( 
.A(n_5069),
.Y(n_5184)
);

AND2x2_ASAP7_75t_L g5185 ( 
.A(n_5073),
.B(n_5028),
.Y(n_5185)
);

AO31x2_ASAP7_75t_L g5186 ( 
.A1(n_5140),
.A2(n_5147),
.A3(n_5139),
.B(n_5136),
.Y(n_5186)
);

INVx2_ASAP7_75t_L g5187 ( 
.A(n_5094),
.Y(n_5187)
);

INVx2_ASAP7_75t_L g5188 ( 
.A(n_5095),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_5114),
.Y(n_5189)
);

OAI21x1_ASAP7_75t_L g5190 ( 
.A1(n_5071),
.A2(n_5146),
.B(n_5092),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_5123),
.Y(n_5191)
);

INVx2_ASAP7_75t_L g5192 ( 
.A(n_5100),
.Y(n_5192)
);

INVxp67_ASAP7_75t_SL g5193 ( 
.A(n_5111),
.Y(n_5193)
);

INVx2_ASAP7_75t_L g5194 ( 
.A(n_5101),
.Y(n_5194)
);

BUFx3_ASAP7_75t_L g5195 ( 
.A(n_5103),
.Y(n_5195)
);

OA21x2_ASAP7_75t_L g5196 ( 
.A1(n_5117),
.A2(n_5081),
.B(n_5135),
.Y(n_5196)
);

AND2x4_ASAP7_75t_L g5197 ( 
.A(n_5097),
.B(n_5135),
.Y(n_5197)
);

BUFx6f_ASAP7_75t_L g5198 ( 
.A(n_5115),
.Y(n_5198)
);

AND2x2_ASAP7_75t_L g5199 ( 
.A(n_5118),
.B(n_4868),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_5077),
.B(n_4870),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_5132),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_5078),
.Y(n_5202)
);

AOI211x1_ASAP7_75t_L g5203 ( 
.A1(n_5116),
.A2(n_4798),
.B(n_4818),
.C(n_4460),
.Y(n_5203)
);

INVx2_ASAP7_75t_L g5204 ( 
.A(n_5083),
.Y(n_5204)
);

AND2x2_ASAP7_75t_L g5205 ( 
.A(n_5158),
.B(n_5152),
.Y(n_5205)
);

AOI22xp33_ASAP7_75t_L g5206 ( 
.A1(n_5161),
.A2(n_5142),
.B1(n_5118),
.B2(n_5066),
.Y(n_5206)
);

AOI221xp5_ASAP7_75t_L g5207 ( 
.A1(n_5155),
.A2(n_5099),
.B1(n_5102),
.B2(n_5126),
.C(n_5108),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_5170),
.Y(n_5208)
);

AND2x2_ASAP7_75t_L g5209 ( 
.A(n_5193),
.B(n_5106),
.Y(n_5209)
);

INVx2_ASAP7_75t_L g5210 ( 
.A(n_5177),
.Y(n_5210)
);

BUFx2_ASAP7_75t_L g5211 ( 
.A(n_5179),
.Y(n_5211)
);

INVx2_ASAP7_75t_L g5212 ( 
.A(n_5150),
.Y(n_5212)
);

NOR2xp33_ASAP7_75t_L g5213 ( 
.A(n_5169),
.B(n_5124),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_5162),
.Y(n_5214)
);

NAND2xp5_ASAP7_75t_L g5215 ( 
.A(n_5167),
.B(n_5087),
.Y(n_5215)
);

OAI221xp5_ASAP7_75t_L g5216 ( 
.A1(n_5149),
.A2(n_5142),
.B1(n_5109),
.B2(n_5120),
.C(n_5133),
.Y(n_5216)
);

NAND2xp5_ASAP7_75t_L g5217 ( 
.A(n_5154),
.B(n_5070),
.Y(n_5217)
);

AND2x2_ASAP7_75t_L g5218 ( 
.A(n_5185),
.B(n_5105),
.Y(n_5218)
);

OR2x2_ASAP7_75t_L g5219 ( 
.A(n_5184),
.B(n_5134),
.Y(n_5219)
);

AOI21xp33_ASAP7_75t_L g5220 ( 
.A1(n_5163),
.A2(n_4838),
.B(n_4776),
.Y(n_5220)
);

AND2x2_ASAP7_75t_L g5221 ( 
.A(n_5197),
.B(n_5145),
.Y(n_5221)
);

OR2x2_ASAP7_75t_L g5222 ( 
.A(n_5176),
.B(n_5137),
.Y(n_5222)
);

AND2x2_ASAP7_75t_L g5223 ( 
.A(n_5196),
.B(n_5113),
.Y(n_5223)
);

NAND3x1_ASAP7_75t_SL g5224 ( 
.A(n_5179),
.B(n_4699),
.C(n_4990),
.Y(n_5224)
);

AND2x4_ASAP7_75t_L g5225 ( 
.A(n_5159),
.B(n_5081),
.Y(n_5225)
);

OR2x6_ASAP7_75t_SL g5226 ( 
.A(n_5151),
.B(n_4477),
.Y(n_5226)
);

AND2x2_ASAP7_75t_L g5227 ( 
.A(n_5196),
.B(n_5166),
.Y(n_5227)
);

INVx2_ASAP7_75t_L g5228 ( 
.A(n_5156),
.Y(n_5228)
);

HB1xp67_ASAP7_75t_L g5229 ( 
.A(n_5186),
.Y(n_5229)
);

NAND2xp5_ASAP7_75t_L g5230 ( 
.A(n_5181),
.B(n_5121),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_5168),
.Y(n_5231)
);

AND2x2_ASAP7_75t_L g5232 ( 
.A(n_5160),
.B(n_5090),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5172),
.Y(n_5233)
);

HB1xp67_ASAP7_75t_L g5234 ( 
.A(n_5186),
.Y(n_5234)
);

AND2x2_ASAP7_75t_L g5235 ( 
.A(n_5190),
.B(n_4874),
.Y(n_5235)
);

BUFx3_ASAP7_75t_L g5236 ( 
.A(n_5195),
.Y(n_5236)
);

AND2x2_ASAP7_75t_L g5237 ( 
.A(n_5199),
.B(n_4877),
.Y(n_5237)
);

AND2x2_ASAP7_75t_L g5238 ( 
.A(n_5153),
.B(n_4882),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_5174),
.Y(n_5239)
);

NAND2xp5_ASAP7_75t_SL g5240 ( 
.A(n_5175),
.B(n_4154),
.Y(n_5240)
);

OR2x2_ASAP7_75t_L g5241 ( 
.A(n_5200),
.B(n_4678),
.Y(n_5241)
);

INVx2_ASAP7_75t_L g5242 ( 
.A(n_5165),
.Y(n_5242)
);

BUFx3_ASAP7_75t_L g5243 ( 
.A(n_5157),
.Y(n_5243)
);

AND2x2_ASAP7_75t_L g5244 ( 
.A(n_5164),
.B(n_4154),
.Y(n_5244)
);

INVx2_ASAP7_75t_L g5245 ( 
.A(n_5171),
.Y(n_5245)
);

NAND2xp5_ASAP7_75t_L g5246 ( 
.A(n_5178),
.B(n_4634),
.Y(n_5246)
);

INVx2_ASAP7_75t_L g5247 ( 
.A(n_5188),
.Y(n_5247)
);

OR2x2_ASAP7_75t_L g5248 ( 
.A(n_5180),
.B(n_4678),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_5189),
.Y(n_5249)
);

INVx2_ASAP7_75t_L g5250 ( 
.A(n_5192),
.Y(n_5250)
);

AND2x4_ASAP7_75t_SL g5251 ( 
.A(n_5157),
.B(n_5198),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_5191),
.Y(n_5252)
);

INVx1_ASAP7_75t_L g5253 ( 
.A(n_5201),
.Y(n_5253)
);

AND2x2_ASAP7_75t_L g5254 ( 
.A(n_5202),
.B(n_4158),
.Y(n_5254)
);

OR2x2_ASAP7_75t_L g5255 ( 
.A(n_5187),
.B(n_4650),
.Y(n_5255)
);

INVx2_ASAP7_75t_L g5256 ( 
.A(n_5194),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_5182),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_5182),
.Y(n_5258)
);

INVx3_ASAP7_75t_L g5259 ( 
.A(n_5173),
.Y(n_5259)
);

OR2x2_ASAP7_75t_L g5260 ( 
.A(n_5210),
.B(n_5204),
.Y(n_5260)
);

AND3x2_ASAP7_75t_L g5261 ( 
.A(n_5213),
.B(n_5203),
.C(n_4792),
.Y(n_5261)
);

INVx1_ASAP7_75t_SL g5262 ( 
.A(n_5251),
.Y(n_5262)
);

AND2x2_ASAP7_75t_L g5263 ( 
.A(n_5211),
.B(n_5173),
.Y(n_5263)
);

NAND2xp5_ASAP7_75t_L g5264 ( 
.A(n_5226),
.B(n_5183),
.Y(n_5264)
);

AND2x2_ASAP7_75t_L g5265 ( 
.A(n_5205),
.B(n_4749),
.Y(n_5265)
);

NAND2xp5_ASAP7_75t_L g5266 ( 
.A(n_5206),
.B(n_4777),
.Y(n_5266)
);

INVx4_ASAP7_75t_L g5267 ( 
.A(n_5243),
.Y(n_5267)
);

AOI22xp33_ASAP7_75t_L g5268 ( 
.A1(n_5227),
.A2(n_4313),
.B1(n_4778),
.B2(n_4803),
.Y(n_5268)
);

OR2x2_ASAP7_75t_L g5269 ( 
.A(n_5214),
.B(n_4788),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_5209),
.Y(n_5270)
);

OR2x2_ASAP7_75t_L g5271 ( 
.A(n_5241),
.B(n_4788),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_5212),
.Y(n_5272)
);

AOI22xp33_ASAP7_75t_L g5273 ( 
.A1(n_5207),
.A2(n_4816),
.B1(n_4812),
.B2(n_4461),
.Y(n_5273)
);

INVx2_ASAP7_75t_L g5274 ( 
.A(n_5219),
.Y(n_5274)
);

NAND2xp5_ASAP7_75t_L g5275 ( 
.A(n_5208),
.B(n_4695),
.Y(n_5275)
);

INVx2_ASAP7_75t_L g5276 ( 
.A(n_5236),
.Y(n_5276)
);

NAND2xp5_ASAP7_75t_L g5277 ( 
.A(n_5208),
.B(n_4695),
.Y(n_5277)
);

NAND2xp5_ASAP7_75t_L g5278 ( 
.A(n_5220),
.B(n_4707),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5217),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_L g5280 ( 
.A(n_5230),
.B(n_5215),
.Y(n_5280)
);

NAND2xp5_ASAP7_75t_L g5281 ( 
.A(n_5232),
.B(n_4707),
.Y(n_5281)
);

OR2x2_ASAP7_75t_L g5282 ( 
.A(n_5248),
.B(n_4758),
.Y(n_5282)
);

AND2x2_ASAP7_75t_L g5283 ( 
.A(n_5223),
.B(n_4327),
.Y(n_5283)
);

AND2x2_ASAP7_75t_L g5284 ( 
.A(n_5225),
.B(n_4231),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_5255),
.Y(n_5285)
);

AND2x2_ASAP7_75t_L g5286 ( 
.A(n_5225),
.B(n_4274),
.Y(n_5286)
);

INVx1_ASAP7_75t_L g5287 ( 
.A(n_5229),
.Y(n_5287)
);

INVx1_ASAP7_75t_L g5288 ( 
.A(n_5249),
.Y(n_5288)
);

AND2x2_ASAP7_75t_L g5289 ( 
.A(n_5244),
.B(n_4208),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_5249),
.Y(n_5290)
);

AND2x2_ASAP7_75t_L g5291 ( 
.A(n_5221),
.B(n_4573),
.Y(n_5291)
);

INVx1_ASAP7_75t_SL g5292 ( 
.A(n_5240),
.Y(n_5292)
);

NAND2xp5_ASAP7_75t_L g5293 ( 
.A(n_5252),
.B(n_4652),
.Y(n_5293)
);

AND2x2_ASAP7_75t_L g5294 ( 
.A(n_5218),
.B(n_4326),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_5252),
.B(n_4659),
.Y(n_5295)
);

OR2x2_ASAP7_75t_L g5296 ( 
.A(n_5253),
.B(n_4595),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_5234),
.Y(n_5297)
);

INVxp67_ASAP7_75t_L g5298 ( 
.A(n_5276),
.Y(n_5298)
);

INVx2_ASAP7_75t_L g5299 ( 
.A(n_5272),
.Y(n_5299)
);

INVx2_ASAP7_75t_L g5300 ( 
.A(n_5267),
.Y(n_5300)
);

HB1xp67_ASAP7_75t_L g5301 ( 
.A(n_5287),
.Y(n_5301)
);

NOR2xp33_ASAP7_75t_L g5302 ( 
.A(n_5267),
.B(n_5216),
.Y(n_5302)
);

OR2x2_ASAP7_75t_L g5303 ( 
.A(n_5296),
.B(n_5246),
.Y(n_5303)
);

INVx2_ASAP7_75t_L g5304 ( 
.A(n_5274),
.Y(n_5304)
);

OR2x6_ASAP7_75t_L g5305 ( 
.A(n_5297),
.B(n_5224),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_5270),
.B(n_5231),
.Y(n_5306)
);

INVx3_ASAP7_75t_L g5307 ( 
.A(n_5262),
.Y(n_5307)
);

INVx3_ASAP7_75t_L g5308 ( 
.A(n_5283),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_5288),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_5288),
.Y(n_5310)
);

INVx2_ASAP7_75t_L g5311 ( 
.A(n_5260),
.Y(n_5311)
);

NAND2xp5_ASAP7_75t_L g5312 ( 
.A(n_5261),
.B(n_5233),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_5290),
.Y(n_5313)
);

AND2x2_ASAP7_75t_L g5314 ( 
.A(n_5292),
.B(n_5238),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_5279),
.B(n_5239),
.Y(n_5315)
);

AND2x2_ASAP7_75t_L g5316 ( 
.A(n_5263),
.B(n_5235),
.Y(n_5316)
);

NAND2xp5_ASAP7_75t_L g5317 ( 
.A(n_5268),
.B(n_5273),
.Y(n_5317)
);

INVx1_ASAP7_75t_L g5318 ( 
.A(n_5290),
.Y(n_5318)
);

OR2x2_ASAP7_75t_L g5319 ( 
.A(n_5271),
.B(n_5228),
.Y(n_5319)
);

AND2x2_ASAP7_75t_L g5320 ( 
.A(n_5265),
.B(n_5237),
.Y(n_5320)
);

NAND2xp5_ASAP7_75t_L g5321 ( 
.A(n_5266),
.B(n_5250),
.Y(n_5321)
);

AND2x2_ASAP7_75t_L g5322 ( 
.A(n_5291),
.B(n_5254),
.Y(n_5322)
);

OR2x2_ASAP7_75t_L g5323 ( 
.A(n_5275),
.B(n_5256),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_5285),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_5295),
.Y(n_5325)
);

OAI22xp33_ASAP7_75t_SL g5326 ( 
.A1(n_5264),
.A2(n_5259),
.B1(n_5257),
.B2(n_5258),
.Y(n_5326)
);

NAND2xp5_ASAP7_75t_L g5327 ( 
.A(n_5280),
.B(n_5247),
.Y(n_5327)
);

INVx3_ASAP7_75t_L g5328 ( 
.A(n_5294),
.Y(n_5328)
);

INVxp67_ASAP7_75t_L g5329 ( 
.A(n_5278),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_5277),
.Y(n_5330)
);

NAND2xp5_ASAP7_75t_L g5331 ( 
.A(n_5281),
.B(n_5242),
.Y(n_5331)
);

AND2x4_ASAP7_75t_L g5332 ( 
.A(n_5307),
.B(n_5284),
.Y(n_5332)
);

INVxp67_ASAP7_75t_L g5333 ( 
.A(n_5307),
.Y(n_5333)
);

AND2x2_ASAP7_75t_L g5334 ( 
.A(n_5300),
.B(n_5286),
.Y(n_5334)
);

AND2x2_ASAP7_75t_L g5335 ( 
.A(n_5298),
.B(n_5289),
.Y(n_5335)
);

AND2x2_ASAP7_75t_L g5336 ( 
.A(n_5314),
.B(n_5282),
.Y(n_5336)
);

INVx2_ASAP7_75t_L g5337 ( 
.A(n_5311),
.Y(n_5337)
);

INVx2_ASAP7_75t_L g5338 ( 
.A(n_5304),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_5301),
.Y(n_5339)
);

INVx1_ASAP7_75t_SL g5340 ( 
.A(n_5299),
.Y(n_5340)
);

INVx4_ASAP7_75t_L g5341 ( 
.A(n_5305),
.Y(n_5341)
);

NAND2xp5_ASAP7_75t_L g5342 ( 
.A(n_5317),
.B(n_5325),
.Y(n_5342)
);

INVx1_ASAP7_75t_SL g5343 ( 
.A(n_5312),
.Y(n_5343)
);

INVx2_ASAP7_75t_L g5344 ( 
.A(n_5319),
.Y(n_5344)
);

OR2x2_ASAP7_75t_L g5345 ( 
.A(n_5327),
.B(n_5269),
.Y(n_5345)
);

AND2x2_ASAP7_75t_L g5346 ( 
.A(n_5316),
.B(n_5293),
.Y(n_5346)
);

AND2x2_ASAP7_75t_L g5347 ( 
.A(n_5308),
.B(n_5245),
.Y(n_5347)
);

AND2x2_ASAP7_75t_L g5348 ( 
.A(n_5308),
.B(n_5328),
.Y(n_5348)
);

AND2x2_ASAP7_75t_L g5349 ( 
.A(n_5320),
.B(n_5222),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_5324),
.Y(n_5350)
);

INVx2_ASAP7_75t_L g5351 ( 
.A(n_5323),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_5306),
.Y(n_5352)
);

INVx1_ASAP7_75t_SL g5353 ( 
.A(n_5302),
.Y(n_5353)
);

INVx1_ASAP7_75t_SL g5354 ( 
.A(n_5315),
.Y(n_5354)
);

INVx2_ASAP7_75t_L g5355 ( 
.A(n_5322),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_5309),
.Y(n_5356)
);

INVx2_ASAP7_75t_L g5357 ( 
.A(n_5303),
.Y(n_5357)
);

AND2x2_ASAP7_75t_L g5358 ( 
.A(n_5330),
.B(n_4717),
.Y(n_5358)
);

INVx2_ASAP7_75t_L g5359 ( 
.A(n_5310),
.Y(n_5359)
);

INVx1_ASAP7_75t_SL g5360 ( 
.A(n_5321),
.Y(n_5360)
);

AOI22xp33_ASAP7_75t_SL g5361 ( 
.A1(n_5326),
.A2(n_4557),
.B1(n_4527),
.B2(n_4520),
.Y(n_5361)
);

NAND2xp5_ASAP7_75t_L g5362 ( 
.A(n_5329),
.B(n_4499),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_5313),
.Y(n_5363)
);

AND2x2_ASAP7_75t_L g5364 ( 
.A(n_5331),
.B(n_4717),
.Y(n_5364)
);

HB1xp67_ASAP7_75t_L g5365 ( 
.A(n_5318),
.Y(n_5365)
);

INVx1_ASAP7_75t_L g5366 ( 
.A(n_5301),
.Y(n_5366)
);

INVx1_ASAP7_75t_L g5367 ( 
.A(n_5307),
.Y(n_5367)
);

NAND2xp5_ASAP7_75t_L g5368 ( 
.A(n_5333),
.B(n_639),
.Y(n_5368)
);

OR2x2_ASAP7_75t_L g5369 ( 
.A(n_5367),
.B(n_640),
.Y(n_5369)
);

NOR2xp33_ASAP7_75t_L g5370 ( 
.A(n_5341),
.B(n_4261),
.Y(n_5370)
);

INVx2_ASAP7_75t_L g5371 ( 
.A(n_5344),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_L g5372 ( 
.A(n_5338),
.B(n_641),
.Y(n_5372)
);

INVx3_ASAP7_75t_L g5373 ( 
.A(n_5332),
.Y(n_5373)
);

INVxp67_ASAP7_75t_SL g5374 ( 
.A(n_5366),
.Y(n_5374)
);

NOR2x1p5_ASAP7_75t_SL g5375 ( 
.A(n_5339),
.B(n_5337),
.Y(n_5375)
);

NAND4xp25_ASAP7_75t_L g5376 ( 
.A(n_5353),
.B(n_4774),
.C(n_4767),
.D(n_4468),
.Y(n_5376)
);

NAND2xp5_ASAP7_75t_L g5377 ( 
.A(n_5360),
.B(n_5336),
.Y(n_5377)
);

INVx2_ASAP7_75t_L g5378 ( 
.A(n_5348),
.Y(n_5378)
);

OR2x2_ASAP7_75t_L g5379 ( 
.A(n_5357),
.B(n_641),
.Y(n_5379)
);

NAND2xp5_ASAP7_75t_L g5380 ( 
.A(n_5340),
.B(n_5347),
.Y(n_5380)
);

NAND2xp5_ASAP7_75t_L g5381 ( 
.A(n_5351),
.B(n_642),
.Y(n_5381)
);

INVx2_ASAP7_75t_SL g5382 ( 
.A(n_5335),
.Y(n_5382)
);

INVx2_ASAP7_75t_L g5383 ( 
.A(n_5334),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_5365),
.Y(n_5384)
);

NAND2xp5_ASAP7_75t_L g5385 ( 
.A(n_5349),
.B(n_642),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_5355),
.Y(n_5386)
);

INVx1_ASAP7_75t_L g5387 ( 
.A(n_5345),
.Y(n_5387)
);

AND2x4_ASAP7_75t_L g5388 ( 
.A(n_5343),
.B(n_4770),
.Y(n_5388)
);

CKINVDCx5p33_ASAP7_75t_R g5389 ( 
.A(n_5354),
.Y(n_5389)
);

INVx1_ASAP7_75t_L g5390 ( 
.A(n_5350),
.Y(n_5390)
);

NAND2xp5_ASAP7_75t_L g5391 ( 
.A(n_5361),
.B(n_642),
.Y(n_5391)
);

HB1xp67_ASAP7_75t_L g5392 ( 
.A(n_5350),
.Y(n_5392)
);

INVx1_ASAP7_75t_L g5393 ( 
.A(n_5356),
.Y(n_5393)
);

INVx2_ASAP7_75t_SL g5394 ( 
.A(n_5346),
.Y(n_5394)
);

INVxp67_ASAP7_75t_L g5395 ( 
.A(n_5342),
.Y(n_5395)
);

INVx2_ASAP7_75t_L g5396 ( 
.A(n_5359),
.Y(n_5396)
);

HB1xp67_ASAP7_75t_L g5397 ( 
.A(n_5356),
.Y(n_5397)
);

AND2x2_ASAP7_75t_L g5398 ( 
.A(n_5364),
.B(n_4619),
.Y(n_5398)
);

NAND2xp5_ASAP7_75t_L g5399 ( 
.A(n_5352),
.B(n_5358),
.Y(n_5399)
);

BUFx2_ASAP7_75t_L g5400 ( 
.A(n_5352),
.Y(n_5400)
);

AND2x4_ASAP7_75t_L g5401 ( 
.A(n_5363),
.B(n_4485),
.Y(n_5401)
);

NAND2xp5_ASAP7_75t_L g5402 ( 
.A(n_5382),
.B(n_5362),
.Y(n_5402)
);

INVx1_ASAP7_75t_L g5403 ( 
.A(n_5371),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_5374),
.Y(n_5404)
);

INVx2_ASAP7_75t_L g5405 ( 
.A(n_5373),
.Y(n_5405)
);

INVx2_ASAP7_75t_L g5406 ( 
.A(n_5383),
.Y(n_5406)
);

NAND2xp5_ASAP7_75t_L g5407 ( 
.A(n_5389),
.B(n_643),
.Y(n_5407)
);

INVx2_ASAP7_75t_L g5408 ( 
.A(n_5378),
.Y(n_5408)
);

NOR2xp33_ASAP7_75t_L g5409 ( 
.A(n_5370),
.B(n_643),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_5385),
.Y(n_5410)
);

OAI221xp5_ASAP7_75t_L g5411 ( 
.A1(n_5394),
.A2(n_4568),
.B1(n_4260),
.B2(n_4286),
.C(n_4267),
.Y(n_5411)
);

A2O1A1Ixp33_ASAP7_75t_L g5412 ( 
.A1(n_5375),
.A2(n_4800),
.B(n_4785),
.C(n_4801),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_5368),
.Y(n_5413)
);

NOR2x1p5_ASAP7_75t_L g5414 ( 
.A(n_5386),
.B(n_4442),
.Y(n_5414)
);

AOI21xp33_ASAP7_75t_SL g5415 ( 
.A1(n_5381),
.A2(n_644),
.B(n_645),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5379),
.Y(n_5416)
);

OAI22xp33_ASAP7_75t_L g5417 ( 
.A1(n_5399),
.A2(n_5391),
.B1(n_5369),
.B2(n_5387),
.Y(n_5417)
);

NAND2xp5_ASAP7_75t_L g5418 ( 
.A(n_5401),
.B(n_644),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_5372),
.Y(n_5419)
);

OAI21xp33_ASAP7_75t_L g5420 ( 
.A1(n_5395),
.A2(n_4335),
.B(n_4748),
.Y(n_5420)
);

OAI322xp33_ASAP7_75t_L g5421 ( 
.A1(n_5384),
.A2(n_4447),
.A3(n_4442),
.B1(n_4556),
.B2(n_646),
.C1(n_650),
.C2(n_649),
.Y(n_5421)
);

AOI21xp5_ASAP7_75t_L g5422 ( 
.A1(n_5392),
.A2(n_5396),
.B(n_5397),
.Y(n_5422)
);

INVxp67_ASAP7_75t_L g5423 ( 
.A(n_5400),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_5390),
.Y(n_5424)
);

INVx1_ASAP7_75t_SL g5425 ( 
.A(n_5388),
.Y(n_5425)
);

OAI21xp33_ASAP7_75t_SL g5426 ( 
.A1(n_5393),
.A2(n_5398),
.B(n_5376),
.Y(n_5426)
);

AOI21xp33_ASAP7_75t_SL g5427 ( 
.A1(n_5388),
.A2(n_648),
.B(n_646),
.Y(n_5427)
);

INVx1_ASAP7_75t_L g5428 ( 
.A(n_5371),
.Y(n_5428)
);

INVx2_ASAP7_75t_L g5429 ( 
.A(n_5373),
.Y(n_5429)
);

AOI21xp5_ASAP7_75t_L g5430 ( 
.A1(n_5377),
.A2(n_4745),
.B(n_4685),
.Y(n_5430)
);

AND2x2_ASAP7_75t_L g5431 ( 
.A(n_5382),
.B(n_645),
.Y(n_5431)
);

AOI22xp33_ASAP7_75t_L g5432 ( 
.A1(n_5373),
.A2(n_4447),
.B1(n_4556),
.B2(n_4647),
.Y(n_5432)
);

HB1xp67_ASAP7_75t_L g5433 ( 
.A(n_5371),
.Y(n_5433)
);

OR2x2_ASAP7_75t_L g5434 ( 
.A(n_5385),
.B(n_645),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5371),
.Y(n_5435)
);

AOI22xp5_ASAP7_75t_L g5436 ( 
.A1(n_5370),
.A2(n_4720),
.B1(n_4743),
.B2(n_4727),
.Y(n_5436)
);

INVxp67_ASAP7_75t_L g5437 ( 
.A(n_5380),
.Y(n_5437)
);

AOI22xp33_ASAP7_75t_L g5438 ( 
.A1(n_5373),
.A2(n_4590),
.B1(n_4357),
.B2(n_4247),
.Y(n_5438)
);

OR2x2_ASAP7_75t_L g5439 ( 
.A(n_5385),
.B(n_646),
.Y(n_5439)
);

NAND2x1_ASAP7_75t_L g5440 ( 
.A(n_5373),
.B(n_4357),
.Y(n_5440)
);

AOI22xp5_ASAP7_75t_L g5441 ( 
.A1(n_5370),
.A2(n_4633),
.B1(n_4643),
.B2(n_4706),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_5371),
.Y(n_5442)
);

AOI21xp5_ASAP7_75t_L g5443 ( 
.A1(n_5377),
.A2(n_4671),
.B(n_4668),
.Y(n_5443)
);

INVxp67_ASAP7_75t_L g5444 ( 
.A(n_5433),
.Y(n_5444)
);

INVx1_ASAP7_75t_L g5445 ( 
.A(n_5407),
.Y(n_5445)
);

INVx1_ASAP7_75t_SL g5446 ( 
.A(n_5405),
.Y(n_5446)
);

AND2x2_ASAP7_75t_L g5447 ( 
.A(n_5431),
.B(n_5408),
.Y(n_5447)
);

NAND2xp5_ASAP7_75t_L g5448 ( 
.A(n_5429),
.B(n_5403),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_5428),
.Y(n_5449)
);

AND2x2_ASAP7_75t_L g5450 ( 
.A(n_5406),
.B(n_649),
.Y(n_5450)
);

INVx1_ASAP7_75t_L g5451 ( 
.A(n_5435),
.Y(n_5451)
);

NAND2xp5_ASAP7_75t_SL g5452 ( 
.A(n_5427),
.B(n_4244),
.Y(n_5452)
);

INVx1_ASAP7_75t_L g5453 ( 
.A(n_5442),
.Y(n_5453)
);

NAND2xp5_ASAP7_75t_L g5454 ( 
.A(n_5404),
.B(n_649),
.Y(n_5454)
);

AO22x1_ASAP7_75t_L g5455 ( 
.A1(n_5409),
.A2(n_4547),
.B1(n_4283),
.B2(n_4287),
.Y(n_5455)
);

OR2x2_ASAP7_75t_L g5456 ( 
.A(n_5425),
.B(n_650),
.Y(n_5456)
);

NAND2xp5_ASAP7_75t_L g5457 ( 
.A(n_5437),
.B(n_651),
.Y(n_5457)
);

AND3x2_ASAP7_75t_L g5458 ( 
.A(n_5423),
.B(n_651),
.C(n_652),
.Y(n_5458)
);

NOR2xp33_ASAP7_75t_L g5459 ( 
.A(n_5426),
.B(n_652),
.Y(n_5459)
);

INVx1_ASAP7_75t_SL g5460 ( 
.A(n_5418),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_5402),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_5434),
.Y(n_5462)
);

INVx1_ASAP7_75t_SL g5463 ( 
.A(n_5439),
.Y(n_5463)
);

NAND2xp5_ASAP7_75t_SL g5464 ( 
.A(n_5417),
.B(n_4282),
.Y(n_5464)
);

INVx1_ASAP7_75t_L g5465 ( 
.A(n_5416),
.Y(n_5465)
);

OAI22xp5_ASAP7_75t_L g5466 ( 
.A1(n_5411),
.A2(n_4547),
.B1(n_4411),
.B2(n_4465),
.Y(n_5466)
);

AND2x2_ASAP7_75t_L g5467 ( 
.A(n_5410),
.B(n_653),
.Y(n_5467)
);

INVx1_ASAP7_75t_L g5468 ( 
.A(n_5422),
.Y(n_5468)
);

INVx2_ASAP7_75t_L g5469 ( 
.A(n_5414),
.Y(n_5469)
);

NAND2xp5_ASAP7_75t_L g5470 ( 
.A(n_5430),
.B(n_653),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_5421),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_5424),
.Y(n_5472)
);

NAND2xp5_ASAP7_75t_L g5473 ( 
.A(n_5443),
.B(n_653),
.Y(n_5473)
);

NAND3xp33_ASAP7_75t_L g5474 ( 
.A(n_5413),
.B(n_654),
.C(n_655),
.Y(n_5474)
);

INVx1_ASAP7_75t_L g5475 ( 
.A(n_5419),
.Y(n_5475)
);

NAND2xp5_ASAP7_75t_L g5476 ( 
.A(n_5415),
.B(n_654),
.Y(n_5476)
);

NAND2xp5_ASAP7_75t_L g5477 ( 
.A(n_5415),
.B(n_654),
.Y(n_5477)
);

OAI221xp5_ASAP7_75t_SL g5478 ( 
.A1(n_5420),
.A2(n_657),
.B1(n_655),
.B2(n_656),
.C(n_658),
.Y(n_5478)
);

NAND2xp5_ASAP7_75t_L g5479 ( 
.A(n_5432),
.B(n_655),
.Y(n_5479)
);

NAND2xp5_ASAP7_75t_L g5480 ( 
.A(n_5412),
.B(n_656),
.Y(n_5480)
);

NOR2xp33_ASAP7_75t_L g5481 ( 
.A(n_5446),
.B(n_5440),
.Y(n_5481)
);

NAND2xp5_ASAP7_75t_L g5482 ( 
.A(n_5459),
.B(n_5436),
.Y(n_5482)
);

NAND2xp5_ASAP7_75t_L g5483 ( 
.A(n_5468),
.B(n_5471),
.Y(n_5483)
);

INVx1_ASAP7_75t_L g5484 ( 
.A(n_5450),
.Y(n_5484)
);

NAND2xp5_ASAP7_75t_L g5485 ( 
.A(n_5444),
.B(n_5438),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_5447),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_5456),
.Y(n_5487)
);

NAND2xp5_ASAP7_75t_SL g5488 ( 
.A(n_5474),
.B(n_5441),
.Y(n_5488)
);

CKINVDCx5p33_ASAP7_75t_R g5489 ( 
.A(n_5461),
.Y(n_5489)
);

NAND2xp5_ASAP7_75t_L g5490 ( 
.A(n_5449),
.B(n_657),
.Y(n_5490)
);

AND2x2_ASAP7_75t_L g5491 ( 
.A(n_5467),
.B(n_657),
.Y(n_5491)
);

NAND2xp5_ASAP7_75t_L g5492 ( 
.A(n_5451),
.B(n_658),
.Y(n_5492)
);

INVx2_ASAP7_75t_L g5493 ( 
.A(n_5453),
.Y(n_5493)
);

NOR2xp33_ASAP7_75t_L g5494 ( 
.A(n_5476),
.B(n_658),
.Y(n_5494)
);

INVx1_ASAP7_75t_L g5495 ( 
.A(n_5479),
.Y(n_5495)
);

NAND2xp5_ASAP7_75t_L g5496 ( 
.A(n_5463),
.B(n_659),
.Y(n_5496)
);

AND2x2_ASAP7_75t_L g5497 ( 
.A(n_5469),
.B(n_659),
.Y(n_5497)
);

NOR2xp33_ASAP7_75t_L g5498 ( 
.A(n_5477),
.B(n_660),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5454),
.Y(n_5499)
);

OR2x2_ASAP7_75t_L g5500 ( 
.A(n_5457),
.B(n_660),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_L g5501 ( 
.A(n_5462),
.B(n_5460),
.Y(n_5501)
);

NAND2xp5_ASAP7_75t_L g5502 ( 
.A(n_5445),
.B(n_660),
.Y(n_5502)
);

INVx2_ASAP7_75t_L g5503 ( 
.A(n_5465),
.Y(n_5503)
);

NAND2xp5_ASAP7_75t_L g5504 ( 
.A(n_5474),
.B(n_661),
.Y(n_5504)
);

AND2x2_ASAP7_75t_L g5505 ( 
.A(n_5464),
.B(n_662),
.Y(n_5505)
);

INVx2_ASAP7_75t_L g5506 ( 
.A(n_5452),
.Y(n_5506)
);

NAND2xp5_ASAP7_75t_L g5507 ( 
.A(n_5470),
.B(n_662),
.Y(n_5507)
);

AND2x2_ASAP7_75t_L g5508 ( 
.A(n_5475),
.B(n_663),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_5473),
.Y(n_5509)
);

NAND2xp5_ASAP7_75t_L g5510 ( 
.A(n_5480),
.B(n_5472),
.Y(n_5510)
);

INVx2_ASAP7_75t_L g5511 ( 
.A(n_5455),
.Y(n_5511)
);

NOR2x1_ASAP7_75t_L g5512 ( 
.A(n_5478),
.B(n_663),
.Y(n_5512)
);

OR2x2_ASAP7_75t_L g5513 ( 
.A(n_5466),
.B(n_664),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_5448),
.Y(n_5514)
);

NAND2xp5_ASAP7_75t_L g5515 ( 
.A(n_5458),
.B(n_664),
.Y(n_5515)
);

OR2x2_ASAP7_75t_L g5516 ( 
.A(n_5446),
.B(n_665),
.Y(n_5516)
);

NAND2xp5_ASAP7_75t_L g5517 ( 
.A(n_5497),
.B(n_665),
.Y(n_5517)
);

NAND2xp5_ASAP7_75t_L g5518 ( 
.A(n_5491),
.B(n_665),
.Y(n_5518)
);

NAND3xp33_ASAP7_75t_SL g5519 ( 
.A(n_5483),
.B(n_5489),
.C(n_5515),
.Y(n_5519)
);

NAND2xp5_ASAP7_75t_SL g5520 ( 
.A(n_5512),
.B(n_4282),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_5505),
.Y(n_5521)
);

AND2x2_ASAP7_75t_L g5522 ( 
.A(n_5486),
.B(n_666),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_5516),
.Y(n_5523)
);

NAND2xp5_ASAP7_75t_L g5524 ( 
.A(n_5481),
.B(n_666),
.Y(n_5524)
);

AND5x1_ASAP7_75t_L g5525 ( 
.A(n_5494),
.B(n_669),
.C(n_667),
.D(n_668),
.E(n_670),
.Y(n_5525)
);

AOI211xp5_ASAP7_75t_L g5526 ( 
.A1(n_5514),
.A2(n_4663),
.B(n_4814),
.C(n_4811),
.Y(n_5526)
);

AOI211xp5_ASAP7_75t_L g5527 ( 
.A1(n_5498),
.A2(n_671),
.B(n_669),
.C(n_670),
.Y(n_5527)
);

NOR2xp67_ASAP7_75t_L g5528 ( 
.A(n_5511),
.B(n_670),
.Y(n_5528)
);

NAND2xp5_ASAP7_75t_L g5529 ( 
.A(n_5508),
.B(n_5512),
.Y(n_5529)
);

NAND4xp75_ASAP7_75t_L g5530 ( 
.A(n_5496),
.B(n_673),
.C(n_671),
.D(n_672),
.Y(n_5530)
);

OR2x2_ASAP7_75t_L g5531 ( 
.A(n_5485),
.B(n_671),
.Y(n_5531)
);

AND2x2_ASAP7_75t_L g5532 ( 
.A(n_5484),
.B(n_672),
.Y(n_5532)
);

AND4x1_ASAP7_75t_L g5533 ( 
.A(n_5507),
.B(n_5501),
.C(n_5504),
.D(n_5487),
.Y(n_5533)
);

NOR2xp33_ASAP7_75t_L g5534 ( 
.A(n_5506),
.B(n_672),
.Y(n_5534)
);

AO21x1_ASAP7_75t_L g5535 ( 
.A1(n_5490),
.A2(n_4688),
.B(n_673),
.Y(n_5535)
);

NAND2xp5_ASAP7_75t_L g5536 ( 
.A(n_5493),
.B(n_674),
.Y(n_5536)
);

INVx2_ASAP7_75t_L g5537 ( 
.A(n_5513),
.Y(n_5537)
);

NOR4xp25_ASAP7_75t_SL g5538 ( 
.A(n_5488),
.B(n_677),
.C(n_675),
.D(n_676),
.Y(n_5538)
);

NOR3xp33_ASAP7_75t_L g5539 ( 
.A(n_5503),
.B(n_675),
.C(n_677),
.Y(n_5539)
);

NAND2xp5_ASAP7_75t_L g5540 ( 
.A(n_5509),
.B(n_677),
.Y(n_5540)
);

NOR3xp33_ASAP7_75t_L g5541 ( 
.A(n_5492),
.B(n_678),
.C(n_679),
.Y(n_5541)
);

NOR3xp33_ASAP7_75t_L g5542 ( 
.A(n_5502),
.B(n_678),
.C(n_680),
.Y(n_5542)
);

NOR2xp33_ASAP7_75t_L g5543 ( 
.A(n_5482),
.B(n_678),
.Y(n_5543)
);

NAND2xp5_ASAP7_75t_SL g5544 ( 
.A(n_5510),
.B(n_4320),
.Y(n_5544)
);

NAND4xp25_ASAP7_75t_L g5545 ( 
.A(n_5495),
.B(n_682),
.C(n_680),
.D(n_681),
.Y(n_5545)
);

NOR3x1_ASAP7_75t_L g5546 ( 
.A(n_5500),
.B(n_4632),
.C(n_680),
.Y(n_5546)
);

NAND2xp5_ASAP7_75t_SL g5547 ( 
.A(n_5499),
.B(n_4328),
.Y(n_5547)
);

INVxp67_ASAP7_75t_L g5548 ( 
.A(n_5481),
.Y(n_5548)
);

AOI21xp33_ASAP7_75t_L g5549 ( 
.A1(n_5543),
.A2(n_681),
.B(n_682),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_5524),
.Y(n_5550)
);

O2A1O1Ixp33_ASAP7_75t_L g5551 ( 
.A1(n_5548),
.A2(n_684),
.B(n_681),
.C(n_683),
.Y(n_5551)
);

AOI221xp5_ASAP7_75t_L g5552 ( 
.A1(n_5545),
.A2(n_4328),
.B1(n_687),
.B2(n_685),
.C(n_686),
.Y(n_5552)
);

NOR2xp33_ASAP7_75t_L g5553 ( 
.A(n_5517),
.B(n_685),
.Y(n_5553)
);

OAI21xp5_ASAP7_75t_L g5554 ( 
.A1(n_5520),
.A2(n_4644),
.B(n_4636),
.Y(n_5554)
);

OAI211xp5_ASAP7_75t_L g5555 ( 
.A1(n_5527),
.A2(n_689),
.B(n_687),
.C(n_688),
.Y(n_5555)
);

XOR2xp5_ASAP7_75t_L g5556 ( 
.A(n_5530),
.B(n_689),
.Y(n_5556)
);

NOR2xp33_ASAP7_75t_R g5557 ( 
.A(n_5519),
.B(n_690),
.Y(n_5557)
);

AOI22xp33_ASAP7_75t_SL g5558 ( 
.A1(n_5522),
.A2(n_4369),
.B1(n_4626),
.B2(n_4617),
.Y(n_5558)
);

AOI221xp5_ASAP7_75t_L g5559 ( 
.A1(n_5539),
.A2(n_692),
.B1(n_690),
.B2(n_691),
.C(n_693),
.Y(n_5559)
);

INVxp67_ASAP7_75t_L g5560 ( 
.A(n_5534),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_5531),
.Y(n_5561)
);

AOI211x1_ASAP7_75t_SL g5562 ( 
.A1(n_5528),
.A2(n_5529),
.B(n_5537),
.C(n_5544),
.Y(n_5562)
);

AOI221xp5_ASAP7_75t_SL g5563 ( 
.A1(n_5547),
.A2(n_696),
.B1(n_694),
.B2(n_695),
.C(n_697),
.Y(n_5563)
);

AOI221xp5_ASAP7_75t_L g5564 ( 
.A1(n_5542),
.A2(n_696),
.B1(n_694),
.B2(n_695),
.C(n_697),
.Y(n_5564)
);

O2A1O1Ixp33_ASAP7_75t_L g5565 ( 
.A1(n_5536),
.A2(n_698),
.B(n_695),
.C(n_697),
.Y(n_5565)
);

AOI221xp5_ASAP7_75t_L g5566 ( 
.A1(n_5541),
.A2(n_700),
.B1(n_698),
.B2(n_699),
.C(n_701),
.Y(n_5566)
);

OAI211xp5_ASAP7_75t_L g5567 ( 
.A1(n_5518),
.A2(n_5538),
.B(n_5540),
.C(n_5523),
.Y(n_5567)
);

CKINVDCx5p33_ASAP7_75t_R g5568 ( 
.A(n_5532),
.Y(n_5568)
);

AOI321xp33_ASAP7_75t_L g5569 ( 
.A1(n_5521),
.A2(n_702),
.A3(n_704),
.B1(n_700),
.B2(n_701),
.C(n_703),
.Y(n_5569)
);

NOR2xp33_ASAP7_75t_R g5570 ( 
.A(n_5525),
.B(n_704),
.Y(n_5570)
);

OAI21xp5_ASAP7_75t_L g5571 ( 
.A1(n_5533),
.A2(n_704),
.B(n_705),
.Y(n_5571)
);

AOI21xp33_ASAP7_75t_SL g5572 ( 
.A1(n_5546),
.A2(n_705),
.B(n_706),
.Y(n_5572)
);

O2A1O1Ixp33_ASAP7_75t_L g5573 ( 
.A1(n_5535),
.A2(n_708),
.B(n_706),
.C(n_707),
.Y(n_5573)
);

NAND2xp5_ASAP7_75t_L g5574 ( 
.A(n_5526),
.B(n_707),
.Y(n_5574)
);

XNOR2xp5_ASAP7_75t_L g5575 ( 
.A(n_5556),
.B(n_708),
.Y(n_5575)
);

AOI211xp5_ASAP7_75t_L g5576 ( 
.A1(n_5549),
.A2(n_713),
.B(n_710),
.C(n_712),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_5551),
.Y(n_5577)
);

AOI221xp5_ASAP7_75t_L g5578 ( 
.A1(n_5572),
.A2(n_5552),
.B1(n_5565),
.B2(n_5559),
.C(n_5573),
.Y(n_5578)
);

AOI221x1_ASAP7_75t_L g5579 ( 
.A1(n_5571),
.A2(n_5550),
.B1(n_5561),
.B2(n_5553),
.C(n_5574),
.Y(n_5579)
);

XNOR2x2_ASAP7_75t_L g5580 ( 
.A(n_5564),
.B(n_714),
.Y(n_5580)
);

AOI221xp5_ASAP7_75t_L g5581 ( 
.A1(n_5566),
.A2(n_717),
.B1(n_715),
.B2(n_716),
.C(n_718),
.Y(n_5581)
);

AOI211xp5_ASAP7_75t_L g5582 ( 
.A1(n_5555),
.A2(n_717),
.B(n_715),
.C(n_716),
.Y(n_5582)
);

AOI221x1_ASAP7_75t_L g5583 ( 
.A1(n_5557),
.A2(n_720),
.B1(n_718),
.B2(n_719),
.C(n_721),
.Y(n_5583)
);

AOI221xp5_ASAP7_75t_L g5584 ( 
.A1(n_5563),
.A2(n_721),
.B1(n_719),
.B2(n_720),
.C(n_722),
.Y(n_5584)
);

AOI221xp5_ASAP7_75t_L g5585 ( 
.A1(n_5560),
.A2(n_722),
.B1(n_723),
.B2(n_790),
.C(n_791),
.Y(n_5585)
);

BUFx6f_ASAP7_75t_L g5586 ( 
.A(n_5568),
.Y(n_5586)
);

AOI21xp5_ASAP7_75t_L g5587 ( 
.A1(n_5567),
.A2(n_723),
.B(n_791),
.Y(n_5587)
);

INVx1_ASAP7_75t_L g5588 ( 
.A(n_5569),
.Y(n_5588)
);

AOI221xp5_ASAP7_75t_L g5589 ( 
.A1(n_5570),
.A2(n_794),
.B1(n_792),
.B2(n_793),
.C(n_795),
.Y(n_5589)
);

NAND4xp25_ASAP7_75t_L g5590 ( 
.A(n_5562),
.B(n_796),
.C(n_794),
.D(n_795),
.Y(n_5590)
);

OAI22x1_ASAP7_75t_L g5591 ( 
.A1(n_5558),
.A2(n_5554),
.B1(n_799),
.B2(n_796),
.Y(n_5591)
);

AND2x2_ASAP7_75t_L g5592 ( 
.A(n_5588),
.B(n_797),
.Y(n_5592)
);

AND2x2_ASAP7_75t_L g5593 ( 
.A(n_5577),
.B(n_797),
.Y(n_5593)
);

AOI21xp5_ASAP7_75t_L g5594 ( 
.A1(n_5587),
.A2(n_800),
.B(n_801),
.Y(n_5594)
);

NAND2x1p5_ASAP7_75t_L g5595 ( 
.A(n_5586),
.B(n_802),
.Y(n_5595)
);

OR2x2_ASAP7_75t_L g5596 ( 
.A(n_5590),
.B(n_803),
.Y(n_5596)
);

XNOR2xp5_ASAP7_75t_L g5597 ( 
.A(n_5575),
.B(n_805),
.Y(n_5597)
);

AOI22xp5_ASAP7_75t_L g5598 ( 
.A1(n_5578),
.A2(n_4501),
.B1(n_4416),
.B2(n_807),
.Y(n_5598)
);

AND3x1_ASAP7_75t_L g5599 ( 
.A(n_5589),
.B(n_808),
.C(n_809),
.Y(n_5599)
);

AOI22xp33_ASAP7_75t_L g5600 ( 
.A1(n_5584),
.A2(n_4416),
.B1(n_4501),
.B2(n_810),
.Y(n_5600)
);

OAI321xp33_ASAP7_75t_L g5601 ( 
.A1(n_5582),
.A2(n_810),
.A3(n_812),
.B1(n_808),
.B2(n_809),
.C(n_811),
.Y(n_5601)
);

OAI221xp5_ASAP7_75t_SL g5602 ( 
.A1(n_5581),
.A2(n_814),
.B1(n_811),
.B2(n_813),
.C(n_815),
.Y(n_5602)
);

AOI21xp5_ASAP7_75t_L g5603 ( 
.A1(n_5591),
.A2(n_813),
.B(n_814),
.Y(n_5603)
);

AOI32xp33_ASAP7_75t_L g5604 ( 
.A1(n_5576),
.A2(n_817),
.A3(n_815),
.B1(n_816),
.B2(n_818),
.Y(n_5604)
);

AOI221x1_ASAP7_75t_L g5605 ( 
.A1(n_5586),
.A2(n_821),
.B1(n_818),
.B2(n_819),
.C(n_822),
.Y(n_5605)
);

AOI32xp33_ASAP7_75t_L g5606 ( 
.A1(n_5585),
.A2(n_822),
.A3(n_819),
.B1(n_821),
.B2(n_823),
.Y(n_5606)
);

AND2x2_ASAP7_75t_L g5607 ( 
.A(n_5586),
.B(n_824),
.Y(n_5607)
);

AND2x2_ASAP7_75t_L g5608 ( 
.A(n_5592),
.B(n_5580),
.Y(n_5608)
);

OR2x2_ASAP7_75t_L g5609 ( 
.A(n_5596),
.B(n_5583),
.Y(n_5609)
);

AND2x2_ASAP7_75t_L g5610 ( 
.A(n_5593),
.B(n_5579),
.Y(n_5610)
);

NAND2xp33_ASAP7_75t_SL g5611 ( 
.A(n_5597),
.B(n_5607),
.Y(n_5611)
);

NAND3xp33_ASAP7_75t_L g5612 ( 
.A(n_5604),
.B(n_825),
.C(n_826),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_5595),
.Y(n_5613)
);

OR2x2_ASAP7_75t_L g5614 ( 
.A(n_5602),
.B(n_826),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_5599),
.Y(n_5615)
);

AOI22xp5_ASAP7_75t_L g5616 ( 
.A1(n_5600),
.A2(n_4501),
.B1(n_830),
.B2(n_827),
.Y(n_5616)
);

AOI22xp5_ASAP7_75t_L g5617 ( 
.A1(n_5598),
.A2(n_4501),
.B1(n_832),
.B2(n_829),
.Y(n_5617)
);

NAND3xp33_ASAP7_75t_SL g5618 ( 
.A(n_5606),
.B(n_831),
.C(n_833),
.Y(n_5618)
);

AND4x2_ASAP7_75t_L g5619 ( 
.A(n_5594),
.B(n_835),
.C(n_831),
.D(n_834),
.Y(n_5619)
);

HB1xp67_ASAP7_75t_L g5620 ( 
.A(n_5605),
.Y(n_5620)
);

NOR3x1_ASAP7_75t_L g5621 ( 
.A(n_5601),
.B(n_834),
.C(n_835),
.Y(n_5621)
);

BUFx2_ASAP7_75t_L g5622 ( 
.A(n_5610),
.Y(n_5622)
);

NAND2xp5_ASAP7_75t_L g5623 ( 
.A(n_5608),
.B(n_5603),
.Y(n_5623)
);

BUFx2_ASAP7_75t_L g5624 ( 
.A(n_5609),
.Y(n_5624)
);

INVx1_ASAP7_75t_SL g5625 ( 
.A(n_5611),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_5614),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5619),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_5622),
.Y(n_5628)
);

OA21x2_ASAP7_75t_L g5629 ( 
.A1(n_5623),
.A2(n_5615),
.B(n_5613),
.Y(n_5629)
);

AND2x4_ASAP7_75t_L g5630 ( 
.A(n_5624),
.B(n_5620),
.Y(n_5630)
);

OAI22xp5_ASAP7_75t_L g5631 ( 
.A1(n_5626),
.A2(n_5612),
.B1(n_5616),
.B2(n_5617),
.Y(n_5631)
);

INVx2_ASAP7_75t_L g5632 ( 
.A(n_5627),
.Y(n_5632)
);

OAI22xp5_ASAP7_75t_SL g5633 ( 
.A1(n_5625),
.A2(n_5621),
.B1(n_5618),
.B2(n_838),
.Y(n_5633)
);

HB1xp67_ASAP7_75t_L g5634 ( 
.A(n_5622),
.Y(n_5634)
);

AOI21xp5_ASAP7_75t_L g5635 ( 
.A1(n_5623),
.A2(n_837),
.B(n_839),
.Y(n_5635)
);

OA22x2_ASAP7_75t_L g5636 ( 
.A1(n_5628),
.A2(n_843),
.B1(n_841),
.B2(n_842),
.Y(n_5636)
);

AND2x4_ASAP7_75t_L g5637 ( 
.A(n_5630),
.B(n_841),
.Y(n_5637)
);

OAI221xp5_ASAP7_75t_L g5638 ( 
.A1(n_5634),
.A2(n_845),
.B1(n_842),
.B2(n_844),
.C(n_846),
.Y(n_5638)
);

NAND2xp5_ASAP7_75t_L g5639 ( 
.A(n_5635),
.B(n_844),
.Y(n_5639)
);

INVx2_ASAP7_75t_L g5640 ( 
.A(n_5636),
.Y(n_5640)
);

OAI22xp5_ASAP7_75t_L g5641 ( 
.A1(n_5640),
.A2(n_5632),
.B1(n_5629),
.B2(n_5639),
.Y(n_5641)
);

AOI21xp5_ASAP7_75t_L g5642 ( 
.A1(n_5641),
.A2(n_5633),
.B(n_5631),
.Y(n_5642)
);

INVx4_ASAP7_75t_L g5643 ( 
.A(n_5642),
.Y(n_5643)
);

AOI21xp33_ASAP7_75t_SL g5644 ( 
.A1(n_5643),
.A2(n_5637),
.B(n_5638),
.Y(n_5644)
);

AOI22xp5_ASAP7_75t_SL g5645 ( 
.A1(n_5644),
.A2(n_853),
.B1(n_847),
.B2(n_850),
.Y(n_5645)
);

OA22x2_ASAP7_75t_L g5646 ( 
.A1(n_5645),
.A2(n_857),
.B1(n_855),
.B2(n_856),
.Y(n_5646)
);

AOI221xp5_ASAP7_75t_L g5647 ( 
.A1(n_5646),
.A2(n_861),
.B1(n_859),
.B2(n_860),
.C(n_862),
.Y(n_5647)
);

AOI211xp5_ASAP7_75t_L g5648 ( 
.A1(n_5647),
.A2(n_865),
.B(n_863),
.C(n_864),
.Y(n_5648)
);


endmodule