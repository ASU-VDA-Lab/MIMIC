module fake_jpeg_2013_n_147 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_147);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVxp33_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_R g60 ( 
.A(n_36),
.B(n_49),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx2_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_10),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_14),
.B(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_48),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_2),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_31),
.A2(n_16),
.B1(n_20),
.B2(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_51),
.A2(n_57),
.B1(n_61),
.B2(n_73),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_55),
.B(n_71),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_16),
.B1(n_20),
.B2(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_27),
.B1(n_21),
.B2(n_24),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_27),
.B1(n_23),
.B2(n_24),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_23),
.B1(n_3),
.B2(n_4),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

AOI22x1_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_32),
.B(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_76),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_38),
.A2(n_32),
.B1(n_37),
.B2(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_5),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_87),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_39),
.C(n_8),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_91),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_39),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_66),
.B(n_54),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_60),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_SL g98 ( 
.A(n_92),
.B(n_94),
.C(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_84),
.B1(n_92),
.B2(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_62),
.B1(n_73),
.B2(n_64),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_80),
.B1(n_94),
.B2(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_102),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_60),
.B(n_71),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_68),
.B(n_54),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_68),
.B(n_74),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_109),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_80),
.B(n_85),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_119),
.B1(n_77),
.B2(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_113),
.B(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_78),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_67),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_104),
.B(n_102),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_101),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_121),
.C(n_118),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_99),
.B1(n_98),
.B2(n_103),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_105),
.B(n_107),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_98),
.B1(n_90),
.B2(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_69),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_126),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_133),
.A2(n_135),
.B(n_85),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_115),
.C(n_111),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_83),
.C(n_74),
.Y(n_138)
);

AO221x1_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_119),
.B1(n_113),
.B2(n_82),
.C(n_112),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_90),
.B1(n_125),
.B2(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_131),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_139),
.C(n_134),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_141),
.A2(n_142),
.B(n_138),
.Y(n_144)
);

XNOR2x2_ASAP7_75t_SL g143 ( 
.A(n_140),
.B(n_139),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_143),
.A2(n_144),
.B(n_132),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_95),
.B(n_69),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_52),
.Y(n_147)
);


endmodule