module real_aes_7817_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_1), .A2(n_146), .B(n_151), .C(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g258 ( .A(n_2), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_3), .A2(n_141), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_4), .B(n_218), .Y(n_467) );
AOI21xp33_ASAP7_75t_L g219 ( .A1(n_5), .A2(n_141), .B(n_220), .Y(n_219) );
AND2x6_ASAP7_75t_L g146 ( .A(n_6), .B(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_7), .A2(n_140), .B(n_148), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_8), .B(n_40), .Y(n_112) );
INVx1_ASAP7_75t_L g556 ( .A(n_9), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_10), .B(n_190), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_11), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g225 ( .A(n_12), .Y(n_225) );
INVx1_ASAP7_75t_L g138 ( .A(n_13), .Y(n_138) );
INVx1_ASAP7_75t_L g158 ( .A(n_14), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_15), .A2(n_159), .B(n_173), .C(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_16), .B(n_218), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_17), .B(n_175), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_18), .B(n_141), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_19), .B(n_480), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_20), .A2(n_206), .B(n_232), .C(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_21), .B(n_218), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_22), .B(n_190), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_23), .A2(n_155), .B(n_157), .C(n_159), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_24), .B(n_190), .Y(n_453) );
CKINVDCx16_ASAP7_75t_R g484 ( .A(n_25), .Y(n_484) );
INVx1_ASAP7_75t_L g452 ( .A(n_26), .Y(n_452) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_27), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_28), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_29), .B(n_190), .Y(n_259) );
INVx1_ASAP7_75t_L g477 ( .A(n_30), .Y(n_477) );
INVx1_ASAP7_75t_L g237 ( .A(n_31), .Y(n_237) );
INVx2_ASAP7_75t_L g144 ( .A(n_32), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_33), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_34), .A2(n_206), .B(n_226), .C(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_L g478 ( .A(n_35), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_36), .A2(n_146), .B(n_151), .C(n_170), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_37), .A2(n_151), .B(n_451), .C(n_456), .Y(n_450) );
CKINVDCx14_ASAP7_75t_R g463 ( .A(n_38), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_39), .A2(n_68), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_39), .Y(n_123) );
INVx1_ASAP7_75t_L g235 ( .A(n_41), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_42), .A2(n_177), .B(n_223), .C(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_43), .B(n_190), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g715 ( .A1(n_44), .A2(n_84), .B1(n_716), .B2(n_717), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_44), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_45), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_46), .Y(n_474) );
INVx1_ASAP7_75t_L g522 ( .A(n_47), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g238 ( .A(n_48), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_49), .B(n_141), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_50), .A2(n_151), .B1(n_232), .B2(n_234), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_51), .Y(n_181) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_52), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_53), .A2(n_223), .B(n_224), .C(n_226), .Y(n_222) );
CKINVDCx14_ASAP7_75t_R g553 ( .A(n_54), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_55), .Y(n_194) );
INVx1_ASAP7_75t_L g221 ( .A(n_56), .Y(n_221) );
AOI222xp33_ASAP7_75t_SL g121 ( .A1(n_57), .A2(n_122), .B1(n_125), .B2(n_706), .C1(n_707), .C2(n_708), .Y(n_121) );
INVx1_ASAP7_75t_L g147 ( .A(n_58), .Y(n_147) );
INVx1_ASAP7_75t_L g137 ( .A(n_59), .Y(n_137) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_60), .A2(n_102), .B1(n_113), .B2(n_719), .Y(n_101) );
INVx1_ASAP7_75t_SL g466 ( .A(n_61), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_62), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_63), .B(n_218), .Y(n_526) );
INVx1_ASAP7_75t_L g487 ( .A(n_64), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_SL g245 ( .A1(n_65), .A2(n_175), .B(n_226), .C(n_246), .Y(n_245) );
INVxp67_ASAP7_75t_L g247 ( .A(n_66), .Y(n_247) );
INVx1_ASAP7_75t_L g106 ( .A(n_67), .Y(n_106) );
INVx1_ASAP7_75t_L g124 ( .A(n_68), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_69), .A2(n_141), .B(n_552), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_70), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_71), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_72), .A2(n_141), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g185 ( .A(n_73), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_74), .A2(n_140), .B(n_473), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g449 ( .A(n_75), .Y(n_449) );
INVx1_ASAP7_75t_L g514 ( .A(n_76), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_77), .A2(n_146), .B(n_151), .C(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_78), .A2(n_141), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g517 ( .A(n_79), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_80), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g135 ( .A(n_81), .Y(n_135) );
INVx1_ASAP7_75t_L g506 ( .A(n_82), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_83), .B(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_84), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_85), .A2(n_146), .B(n_151), .C(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g108 ( .A(n_86), .B(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g438 ( .A(n_86), .Y(n_438) );
OR2x2_ASAP7_75t_L g705 ( .A(n_86), .B(n_110), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_87), .A2(n_151), .B(n_486), .C(n_490), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_88), .B(n_134), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_89), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_90), .A2(n_146), .B(n_151), .C(n_203), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_91), .Y(n_211) );
INVx1_ASAP7_75t_L g244 ( .A(n_92), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g149 ( .A(n_93), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_94), .B(n_172), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_95), .B(n_163), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_96), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_97), .B(n_106), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_98), .A2(n_141), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g525 ( .A(n_99), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_100), .Y(n_120) );
CKINVDCx6p67_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g720 ( .A(n_103), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_108), .Y(n_119) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_108), .Y(n_718) );
NOR2x2_ASAP7_75t_L g710 ( .A(n_109), .B(n_438), .Y(n_710) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g437 ( .A(n_110), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AOI22x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_121), .B1(n_711), .B2(n_713), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g712 ( .A(n_117), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_118), .A2(n_714), .B(n_718), .Y(n_713) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVx1_ASAP7_75t_L g706 ( .A(n_122), .Y(n_706) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_435), .B1(n_439), .B2(n_703), .Y(n_125) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g707 ( .A1(n_127), .A2(n_437), .B1(n_440), .B2(n_705), .Y(n_707) );
OR4x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_331), .C(n_390), .D(n_417), .Y(n_127) );
NAND3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_273), .C(n_298), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_196), .B(n_216), .C(n_249), .Y(n_129) );
AOI211xp5_ASAP7_75t_SL g421 ( .A1(n_130), .A2(n_422), .B(n_424), .C(n_427), .Y(n_421) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_165), .Y(n_130) );
INVx1_ASAP7_75t_L g296 ( .A(n_131), .Y(n_296) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OR2x2_ASAP7_75t_L g271 ( .A(n_132), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g303 ( .A(n_132), .Y(n_303) );
AND2x2_ASAP7_75t_L g358 ( .A(n_132), .B(n_327), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_132), .B(n_214), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_132), .B(n_215), .Y(n_416) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g277 ( .A(n_133), .Y(n_277) );
AND2x2_ASAP7_75t_L g320 ( .A(n_133), .B(n_183), .Y(n_320) );
AND2x2_ASAP7_75t_L g338 ( .A(n_133), .B(n_215), .Y(n_338) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_139), .B(n_162), .Y(n_133) );
INVx1_ASAP7_75t_L g195 ( .A(n_134), .Y(n_195) );
INVx2_ASAP7_75t_L g200 ( .A(n_134), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_134), .A2(n_186), .B(n_449), .C(n_450), .Y(n_448) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_134), .A2(n_551), .B(n_557), .Y(n_550) );
AND2x2_ASAP7_75t_SL g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_L g164 ( .A(n_135), .B(n_136), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_142), .B(n_146), .Y(n_186) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g455 ( .A(n_143), .Y(n_455) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
INVx1_ASAP7_75t_L g233 ( .A(n_144), .Y(n_233) );
INVx1_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx3_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_145), .Y(n_190) );
INVx4_ASAP7_75t_SL g161 ( .A(n_146), .Y(n_161) );
BUFx3_ASAP7_75t_L g456 ( .A(n_146), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_154), .C(n_161), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_150), .A2(n_161), .B(n_221), .C(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_150), .A2(n_161), .B(n_244), .C(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_150), .A2(n_161), .B(n_463), .C(n_464), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_SL g473 ( .A1(n_150), .A2(n_161), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_SL g513 ( .A1(n_150), .A2(n_161), .B(n_514), .C(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_SL g521 ( .A1(n_150), .A2(n_161), .B(n_522), .C(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_SL g552 ( .A1(n_150), .A2(n_161), .B(n_553), .C(n_554), .Y(n_552) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx3_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_152), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_155), .B(n_158), .Y(n_157) );
OAI22xp33_ASAP7_75t_L g476 ( .A1(n_155), .A2(n_172), .B1(n_477), .B2(n_478), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_155), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_155), .B(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_156), .A2(n_235), .B1(n_236), .B2(n_237), .Y(n_234) );
INVx2_ASAP7_75t_L g236 ( .A(n_156), .Y(n_236) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
OAI22xp33_ASAP7_75t_L g230 ( .A1(n_161), .A2(n_186), .B1(n_231), .B2(n_238), .Y(n_230) );
INVx1_ASAP7_75t_L g490 ( .A(n_161), .Y(n_490) );
INVx4_ASAP7_75t_L g182 ( .A(n_163), .Y(n_182) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_163), .A2(n_242), .B(n_248), .Y(n_241) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_163), .Y(n_460) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
INVx4_ASAP7_75t_L g270 ( .A(n_165), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_165), .A2(n_326), .B(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g406 ( .A(n_165), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_183), .Y(n_165) );
INVx1_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
AND2x2_ASAP7_75t_L g275 ( .A(n_166), .B(n_215), .Y(n_275) );
OR2x2_ASAP7_75t_L g304 ( .A(n_166), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g318 ( .A(n_166), .Y(n_318) );
INVx3_ASAP7_75t_L g327 ( .A(n_166), .Y(n_327) );
AND2x2_ASAP7_75t_L g337 ( .A(n_166), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g370 ( .A(n_166), .B(n_276), .Y(n_370) );
AND2x2_ASAP7_75t_L g394 ( .A(n_166), .B(n_350), .Y(n_394) );
OR2x6_ASAP7_75t_L g166 ( .A(n_167), .B(n_180), .Y(n_166) );
AOI21xp5_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B(n_178), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_176), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_172), .A2(n_258), .B(n_259), .C(n_260), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g451 ( .A1(n_172), .A2(n_452), .B(n_453), .C(n_454), .Y(n_451) );
INVx5_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_173), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_173), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_173), .B(n_556), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_176), .A2(n_189), .B(n_191), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_176), .A2(n_487), .B(n_488), .C(n_489), .Y(n_486) );
O2A1O1Ixp5_ASAP7_75t_L g505 ( .A1(n_176), .A2(n_488), .B(n_506), .C(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g192 ( .A(n_178), .Y(n_192) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_179), .A2(n_230), .B(n_239), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_179), .B(n_240), .Y(n_239) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_179), .A2(n_254), .B(n_261), .Y(n_253) );
NOR2xp33_ASAP7_75t_SL g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx3_ASAP7_75t_L g218 ( .A(n_182), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_182), .B(n_458), .Y(n_457) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_182), .A2(n_483), .B(n_491), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_182), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g215 ( .A(n_183), .Y(n_215) );
AND2x2_ASAP7_75t_L g430 ( .A(n_183), .B(n_272), .Y(n_430) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_192), .B(n_193), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_186), .A2(n_255), .B(n_256), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_186), .A2(n_484), .B(n_485), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_186), .A2(n_503), .B(n_504), .Y(n_502) );
INVx4_ASAP7_75t_L g206 ( .A(n_190), .Y(n_206) );
INVx2_ASAP7_75t_L g223 ( .A(n_190), .Y(n_223) );
INVx1_ASAP7_75t_L g471 ( .A(n_192), .Y(n_471) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_192), .A2(n_496), .B(n_497), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_195), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_195), .B(n_262), .Y(n_261) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_195), .A2(n_502), .B(n_508), .Y(n_501) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_212), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_198), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g350 ( .A(n_198), .B(n_338), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_198), .B(n_327), .Y(n_412) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g272 ( .A(n_199), .Y(n_272) );
AND2x2_ASAP7_75t_L g276 ( .A(n_199), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g317 ( .A(n_199), .B(n_318), .Y(n_317) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_210), .Y(n_199) );
INVx1_ASAP7_75t_L g480 ( .A(n_200), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_200), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_209), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_207), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_206), .B(n_466), .Y(n_465) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g226 ( .A(n_208), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_212), .B(n_313), .Y(n_335) );
INVx1_ASAP7_75t_L g374 ( .A(n_212), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_212), .B(n_301), .Y(n_418) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AND2x2_ASAP7_75t_L g281 ( .A(n_213), .B(n_276), .Y(n_281) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_215), .B(n_272), .Y(n_305) );
INVx1_ASAP7_75t_L g384 ( .A(n_215), .Y(n_384) );
AOI322xp5_ASAP7_75t_L g408 ( .A1(n_216), .A2(n_323), .A3(n_383), .B1(n_409), .B2(n_411), .C1(n_413), .C2(n_415), .Y(n_408) );
AND2x2_ASAP7_75t_SL g216 ( .A(n_217), .B(n_228), .Y(n_216) );
AND2x2_ASAP7_75t_L g263 ( .A(n_217), .B(n_241), .Y(n_263) );
INVx1_ASAP7_75t_SL g266 ( .A(n_217), .Y(n_266) );
AND2x2_ASAP7_75t_L g268 ( .A(n_217), .B(n_229), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_217), .B(n_285), .Y(n_291) );
INVx2_ASAP7_75t_L g310 ( .A(n_217), .Y(n_310) );
AND2x2_ASAP7_75t_L g323 ( .A(n_217), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g361 ( .A(n_217), .B(n_285), .Y(n_361) );
BUFx2_ASAP7_75t_L g378 ( .A(n_217), .Y(n_378) );
AND2x2_ASAP7_75t_L g392 ( .A(n_217), .B(n_252), .Y(n_392) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_227), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_228), .B(n_280), .Y(n_307) );
AND2x2_ASAP7_75t_L g434 ( .A(n_228), .B(n_310), .Y(n_434) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_241), .Y(n_228) );
OR2x2_ASAP7_75t_L g279 ( .A(n_229), .B(n_280), .Y(n_279) );
INVx3_ASAP7_75t_L g285 ( .A(n_229), .Y(n_285) );
AND2x2_ASAP7_75t_L g330 ( .A(n_229), .B(n_253), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_229), .B(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_229), .Y(n_414) );
INVx2_ASAP7_75t_L g260 ( .A(n_232), .Y(n_260) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g488 ( .A(n_236), .Y(n_488) );
AND2x2_ASAP7_75t_L g265 ( .A(n_241), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g287 ( .A(n_241), .Y(n_287) );
BUFx2_ASAP7_75t_L g293 ( .A(n_241), .Y(n_293) );
AND2x2_ASAP7_75t_L g312 ( .A(n_241), .B(n_285), .Y(n_312) );
INVx3_ASAP7_75t_L g324 ( .A(n_241), .Y(n_324) );
OR2x2_ASAP7_75t_L g334 ( .A(n_241), .B(n_285), .Y(n_334) );
AOI31xp33_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_264), .A3(n_267), .B(n_269), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_263), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_251), .B(n_286), .Y(n_297) );
OR2x2_ASAP7_75t_L g321 ( .A(n_251), .B(n_291), .Y(n_321) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_252), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g342 ( .A(n_252), .B(n_334), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_252), .B(n_324), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_252), .B(n_360), .Y(n_359) );
NAND2x1_ASAP7_75t_L g387 ( .A(n_252), .B(n_323), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_252), .B(n_378), .Y(n_388) );
AND2x2_ASAP7_75t_L g400 ( .A(n_252), .B(n_285), .Y(n_400) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g280 ( .A(n_253), .Y(n_280) );
INVx1_ASAP7_75t_L g346 ( .A(n_263), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_263), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_265), .B(n_341), .Y(n_375) );
AND2x4_ASAP7_75t_L g286 ( .A(n_266), .B(n_287), .Y(n_286) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g365 ( .A(n_271), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_271), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g313 ( .A(n_272), .B(n_303), .Y(n_313) );
AND2x2_ASAP7_75t_L g407 ( .A(n_272), .B(n_277), .Y(n_407) );
INVx1_ASAP7_75t_L g432 ( .A(n_272), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_278), .B1(n_281), .B2(n_282), .C(n_288), .Y(n_273) );
CKINVDCx14_ASAP7_75t_R g294 ( .A(n_274), .Y(n_294) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_275), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_278), .B(n_329), .Y(n_348) );
INVx3_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g397 ( .A(n_279), .B(n_293), .Y(n_397) );
AND2x2_ASAP7_75t_L g311 ( .A(n_280), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g341 ( .A(n_280), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_280), .B(n_324), .Y(n_369) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_280), .B(n_381), .C(n_412), .Y(n_411) );
AOI211xp5_ASAP7_75t_SL g344 ( .A1(n_281), .A2(n_345), .B(n_347), .C(n_355), .Y(n_344) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_283), .A2(n_334), .B1(n_335), .B2(n_336), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_284), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_284), .B(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g426 ( .A(n_286), .B(n_400), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_294), .B1(n_295), .B2(n_297), .Y(n_288) );
NOR2xp33_ASAP7_75t_SL g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_292), .B(n_341), .Y(n_372) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_295), .A2(n_387), .B1(n_418), .B2(n_425), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_306), .B1(n_308), .B2(n_313), .C(n_314), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI221xp5_ASAP7_75t_L g314 ( .A1(n_304), .A2(n_315), .B1(n_321), .B2(n_322), .C(n_325), .Y(n_314) );
INVx1_ASAP7_75t_L g357 ( .A(n_305), .Y(n_357) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_SL g329 ( .A(n_310), .Y(n_329) );
OR2x2_ASAP7_75t_L g402 ( .A(n_310), .B(n_334), .Y(n_402) );
AND2x2_ASAP7_75t_L g404 ( .A(n_310), .B(n_312), .Y(n_404) );
INVx1_ASAP7_75t_L g343 ( .A(n_313), .Y(n_343) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .Y(n_315) );
AOI21xp33_ASAP7_75t_SL g373 ( .A1(n_316), .A2(n_374), .B(n_375), .Y(n_373) );
OR2x2_ASAP7_75t_L g380 ( .A(n_316), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g354 ( .A(n_317), .B(n_338), .Y(n_354) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp33_ASAP7_75t_SL g371 ( .A(n_322), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_323), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_324), .B(n_360), .Y(n_423) );
O2A1O1Ixp33_ASAP7_75t_L g339 ( .A1(n_327), .A2(n_340), .B(n_342), .C(n_343), .Y(n_339) );
NAND2x1_ASAP7_75t_SL g364 ( .A(n_327), .B(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_328), .A2(n_377), .B1(n_379), .B2(n_382), .Y(n_376) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_330), .B(n_420), .Y(n_419) );
NAND5xp2_ASAP7_75t_L g331 ( .A(n_332), .B(n_344), .C(n_362), .D(n_376), .E(n_385), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_339), .Y(n_332) );
INVx1_ASAP7_75t_L g389 ( .A(n_335), .Y(n_389) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_337), .A2(n_356), .B1(n_396), .B2(n_398), .C(n_401), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_338), .B(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_341), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_341), .B(n_407), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_351), .B2(n_353), .Y(n_347) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_359), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AND2x2_ASAP7_75t_L g429 ( .A(n_358), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B1(n_370), .B2(n_371), .C(n_373), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g413 ( .A(n_368), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g420 ( .A(n_378), .Y(n_420) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI21xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_388), .B(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI211xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_393), .B(n_395), .C(n_408), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
A2O1A1Ixp33_ASAP7_75t_L g417 ( .A1(n_393), .A2(n_418), .B(n_419), .C(n_421), .Y(n_417) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_397), .B(n_399), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_431), .B(n_433), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
XOR2xp5_ASAP7_75t_L g714 ( .A(n_440), .B(n_715), .Y(n_714) );
OR3x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_614), .C(n_661), .Y(n_440) );
NAND3xp33_ASAP7_75t_SL g441 ( .A(n_442), .B(n_560), .C(n_585), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_500), .B1(n_527), .B2(n_530), .C(n_538), .Y(n_442) );
OAI21xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_468), .B(n_493), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_445), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_445), .B(n_543), .Y(n_658) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_459), .Y(n_445) );
AND2x2_ASAP7_75t_L g529 ( .A(n_446), .B(n_499), .Y(n_529) );
AND2x2_ASAP7_75t_L g578 ( .A(n_446), .B(n_498), .Y(n_578) );
AND2x2_ASAP7_75t_L g599 ( .A(n_446), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g604 ( .A(n_446), .B(n_571), .Y(n_604) );
OR2x2_ASAP7_75t_L g612 ( .A(n_446), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g684 ( .A(n_446), .B(n_481), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_446), .B(n_633), .Y(n_698) );
INVx3_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g544 ( .A(n_447), .B(n_459), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_447), .B(n_481), .Y(n_545) );
AND2x4_ASAP7_75t_L g566 ( .A(n_447), .B(n_499), .Y(n_566) );
AND2x2_ASAP7_75t_L g596 ( .A(n_447), .B(n_470), .Y(n_596) );
AND2x2_ASAP7_75t_L g605 ( .A(n_447), .B(n_595), .Y(n_605) );
AND2x2_ASAP7_75t_L g621 ( .A(n_447), .B(n_482), .Y(n_621) );
OR2x2_ASAP7_75t_L g630 ( .A(n_447), .B(n_613), .Y(n_630) );
AND2x2_ASAP7_75t_L g636 ( .A(n_447), .B(n_571), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_447), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g650 ( .A(n_447), .B(n_495), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_447), .B(n_540), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_447), .B(n_600), .Y(n_689) );
OR2x6_ASAP7_75t_L g447 ( .A(n_448), .B(n_457), .Y(n_447) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_455), .B(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g499 ( .A(n_459), .Y(n_499) );
AND2x2_ASAP7_75t_L g595 ( .A(n_459), .B(n_481), .Y(n_595) );
AND2x2_ASAP7_75t_L g600 ( .A(n_459), .B(n_482), .Y(n_600) );
INVx1_ASAP7_75t_L g656 ( .A(n_459), .Y(n_656) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_467), .Y(n_459) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_460), .A2(n_512), .B(n_518), .Y(n_511) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_460), .A2(n_520), .B(n_526), .Y(n_519) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g565 ( .A(n_469), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_481), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_470), .B(n_529), .Y(n_528) );
BUFx3_ASAP7_75t_L g543 ( .A(n_470), .Y(n_543) );
OR2x2_ASAP7_75t_L g613 ( .A(n_470), .B(n_481), .Y(n_613) );
OR2x2_ASAP7_75t_L g674 ( .A(n_470), .B(n_581), .Y(n_674) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_479), .Y(n_470) );
INVx1_ASAP7_75t_L g496 ( .A(n_472), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_479), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_481), .B(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g633 ( .A(n_481), .B(n_495), .Y(n_633) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g572 ( .A(n_482), .Y(n_572) );
INVx1_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_494), .A2(n_678), .B1(n_682), .B2(n_685), .C(n_686), .Y(n_677) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .Y(n_494) );
INVx1_ASAP7_75t_SL g541 ( .A(n_495), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_495), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g672 ( .A(n_495), .B(n_529), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_498), .B(n_543), .Y(n_664) );
AND2x2_ASAP7_75t_L g571 ( .A(n_499), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g575 ( .A(n_500), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_500), .B(n_581), .Y(n_611) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
AND2x2_ASAP7_75t_L g537 ( .A(n_501), .B(n_511), .Y(n_537) );
INVx4_ASAP7_75t_L g549 ( .A(n_501), .Y(n_549) );
BUFx3_ASAP7_75t_L g591 ( .A(n_501), .Y(n_591) );
AND3x2_ASAP7_75t_L g606 ( .A(n_501), .B(n_607), .C(n_608), .Y(n_606) );
AND2x2_ASAP7_75t_L g688 ( .A(n_510), .B(n_602), .Y(n_688) );
AND2x2_ASAP7_75t_L g696 ( .A(n_510), .B(n_581), .Y(n_696) );
INVx1_ASAP7_75t_SL g701 ( .A(n_510), .Y(n_701) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_519), .Y(n_510) );
INVx1_ASAP7_75t_SL g559 ( .A(n_511), .Y(n_559) );
AND2x2_ASAP7_75t_L g582 ( .A(n_511), .B(n_549), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_511), .B(n_533), .Y(n_584) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_511), .Y(n_624) );
OR2x2_ASAP7_75t_L g629 ( .A(n_511), .B(n_549), .Y(n_629) );
INVx2_ASAP7_75t_L g535 ( .A(n_519), .Y(n_535) );
AND2x2_ASAP7_75t_L g569 ( .A(n_519), .B(n_550), .Y(n_569) );
OR2x2_ASAP7_75t_L g589 ( .A(n_519), .B(n_550), .Y(n_589) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_519), .Y(n_609) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_528), .A2(n_568), .B(n_660), .Y(n_659) );
AOI322xp5_ASAP7_75t_L g695 ( .A1(n_530), .A2(n_540), .A3(n_566), .B1(n_696), .B2(n_697), .C1(n_699), .C2(n_702), .Y(n_695) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_536), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_532), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_533), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g558 ( .A(n_534), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g626 ( .A(n_535), .B(n_549), .Y(n_626) );
AND2x2_ASAP7_75t_L g693 ( .A(n_535), .B(n_550), .Y(n_693) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g634 ( .A(n_537), .B(n_588), .Y(n_634) );
AOI31xp33_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_542), .A3(n_545), .B(n_546), .Y(n_538) );
AND2x2_ASAP7_75t_L g593 ( .A(n_540), .B(n_571), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_540), .B(n_563), .Y(n_675) );
AND2x2_ASAP7_75t_L g694 ( .A(n_540), .B(n_599), .Y(n_694) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_543), .B(n_571), .Y(n_583) );
NAND2x1p5_ASAP7_75t_L g617 ( .A(n_543), .B(n_600), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_543), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_543), .B(n_684), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_544), .B(n_600), .Y(n_632) );
INVx1_ASAP7_75t_L g676 ( .A(n_544), .Y(n_676) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_558), .Y(n_547) );
INVxp67_ASAP7_75t_L g628 ( .A(n_548), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_549), .B(n_559), .Y(n_564) );
INVx1_ASAP7_75t_L g670 ( .A(n_549), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_549), .B(n_647), .Y(n_681) );
BUFx3_ASAP7_75t_L g581 ( .A(n_550), .Y(n_581) );
AND2x2_ASAP7_75t_L g607 ( .A(n_550), .B(n_559), .Y(n_607) );
INVx2_ASAP7_75t_L g647 ( .A(n_550), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_558), .B(n_680), .Y(n_679) );
AOI211xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_565), .B(n_567), .C(n_576), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_562), .A2(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_563), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_563), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g643 ( .A(n_564), .B(n_589), .Y(n_643) );
INVx3_ASAP7_75t_L g574 ( .A(n_566), .Y(n_574) );
OAI22xp5_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_570), .B1(n_573), .B2(n_575), .Y(n_567) );
OAI21xp5_ASAP7_75t_SL g592 ( .A1(n_569), .A2(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g618 ( .A(n_569), .B(n_582), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_569), .B(n_670), .Y(n_669) );
INVxp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g573 ( .A(n_572), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g642 ( .A(n_572), .Y(n_642) );
OAI21xp5_ASAP7_75t_SL g586 ( .A1(n_573), .A2(n_587), .B(n_592), .Y(n_586) );
OAI22xp33_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_579), .B1(n_583), .B2(n_584), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_578), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g602 ( .A(n_581), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_581), .B(n_624), .Y(n_623) );
NOR3xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_597), .C(n_610), .Y(n_585) );
OAI22xp5_ASAP7_75t_SL g652 ( .A1(n_587), .A2(n_653), .B1(n_657), .B2(n_658), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g657 ( .A(n_589), .B(n_590), .Y(n_657) );
AND2x2_ASAP7_75t_L g665 ( .A(n_590), .B(n_646), .Y(n_665) );
CKINVDCx16_ASAP7_75t_R g590 ( .A(n_591), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_SL g673 ( .A1(n_591), .A2(n_674), .B(n_675), .C(n_676), .Y(n_673) );
OR2x2_ASAP7_75t_L g700 ( .A(n_591), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
OAI21xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_601), .B(n_603), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_599), .A2(n_636), .B(n_637), .C(n_640), .Y(n_635) );
OAI21xp33_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_605), .B(n_606), .Y(n_603) );
AND2x2_ASAP7_75t_L g668 ( .A(n_607), .B(n_626), .Y(n_668) );
INVxp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g646 ( .A(n_609), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g651 ( .A(n_611), .Y(n_651) );
NAND3xp33_ASAP7_75t_SL g614 ( .A(n_615), .B(n_635), .C(n_648), .Y(n_614) );
AOI211xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B(n_619), .C(n_627), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g685 ( .A(n_622), .Y(n_685) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g645 ( .A(n_624), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_624), .B(n_693), .Y(n_692) );
INVxp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B(n_630), .C(n_631), .Y(n_627) );
INVx2_ASAP7_75t_SL g639 ( .A(n_629), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_630), .A2(n_641), .B1(n_643), .B2(n_644), .Y(n_640) );
OAI21xp33_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_633), .B(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
AOI211xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B(n_652), .C(n_659), .Y(n_648) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVxp33_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g702 ( .A(n_656), .Y(n_702) );
NAND4xp25_ASAP7_75t_L g661 ( .A(n_662), .B(n_677), .C(n_690), .D(n_695), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_665), .B(n_666), .C(n_673), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B(n_671), .Y(n_666) );
AOI21xp33_ASAP7_75t_L g686 ( .A1(n_667), .A2(n_687), .B(n_689), .Y(n_686) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_674), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .Y(n_690) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
endmodule