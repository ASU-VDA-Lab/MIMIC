module fake_jpeg_11574_n_575 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_575);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_575;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_14),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_55),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_57),
.Y(n_148)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_70),
.Y(n_110)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_77),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_30),
.B(n_11),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_80),
.Y(n_121)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_30),
.B(n_11),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_90),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx11_ASAP7_75t_SL g174 ( 
.A(n_87),
.Y(n_174)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx16f_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_34),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_95),
.B(n_97),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_25),
.B(n_10),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_99),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g122 ( 
.A(n_98),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_103),
.Y(n_160)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_54),
.Y(n_135)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_104),
.Y(n_124)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_25),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g131 ( 
.A(n_106),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_38),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_119),
.B(n_127),
.Y(n_203)
);

INVx2_ASAP7_75t_R g120 ( 
.A(n_87),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_120),
.B(n_135),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_69),
.A2(n_53),
.B1(n_51),
.B2(n_32),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_126),
.A2(n_157),
.B1(n_158),
.B2(n_109),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_77),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_23),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_21),
.B(n_43),
.C(n_54),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_58),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_42),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_144),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_89),
.B(n_42),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_50),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_155),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_53),
.C(n_43),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_151),
.B(n_171),
.Y(n_224)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_74),
.B(n_35),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_88),
.A2(n_38),
.B1(n_53),
.B2(n_95),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_82),
.A2(n_20),
.B1(n_23),
.B2(n_38),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_67),
.B(n_50),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_166),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_79),
.B(n_35),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_84),
.B(n_27),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_173),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_98),
.B(n_27),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_56),
.B1(n_60),
.B2(n_59),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_175),
.A2(n_188),
.B1(n_86),
.B2(n_81),
.Y(n_265)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_177),
.A2(n_170),
.B1(n_168),
.B2(n_163),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_179),
.B(n_186),
.Y(n_245)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_181),
.Y(n_260)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_184),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_118),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_83),
.B1(n_107),
.B2(n_99),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_133),
.Y(n_189)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_136),
.B(n_20),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_193),
.B(n_196),
.Y(n_248)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_195),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_121),
.B(n_44),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_124),
.B(n_44),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_198),
.B(n_202),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_131),
.Y(n_199)
);

INVx11_ASAP7_75t_L g289 ( 
.A(n_199),
.Y(n_289)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_46),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_204),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_117),
.B(n_46),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g280 ( 
.A1(n_205),
.A2(n_234),
.B(n_235),
.Y(n_280)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_130),
.Y(n_206)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_206),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_110),
.B(n_33),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_208),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_138),
.B(n_33),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_158),
.A2(n_61),
.B1(n_64),
.B2(n_68),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_209),
.A2(n_214),
.B1(n_76),
.B2(n_91),
.Y(n_255)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_210),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_152),
.B(n_20),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_213),
.Y(n_250)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_147),
.Y(n_212)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_212),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_146),
.Y(n_216)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_217),
.Y(n_291)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_220),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_114),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_221),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_143),
.B(n_97),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_223),
.Y(n_274)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_114),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_132),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_225),
.B(n_226),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_125),
.B(n_94),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_153),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_227),
.Y(n_259)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_228),
.B(n_231),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_111),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_230),
.B1(n_233),
.B2(n_237),
.Y(n_254)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_132),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_125),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_156),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_232),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_128),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_120),
.B(n_156),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_137),
.B(n_0),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_123),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_236),
.Y(n_269)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_128),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_151),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_241),
.B(n_244),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_142),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_246),
.B(n_4),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_193),
.B(n_192),
.C(n_177),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_213),
.C(n_217),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_255),
.A2(n_264),
.B1(n_278),
.B2(n_285),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_234),
.A2(n_170),
.B(n_168),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_258),
.A2(n_178),
.B(n_189),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_192),
.A2(n_116),
.B1(n_167),
.B2(n_163),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_265),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_200),
.B(n_162),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_266),
.B(n_273),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_181),
.A2(n_116),
.B1(n_167),
.B2(n_162),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_270),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_194),
.B(n_142),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_175),
.A2(n_139),
.B1(n_145),
.B2(n_141),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_275),
.A2(n_237),
.B1(n_190),
.B2(n_210),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_187),
.B(n_113),
.CI(n_154),
.CON(n_276),
.SN(n_276)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_290),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_182),
.B(n_139),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_277),
.B(n_8),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_209),
.A2(n_129),
.B1(n_145),
.B2(n_141),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_230),
.A2(n_129),
.B1(n_113),
.B2(n_174),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_188),
.A2(n_174),
.B1(n_37),
.B2(n_22),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_195),
.A2(n_123),
.B1(n_37),
.B2(n_22),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_286),
.A2(n_178),
.B1(n_199),
.B2(n_212),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_203),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_176),
.A2(n_37),
.B1(n_22),
.B2(n_123),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_293),
.A2(n_185),
.B1(n_37),
.B2(n_22),
.Y(n_326)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_305),
.C(n_311),
.Y(n_344)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_296),
.Y(n_371)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_299),
.A2(n_262),
.B1(n_240),
.B2(n_261),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_199),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_301),
.B(n_302),
.Y(n_349)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_241),
.B(n_227),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_253),
.Y(n_306)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_307),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_284),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_315),
.Y(n_356)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_284),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_310),
.B(n_327),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_244),
.B(n_215),
.C(n_221),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_312),
.Y(n_368)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_272),
.Y(n_314)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_314),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_245),
.B(n_178),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_316),
.B(n_317),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_242),
.B(n_233),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_318),
.B(n_321),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_251),
.B(n_229),
.C(n_204),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_319),
.B(n_336),
.C(n_343),
.Y(n_376)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_243),
.Y(n_321)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_240),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_322),
.B(n_325),
.Y(n_384)
);

INVx13_ASAP7_75t_L g323 ( 
.A(n_281),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_323),
.Y(n_350)
);

AND2x6_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_0),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_328),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_268),
.B(n_197),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_326),
.A2(n_259),
.B1(n_247),
.B2(n_291),
.Y(n_360)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_243),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_248),
.B(n_0),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_275),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_329),
.A2(n_331),
.B1(n_340),
.B2(n_341),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_255),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_330),
.A2(n_263),
.B1(n_239),
.B2(n_262),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_281),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_266),
.B(n_1),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_333),
.B(n_335),
.Y(n_370)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_252),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_337),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_284),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_273),
.B(n_3),
.C(n_4),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_293),
.Y(n_351)
);

INVx13_ASAP7_75t_L g340 ( 
.A(n_249),
.Y(n_340)
);

INVx3_ASAP7_75t_SL g341 ( 
.A(n_238),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_288),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_292),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_277),
.B(n_5),
.C(n_6),
.Y(n_343)
);

FAx1_ASAP7_75t_SL g345 ( 
.A(n_313),
.B(n_280),
.CI(n_276),
.CON(n_345),
.SN(n_345)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_345),
.B(n_300),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_346),
.B(n_367),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_305),
.B(n_250),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_347),
.B(n_363),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_351),
.B(n_360),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_320),
.A2(n_303),
.B1(n_295),
.B2(n_310),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_352),
.A2(n_386),
.B(n_314),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_313),
.A2(n_274),
.B1(n_282),
.B2(n_254),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_353),
.A2(n_372),
.B1(n_377),
.B2(n_382),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_339),
.A2(n_239),
.B1(n_263),
.B2(n_261),
.Y(n_358)
);

OA22x2_ASAP7_75t_L g405 ( 
.A1(n_358),
.A2(n_302),
.B1(n_294),
.B2(n_334),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_332),
.B(n_319),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_332),
.B(n_271),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_365),
.B(n_381),
.C(n_385),
.Y(n_415)
);

OAI32xp33_ASAP7_75t_L g367 ( 
.A1(n_298),
.A2(n_257),
.A3(n_247),
.B1(n_267),
.B2(n_291),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_337),
.B(n_292),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_369),
.B(n_326),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_339),
.A2(n_258),
.B1(n_257),
.B2(n_256),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_338),
.A2(n_256),
.B1(n_288),
.B2(n_267),
.Y(n_377)
);

XOR2x2_ASAP7_75t_L g378 ( 
.A(n_311),
.B(n_324),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_343),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_312),
.A2(n_252),
.B(n_283),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_380),
.A2(n_296),
.B(n_297),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_283),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_303),
.A2(n_238),
.B1(n_6),
.B2(n_7),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_304),
.B(n_5),
.C(n_6),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_306),
.B(n_5),
.Y(n_386)
);

INVx13_ASAP7_75t_L g388 ( 
.A(n_371),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_388),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_389),
.B(n_409),
.Y(n_445)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_355),
.Y(n_391)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_391),
.Y(n_435)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_392),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_370),
.B(n_309),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_393),
.B(n_414),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_349),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_395),
.B(n_398),
.Y(n_433)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_364),
.Y(n_396)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_396),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_354),
.A2(n_320),
.B1(n_341),
.B2(n_300),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_397),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_321),
.Y(n_400)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_400),
.Y(n_451)
);

NOR3xp33_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_357),
.C(n_345),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_327),
.Y(n_402)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_402),
.Y(n_455)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_375),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_404),
.B(n_410),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_411),
.Y(n_426)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_356),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_417),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_368),
.A2(n_323),
.B(n_340),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_407),
.A2(n_419),
.B(n_380),
.Y(n_429)
);

CKINVDCx12_ASAP7_75t_R g408 ( 
.A(n_344),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_408),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_383),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_365),
.B(n_322),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_348),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_418),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_330),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_416),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_342),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_315),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_347),
.B(n_318),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_348),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_344),
.B(n_7),
.C(n_8),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_423),
.C(n_424),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_363),
.B(n_8),
.C(n_376),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_376),
.B(n_381),
.C(n_369),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_378),
.B(n_352),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_353),
.C(n_374),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_350),
.Y(n_430)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_447),
.C(n_456),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_403),
.A2(n_368),
.B(n_354),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_437),
.B(n_438),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_361),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_440),
.B(n_442),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_361),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_400),
.B(n_402),
.Y(n_444)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_444),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_374),
.Y(n_446)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_446),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_422),
.B(n_424),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_411),
.B(n_374),
.Y(n_449)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_396),
.B(n_358),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_452),
.B(n_405),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_386),
.Y(n_453)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_453),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_388),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_454),
.B(n_418),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_345),
.C(n_372),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_351),
.C(n_346),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_415),
.C(n_409),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_432),
.B(n_420),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_467),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_461),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_444),
.B(n_390),
.Y(n_462)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_462),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_439),
.A2(n_413),
.B1(n_390),
.B2(n_394),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_464),
.A2(n_477),
.B1(n_457),
.B2(n_456),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_465),
.B(n_470),
.C(n_445),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_432),
.B(n_443),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_439),
.A2(n_399),
.B1(n_403),
.B2(n_394),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_468),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_447),
.B(n_415),
.C(n_389),
.Y(n_470)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_472),
.Y(n_497)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_442),
.Y(n_473)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_473),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_426),
.A2(n_399),
.B1(n_451),
.B2(n_455),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_474),
.Y(n_498)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_430),
.Y(n_475)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_475),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_440),
.B(n_455),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_476),
.B(n_480),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_426),
.A2(n_451),
.B1(n_458),
.B2(n_434),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_443),
.B(n_398),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_452),
.B(n_419),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_481),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_448),
.A2(n_387),
.B1(n_425),
.B2(n_405),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_483),
.B(n_486),
.Y(n_495)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_435),
.Y(n_484)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_484),
.Y(n_500)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_435),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_477),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_489),
.B(n_504),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_445),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_490),
.B(n_505),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_485),
.A2(n_437),
.B(n_429),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_491),
.A2(n_502),
.B(n_407),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_494),
.A2(n_474),
.B1(n_471),
.B2(n_468),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_427),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_499),
.B(n_501),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_485),
.A2(n_481),
.B(n_466),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_470),
.B(n_427),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_463),
.B(n_449),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_466),
.B(n_428),
.C(n_446),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_506),
.B(n_507),
.C(n_501),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_469),
.B(n_428),
.C(n_433),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_511),
.B(n_517),
.Y(n_540)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_508),
.Y(n_512)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_512),
.Y(n_536)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_503),
.Y(n_513)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_513),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_475),
.Y(n_514)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_514),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_493),
.A2(n_478),
.B(n_476),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_515),
.Y(n_533)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_500),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_516),
.B(n_522),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_496),
.A2(n_464),
.B1(n_462),
.B2(n_460),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_487),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_519),
.B(n_509),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_520),
.A2(n_527),
.B1(n_492),
.B2(n_495),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_491),
.Y(n_530)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_488),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_505),
.B(n_489),
.C(n_506),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_523),
.B(n_524),
.C(n_511),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_504),
.B(n_469),
.C(n_471),
.Y(n_524)
);

FAx1_ASAP7_75t_SL g525 ( 
.A(n_502),
.B(n_460),
.CI(n_453),
.CON(n_525),
.SN(n_525)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_525),
.B(n_528),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_498),
.A2(n_473),
.B1(n_461),
.B2(n_486),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_498),
.A2(n_482),
.B1(n_484),
.B2(n_454),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_514),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_529),
.B(n_531),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_530),
.B(n_521),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_534),
.B(n_535),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_490),
.C(n_507),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_538),
.A2(n_541),
.B(n_542),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_510),
.B(n_497),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_526),
.B(n_494),
.C(n_450),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_526),
.B(n_441),
.C(n_405),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_543),
.B(n_528),
.C(n_522),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_540),
.B(n_515),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_545),
.A2(n_539),
.B(n_530),
.Y(n_556)
);

OA21x2_ASAP7_75t_L g546 ( 
.A1(n_533),
.A2(n_517),
.B(n_520),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_546),
.A2(n_555),
.B1(n_544),
.B2(n_545),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_518),
.C(n_524),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_547),
.B(n_548),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_540),
.B(n_518),
.C(n_527),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_549),
.B(n_552),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_542),
.B(n_525),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_554),
.B(n_535),
.C(n_543),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_533),
.A2(n_431),
.B1(n_525),
.B2(n_441),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_556),
.A2(n_551),
.B(n_546),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_558),
.B(n_559),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_550),
.B(n_553),
.C(n_547),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_560),
.B(n_562),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_548),
.B(n_532),
.C(n_536),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_557),
.B(n_554),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_563),
.A2(n_565),
.B(n_561),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_564),
.Y(n_567)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_567),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_566),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_569),
.B(n_561),
.C(n_537),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_570),
.C(n_431),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_572),
.B(n_436),
.C(n_385),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_573),
.B(n_436),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_574),
.A2(n_386),
.B(n_382),
.Y(n_575)
);


endmodule