module fake_jpeg_11946_n_286 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_7),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_0),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_51),
.C(n_36),
.Y(n_88)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_13),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_24),
.B(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_11),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_24),
.B(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_17),
.B1(n_33),
.B2(n_19),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_58),
.A2(n_70),
.B1(n_93),
.B2(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_68),
.Y(n_113)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_64),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_69),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_28),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_35),
.B1(n_34),
.B2(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_30),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_79),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_17),
.B1(n_33),
.B2(n_25),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_23),
.B1(n_27),
.B2(n_47),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_16),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_18),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_17),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_80),
.A2(n_101),
.B(n_1),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_18),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_82),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_18),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_95),
.C(n_21),
.Y(n_104)
);

OA22x2_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_56),
.B1(n_21),
.B2(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_47),
.A2(n_35),
.B1(n_34),
.B2(n_19),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_25),
.C(n_23),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_42),
.B(n_18),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_33),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_58),
.A2(n_55),
.B1(n_23),
.B2(n_25),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_107),
.B1(n_118),
.B2(n_120),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_104),
.B(n_66),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_34),
.B1(n_36),
.B2(n_27),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_45),
.B1(n_25),
.B2(n_23),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_109),
.A2(n_124),
.B1(n_89),
.B2(n_84),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_42),
.C(n_32),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_98),
.C(n_89),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_80),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_66),
.B1(n_86),
.B2(n_92),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_4),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_67),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_133),
.B(n_134),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_63),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_57),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_140),
.B(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_57),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_77),
.A3(n_94),
.B1(n_101),
.B2(n_85),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_149),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_145),
.A2(n_128),
.B(n_5),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_95),
.B1(n_61),
.B2(n_91),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_164),
.B1(n_107),
.B2(n_84),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_147),
.A2(n_156),
.B1(n_132),
.B2(n_115),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_87),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_150),
.B(n_157),
.C(n_158),
.D(n_161),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_87),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_103),
.A2(n_61),
.B1(n_91),
.B2(n_96),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_59),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_59),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_166),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_117),
.B(n_59),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_100),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_110),
.B(n_9),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_163),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_171),
.B(n_183),
.Y(n_202)
);

HAxp5_ASAP7_75t_SL g172 ( 
.A(n_149),
.B(n_102),
.CON(n_172),
.SN(n_172)
);

NOR2x1_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_181),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

OAI22x1_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_121),
.B1(n_83),
.B2(n_62),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_186),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_127),
.B(n_118),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_152),
.B(n_155),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_196),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_SL g181 ( 
.A1(n_138),
.A2(n_130),
.B(n_122),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_146),
.A2(n_115),
.B1(n_106),
.B2(n_132),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_192),
.B1(n_136),
.B2(n_4),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_150),
.B(n_130),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_193),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_148),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_191),
.B(n_194),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_139),
.A2(n_157),
.B1(n_156),
.B2(n_165),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_162),
.B(n_98),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_119),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_145),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_141),
.C(n_159),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_198),
.C(n_168),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_145),
.C(n_147),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_191),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_200),
.B(n_204),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_180),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_201),
.B(n_212),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_144),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_213),
.B(n_205),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_155),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_211),
.Y(n_222)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_119),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_189),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_136),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_215),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_167),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_217),
.A2(n_171),
.B1(n_174),
.B2(n_186),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g218 ( 
.A(n_195),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_170),
.C(n_190),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_221),
.B(n_202),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_169),
.B(n_177),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_179),
.B1(n_185),
.B2(n_5),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_192),
.B1(n_187),
.B2(n_176),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_236),
.B1(n_210),
.B2(n_173),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_169),
.B(n_188),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

AOI221xp5_ASAP7_75t_L g230 ( 
.A1(n_199),
.A2(n_196),
.B1(n_188),
.B2(n_190),
.C(n_176),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_231),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_235),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_168),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_183),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_238),
.C(n_211),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_241),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_228),
.A2(n_203),
.B1(n_205),
.B2(n_198),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_229),
.A2(n_197),
.B1(n_210),
.B2(n_204),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_242),
.A2(n_251),
.B1(n_225),
.B2(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_207),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_SL g255 ( 
.A(n_248),
.B(n_250),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_223),
.B(n_173),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_258),
.B1(n_240),
.B2(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_251),
.Y(n_257)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_257),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_236),
.B1(n_232),
.B2(n_234),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_244),
.A2(n_231),
.B(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_227),
.B(n_238),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_261),
.B(n_247),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_233),
.B(n_220),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_255),
.B(n_248),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_268),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_241),
.C(n_249),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_254),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_246),
.B1(n_221),
.B2(n_185),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_222),
.C(n_223),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_269),
.B(n_237),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_270),
.B(n_272),
.Y(n_276)
);

NAND4xp25_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_256),
.C(n_259),
.D(n_258),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_266),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_250),
.Y(n_272)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_279),
.B(n_274),
.Y(n_280)
);

AOI21x1_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_262),
.B(n_269),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_280),
.A2(n_279),
.B(n_276),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_270),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_272),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_283),
.C(n_246),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_246),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_179),
.Y(n_286)
);


endmodule