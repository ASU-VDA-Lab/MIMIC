module fake_netlist_1_12569_n_728 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_728);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_728;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g103 ( .A(n_47), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_82), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_4), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_74), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_7), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_101), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_87), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_60), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_34), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_28), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_83), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_78), .Y(n_115) );
BUFx5_ASAP7_75t_L g116 ( .A(n_13), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_57), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_58), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_15), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_85), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_97), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_14), .Y(n_122) );
INVxp33_ASAP7_75t_L g123 ( .A(n_91), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_54), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_86), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_53), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_66), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_31), .Y(n_128) );
INVx1_ASAP7_75t_SL g129 ( .A(n_40), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_29), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_63), .Y(n_131) );
BUFx8_ASAP7_75t_SL g132 ( .A(n_46), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_33), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_80), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_9), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_36), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_55), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_41), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_72), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_4), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_51), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_92), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_70), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_115), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_123), .B(n_0), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_116), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_116), .Y(n_148) );
OAI22xp5_ASAP7_75t_SL g149 ( .A1(n_140), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_149) );
BUFx3_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_116), .Y(n_153) );
AND2x2_ASAP7_75t_SL g154 ( .A(n_103), .B(n_20), .Y(n_154) );
CKINVDCx11_ASAP7_75t_R g155 ( .A(n_140), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_115), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_107), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_123), .B(n_1), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_107), .B(n_2), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_115), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_122), .B(n_3), .Y(n_161) );
NOR2x1_ASAP7_75t_L g162 ( .A(n_112), .B(n_3), .Y(n_162) );
BUFx8_ASAP7_75t_SL g163 ( .A(n_155), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_154), .B(n_118), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_159), .A2(n_109), .B1(n_110), .B2(n_121), .Y(n_165) );
INVx2_ASAP7_75t_SL g166 ( .A(n_150), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_144), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_159), .B(n_122), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_150), .B(n_106), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_154), .B(n_120), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_157), .B(n_113), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_144), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_146), .B(n_116), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_158), .B(n_105), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_144), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_159), .B(n_108), .Y(n_183) );
AND2x6_ASAP7_75t_L g184 ( .A(n_159), .B(n_139), .Y(n_184) );
INVx5_ASAP7_75t_L g185 ( .A(n_144), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_147), .B(n_103), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_147), .B(n_126), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_154), .B(n_127), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_161), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_161), .Y(n_190) );
OR2x2_ASAP7_75t_L g191 ( .A(n_165), .B(n_171), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_166), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_175), .B(n_161), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_168), .Y(n_194) );
NOR2x1_ASAP7_75t_L g195 ( .A(n_177), .B(n_161), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_164), .A2(n_153), .B(n_151), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_168), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_168), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_175), .B(n_162), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_177), .B(n_162), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_183), .B(n_114), .Y(n_201) );
OAI22xp5_ASAP7_75t_SL g202 ( .A1(n_165), .A2(n_149), .B1(n_109), .B2(n_110), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_189), .B(n_134), .Y(n_203) );
INVx2_ASAP7_75t_SL g204 ( .A(n_168), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_183), .B(n_151), .Y(n_205) );
NOR2xp67_ASAP7_75t_L g206 ( .A(n_189), .B(n_153), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g207 ( .A(n_189), .B(n_135), .Y(n_207) );
AO22x1_ASAP7_75t_L g208 ( .A1(n_184), .A2(n_132), .B1(n_138), .B2(n_121), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_189), .B(n_136), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_184), .A2(n_152), .B1(n_128), .B2(n_131), .Y(n_210) );
AO221x1_ASAP7_75t_L g211 ( .A1(n_163), .A2(n_149), .B1(n_132), .B2(n_138), .C(n_124), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_190), .B(n_141), .Y(n_212) );
OR2x6_ASAP7_75t_L g213 ( .A(n_190), .B(n_117), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_170), .A2(n_111), .B(n_125), .Y(n_214) );
NAND2x1p5_ASAP7_75t_L g215 ( .A(n_190), .B(n_119), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_190), .B(n_104), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_188), .B(n_129), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_169), .B(n_130), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_186), .A2(n_133), .B1(n_142), .B2(n_143), .Y(n_219) );
NOR3xp33_ASAP7_75t_L g220 ( .A(n_187), .B(n_111), .C(n_125), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_184), .B(n_137), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_184), .B(n_137), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_184), .A2(n_124), .B1(n_115), .B2(n_160), .Y(n_223) );
INVxp67_ASAP7_75t_L g224 ( .A(n_186), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_166), .B(n_124), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_184), .Y(n_226) );
AOI22xp5_ASAP7_75t_SL g227 ( .A1(n_184), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_184), .B(n_124), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_224), .B(n_172), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_226), .B(n_172), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_196), .A2(n_176), .B(n_178), .Y(n_231) );
CKINVDCx6p67_ASAP7_75t_R g232 ( .A(n_213), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_200), .B(n_176), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_200), .B(n_178), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_194), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_201), .A2(n_181), .B(n_180), .C(n_156), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_204), .Y(n_237) );
OR2x6_ASAP7_75t_L g238 ( .A(n_208), .B(n_180), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_201), .B(n_181), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_193), .A2(n_173), .B(n_182), .Y(n_240) );
INVx4_ASAP7_75t_L g241 ( .A(n_213), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_205), .A2(n_173), .B(n_182), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_199), .A2(n_206), .B(n_216), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_191), .B(n_5), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_195), .B(n_6), .Y(n_245) );
BUFx4f_ASAP7_75t_L g246 ( .A(n_215), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_213), .A2(n_160), .B1(n_156), .B2(n_185), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_197), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_212), .A2(n_173), .B(n_182), .Y(n_249) );
O2A1O1Ixp5_ASAP7_75t_L g250 ( .A1(n_203), .A2(n_179), .B(n_174), .C(n_185), .Y(n_250) );
OR2x6_ASAP7_75t_L g251 ( .A(n_202), .B(n_156), .Y(n_251) );
AOI21x1_ASAP7_75t_L g252 ( .A1(n_221), .A2(n_179), .B(n_174), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_210), .B(n_185), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_215), .B(n_8), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_207), .B(n_9), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_207), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_209), .A2(n_179), .B(n_174), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_227), .Y(n_258) );
NOR2xp67_ASAP7_75t_L g259 ( .A(n_214), .B(n_10), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_211), .B(n_10), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_244), .A2(n_220), .B(n_219), .C(n_218), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_232), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_258), .B(n_217), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_229), .B(n_198), .Y(n_264) );
INVx2_ASAP7_75t_SL g265 ( .A(n_246), .Y(n_265) );
AO22x1_ASAP7_75t_L g266 ( .A1(n_258), .A2(n_228), .B1(n_218), .B2(n_222), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_248), .Y(n_267) );
NOR2x1_ASAP7_75t_SL g268 ( .A(n_241), .B(n_192), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_246), .B(n_210), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_238), .Y(n_270) );
AND2x6_ASAP7_75t_L g271 ( .A(n_256), .B(n_228), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_241), .B(n_225), .Y(n_272) );
INVxp67_ASAP7_75t_L g273 ( .A(n_244), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_243), .A2(n_223), .B(n_160), .C(n_156), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_239), .A2(n_223), .B1(n_160), .B2(n_156), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_241), .B(n_11), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_251), .A2(n_160), .B1(n_156), .B2(n_185), .Y(n_277) );
NAND3x1_ASAP7_75t_L g278 ( .A(n_260), .B(n_11), .C(n_12), .Y(n_278) );
AO31x2_ASAP7_75t_L g279 ( .A1(n_236), .A2(n_160), .A3(n_167), .B(n_14), .Y(n_279) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_252), .A2(n_59), .B(n_94), .Y(n_280) );
AO31x2_ASAP7_75t_L g281 ( .A1(n_236), .A2(n_167), .A3(n_13), .B(n_15), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_240), .A2(n_167), .B(n_185), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_251), .B(n_12), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_267), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_273), .B(n_251), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_279), .Y(n_286) );
BUFx12f_ASAP7_75t_L g287 ( .A(n_262), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_264), .B(n_256), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_270), .A2(n_238), .B1(n_256), .B2(n_255), .Y(n_289) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_280), .A2(n_259), .B(n_231), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_282), .A2(n_249), .B(n_257), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_279), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_281), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_261), .A2(n_242), .B(n_230), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_283), .A2(n_254), .B(n_245), .C(n_233), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_279), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_281), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_274), .A2(n_230), .B(n_250), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_281), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_268), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_265), .B(n_256), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_276), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_271), .Y(n_303) );
AOI21x1_ASAP7_75t_L g304 ( .A1(n_266), .A2(n_247), .B(n_253), .Y(n_304) );
AO31x2_ASAP7_75t_L g305 ( .A1(n_275), .A2(n_248), .A3(n_234), .B(n_237), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_300), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_293), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_302), .B(n_271), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_293), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_302), .B(n_238), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_286), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_291), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_286), .Y(n_315) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_292), .A2(n_277), .B(n_253), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_287), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_292), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_305), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_296), .A2(n_277), .B(n_278), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_296), .Y(n_321) );
AOI21x1_ASAP7_75t_L g322 ( .A1(n_297), .A2(n_269), .B(n_272), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_300), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_288), .B(n_271), .Y(n_324) );
OA21x2_ASAP7_75t_L g325 ( .A1(n_297), .A2(n_235), .B(n_272), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_305), .Y(n_326) );
OR2x6_ASAP7_75t_L g327 ( .A(n_303), .B(n_271), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_299), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_303), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_285), .B(n_263), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_299), .B(n_61), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_288), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_291), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_290), .A2(n_167), .B(n_62), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_313), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_309), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_307), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_309), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_325), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_313), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_325), .Y(n_342) );
INVx4_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_311), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_332), .B(n_289), .Y(n_345) );
INVx5_ASAP7_75t_L g346 ( .A(n_331), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_307), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_332), .B(n_289), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_306), .B(n_305), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_313), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_315), .B(n_305), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_306), .B(n_295), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_308), .B(n_305), .Y(n_353) );
INVx5_ASAP7_75t_L g354 ( .A(n_331), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_307), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_313), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_315), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_318), .B(n_321), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_328), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_331), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_323), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_328), .Y(n_362) );
INVx4_ASAP7_75t_L g363 ( .A(n_323), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_308), .B(n_294), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_326), .Y(n_365) );
INVx5_ASAP7_75t_L g366 ( .A(n_331), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_318), .B(n_290), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_321), .B(n_290), .Y(n_368) );
NOR2x1p5_ASAP7_75t_L g369 ( .A(n_323), .B(n_287), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_328), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_328), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_325), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_312), .B(n_298), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_331), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_333), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_333), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_326), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_325), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_319), .B(n_290), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_319), .B(n_304), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_319), .B(n_304), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_331), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_323), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_346), .B(n_329), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_346), .B(n_329), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_336), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_343), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_336), .B(n_312), .Y(n_388) );
AND2x4_ASAP7_75t_SL g389 ( .A(n_343), .B(n_324), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_373), .B(n_325), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_358), .B(n_325), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_358), .B(n_316), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_335), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_358), .B(n_316), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_373), .B(n_330), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_338), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_351), .B(n_316), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_351), .B(n_316), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_369), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_351), .B(n_338), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_377), .B(n_330), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_346), .B(n_329), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_341), .B(n_316), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_335), .Y(n_404) );
INVx3_ASAP7_75t_L g405 ( .A(n_343), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_377), .B(n_330), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_349), .B(n_310), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_341), .B(n_344), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_345), .B(n_317), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_344), .B(n_333), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_357), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_352), .B(n_312), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_335), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_349), .B(n_310), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_357), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_340), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_340), .Y(n_417) );
NOR2x1_ASAP7_75t_L g418 ( .A(n_369), .B(n_327), .Y(n_418) );
OR2x6_ASAP7_75t_L g419 ( .A(n_343), .B(n_320), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_340), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_379), .B(n_333), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_347), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_352), .B(n_324), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_343), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_379), .B(n_324), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_379), .B(n_322), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_345), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_380), .B(n_322), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_380), .B(n_322), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_350), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_349), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_371), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_380), .B(n_314), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_337), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_347), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_346), .B(n_329), .Y(n_436) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_339), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_345), .B(n_320), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_381), .B(n_314), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_371), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_350), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_381), .B(n_314), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_350), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_348), .B(n_320), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_381), .B(n_314), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_347), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_348), .B(n_314), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_356), .B(n_314), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_339), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_348), .B(n_317), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_356), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_363), .B(n_16), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_353), .B(n_314), .Y(n_453) );
NAND2x1p5_ASAP7_75t_L g454 ( .A(n_346), .B(n_334), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_356), .B(n_327), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_359), .B(n_314), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_359), .B(n_327), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_408), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_409), .B(n_363), .Y(n_459) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_399), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_395), .B(n_378), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_400), .B(n_342), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_400), .B(n_342), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_425), .B(n_361), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_393), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_395), .B(n_378), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_401), .B(n_372), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_408), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_389), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_387), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g471 ( .A(n_418), .B(n_346), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_397), .B(n_368), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_386), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_397), .B(n_368), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_398), .B(n_368), .Y(n_475) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_452), .B(n_363), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_386), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_396), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_398), .B(n_372), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_401), .B(n_359), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_393), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_404), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_433), .B(n_360), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_406), .B(n_362), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_406), .B(n_365), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_396), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_433), .B(n_360), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_411), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_411), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_450), .B(n_353), .C(n_364), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_425), .B(n_361), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_391), .B(n_361), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_423), .A2(n_360), .B1(n_382), .B2(n_374), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_412), .A2(n_382), .B1(n_374), .B2(n_360), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_391), .B(n_383), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_407), .B(n_414), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_404), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_439), .B(n_374), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_427), .B(n_365), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_415), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_413), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_407), .B(n_362), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_413), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_405), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_389), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_392), .B(n_383), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_392), .B(n_383), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_387), .B(n_363), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_415), .Y(n_509) );
AND2x4_ASAP7_75t_SL g510 ( .A(n_405), .B(n_363), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_405), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_432), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_424), .A2(n_382), .B1(n_374), .B2(n_355), .Y(n_513) );
NAND4xp25_ASAP7_75t_L g514 ( .A(n_388), .B(n_382), .C(n_364), .D(n_367), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_432), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_414), .B(n_362), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_431), .B(n_370), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_440), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_422), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_439), .B(n_370), .Y(n_520) );
INVx3_ASAP7_75t_SL g521 ( .A(n_435), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_416), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_440), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_431), .B(n_370), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_449), .Y(n_525) );
INVx2_ASAP7_75t_SL g526 ( .A(n_424), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_416), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_446), .B(n_354), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_394), .B(n_355), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_437), .Y(n_530) );
AND2x2_ASAP7_75t_SL g531 ( .A(n_384), .B(n_367), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_390), .B(n_355), .Y(n_532) );
INVxp67_ASAP7_75t_SL g533 ( .A(n_454), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_390), .B(n_337), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_394), .B(n_337), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_421), .B(n_367), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_442), .B(n_445), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_421), .B(n_376), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_410), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_442), .B(n_366), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_445), .B(n_366), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_410), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_426), .B(n_376), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_417), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_417), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_531), .B(n_426), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_479), .B(n_403), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_536), .B(n_447), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_479), .B(n_403), .Y(n_549) );
NAND2x1_ASAP7_75t_L g550 ( .A(n_476), .B(n_419), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_525), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_470), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_458), .Y(n_553) );
OAI21xp33_ASAP7_75t_L g554 ( .A1(n_531), .A2(n_444), .B(n_438), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_468), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_510), .B(n_419), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_537), .B(n_446), .Y(n_557) );
INVxp67_ASAP7_75t_SL g558 ( .A(n_470), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_462), .B(n_447), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_463), .B(n_453), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_496), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_472), .B(n_443), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_526), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_519), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_472), .B(n_453), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_537), .B(n_428), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_526), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_473), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_474), .B(n_428), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_474), .B(n_429), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_532), .Y(n_571) );
AND2x4_ASAP7_75t_SL g572 ( .A(n_464), .B(n_384), .Y(n_572) );
AOI321xp33_ASAP7_75t_L g573 ( .A1(n_459), .A2(n_429), .A3(n_457), .B1(n_455), .B2(n_456), .C(n_448), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_521), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_475), .B(n_434), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_477), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_478), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_486), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_488), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_460), .A2(n_346), .B1(n_366), .B2(n_354), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_475), .B(n_448), .Y(n_581) );
NAND2x1p5_ASAP7_75t_L g582 ( .A(n_469), .B(n_346), .Y(n_582) );
NOR2xp33_ASAP7_75t_SL g583 ( .A(n_521), .B(n_354), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_467), .B(n_443), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_505), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_491), .B(n_457), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_506), .B(n_419), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_489), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_500), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_507), .B(n_419), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_510), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_509), .Y(n_592) );
AND3x1_ASAP7_75t_L g593 ( .A(n_459), .B(n_451), .C(n_420), .Y(n_593) );
AOI211xp5_ASAP7_75t_L g594 ( .A1(n_490), .A2(n_385), .B(n_384), .C(n_436), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_535), .B(n_385), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_461), .B(n_451), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_539), .B(n_456), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_466), .B(n_16), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_512), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_492), .B(n_385), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_515), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_529), .B(n_420), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_495), .B(n_436), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_518), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_542), .B(n_441), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_483), .B(n_436), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_485), .B(n_17), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_483), .B(n_402), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_534), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_508), .B(n_402), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_471), .A2(n_354), .B1(n_366), .B2(n_402), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_480), .B(n_441), .Y(n_612) );
OAI322xp33_ASAP7_75t_L g613 ( .A1(n_502), .A2(n_454), .A3(n_430), .B1(n_376), .B2(n_375), .C1(n_301), .C2(n_17), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_523), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_465), .Y(n_615) );
NAND2x1_ASAP7_75t_L g616 ( .A(n_508), .B(n_430), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_530), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_465), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_487), .B(n_366), .Y(n_619) );
BUFx2_ASAP7_75t_L g620 ( .A(n_508), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_574), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_574), .Y(n_622) );
NAND3xp33_ASAP7_75t_SL g623 ( .A(n_594), .B(n_471), .C(n_528), .Y(n_623) );
OAI22xp33_ASAP7_75t_SL g624 ( .A1(n_616), .A2(n_550), .B1(n_591), .B2(n_585), .Y(n_624) );
OAI322xp33_ASAP7_75t_L g625 ( .A1(n_607), .A2(n_516), .A3(n_484), .B1(n_499), .B2(n_538), .C1(n_493), .C2(n_524), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_584), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_620), .B(n_557), .Y(n_627) );
OAI21xp5_ASAP7_75t_SL g628 ( .A1(n_591), .A2(n_514), .B(n_528), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_593), .A2(n_511), .B1(n_504), .B2(n_354), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_593), .A2(n_487), .B1(n_498), .B2(n_543), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_594), .A2(n_585), .B1(n_556), .B2(n_564), .Y(n_631) );
OAI21xp5_ASAP7_75t_SL g632 ( .A1(n_556), .A2(n_504), .B(n_511), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_606), .B(n_520), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_608), .B(n_520), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_547), .B(n_543), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_561), .B(n_517), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_562), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_573), .A2(n_494), .B1(n_533), .B2(n_513), .C(n_498), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_562), .Y(n_639) );
AOI31xp33_ASAP7_75t_L g640 ( .A1(n_580), .A2(n_533), .A3(n_454), .B(n_494), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_547), .B(n_481), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_613), .A2(n_545), .B1(n_544), .B2(n_481), .C(n_482), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_558), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_617), .Y(n_644) );
OAI32xp33_ASAP7_75t_L g645 ( .A1(n_582), .A2(n_540), .A3(n_541), .B1(n_544), .B2(n_545), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_568), .Y(n_646) );
INVxp33_ASAP7_75t_L g647 ( .A(n_598), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_554), .A2(n_527), .B1(n_522), .B2(n_503), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_615), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_566), .B(n_527), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_551), .Y(n_651) );
AOI32xp33_ASAP7_75t_L g652 ( .A1(n_546), .A2(n_503), .A3(n_501), .B1(n_497), .B2(n_482), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_600), .B(n_522), .Y(n_653) );
O2A1O1Ixp5_ASAP7_75t_L g654 ( .A1(n_613), .A2(n_501), .B(n_497), .C(n_375), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g655 ( .A1(n_580), .A2(n_334), .B(n_366), .C(n_354), .Y(n_655) );
INVx2_ASAP7_75t_SL g656 ( .A(n_572), .Y(n_656) );
OAI32xp33_ASAP7_75t_L g657 ( .A1(n_582), .A2(n_375), .A3(n_366), .B1(n_354), .B2(n_327), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_554), .A2(n_366), .B1(n_354), .B2(n_327), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_603), .B(n_327), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_573), .B(n_327), .C(n_167), .Y(n_660) );
OAI211xp5_ASAP7_75t_SL g661 ( .A1(n_553), .A2(n_18), .B(n_19), .C(n_21), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_587), .A2(n_334), .B1(n_167), .B2(n_18), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_555), .B(n_19), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_549), .B(n_22), .Y(n_664) );
INVx2_ASAP7_75t_SL g665 ( .A(n_610), .Y(n_665) );
OAI21xp33_ASAP7_75t_L g666 ( .A1(n_597), .A2(n_23), .B(n_24), .Y(n_666) );
OAI21xp33_ASAP7_75t_L g667 ( .A1(n_575), .A2(n_25), .B(n_26), .Y(n_667) );
INVx2_ASAP7_75t_SL g668 ( .A(n_656), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_631), .A2(n_590), .B1(n_571), .B2(n_609), .Y(n_669) );
OAI22xp5_ASAP7_75t_SL g670 ( .A1(n_660), .A2(n_610), .B1(n_611), .B2(n_552), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_624), .A2(n_583), .B(n_611), .Y(n_671) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_660), .A2(n_599), .B1(n_579), .B2(n_614), .C1(n_578), .C2(n_588), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_621), .A2(n_619), .B1(n_563), .B2(n_567), .Y(n_673) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_628), .A2(n_605), .B1(n_583), .B2(n_589), .C(n_604), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_622), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_654), .A2(n_605), .B(n_569), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_637), .B(n_576), .Y(n_677) );
OAI21xp33_ASAP7_75t_SL g678 ( .A1(n_640), .A2(n_570), .B(n_595), .Y(n_678) );
NAND3xp33_ASAP7_75t_SL g679 ( .A(n_632), .B(n_596), .C(n_565), .Y(n_679) );
AOI21xp33_ASAP7_75t_L g680 ( .A1(n_647), .A2(n_601), .B(n_592), .Y(n_680) );
NAND4xp25_ASAP7_75t_L g681 ( .A(n_623), .B(n_602), .C(n_560), .D(n_577), .Y(n_681) );
NAND4xp25_ASAP7_75t_SL g682 ( .A(n_630), .B(n_581), .C(n_548), .D(n_586), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_639), .B(n_559), .Y(n_683) );
NOR4xp25_ASAP7_75t_SL g684 ( .A(n_638), .B(n_612), .C(n_618), .D(n_32), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g685 ( .A1(n_665), .A2(n_185), .B1(n_30), .B2(n_35), .Y(n_685) );
AOI311xp33_ASAP7_75t_L g686 ( .A1(n_624), .A2(n_27), .A3(n_37), .B(n_38), .C(n_39), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_649), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_625), .A2(n_42), .B1(n_43), .B2(n_44), .C(n_45), .Y(n_688) );
O2A1O1Ixp33_ASAP7_75t_SL g689 ( .A1(n_643), .A2(n_48), .B(n_49), .C(n_50), .Y(n_689) );
OAI21xp33_ASAP7_75t_L g690 ( .A1(n_652), .A2(n_52), .B(n_56), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_646), .Y(n_691) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_663), .A2(n_64), .B(n_65), .C(n_67), .Y(n_692) );
NOR5xp2_ASAP7_75t_L g693 ( .A(n_645), .B(n_68), .C(n_69), .D(n_71), .E(n_73), .Y(n_693) );
NAND4xp25_ASAP7_75t_SL g694 ( .A(n_655), .B(n_75), .C(n_76), .D(n_77), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_625), .A2(n_79), .B1(n_81), .B2(n_84), .C(n_88), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_651), .B(n_89), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_626), .B(n_90), .Y(n_697) );
OAI21xp33_ASAP7_75t_L g698 ( .A1(n_636), .A2(n_93), .B(n_95), .Y(n_698) );
O2A1O1Ixp5_ASAP7_75t_SL g699 ( .A1(n_644), .A2(n_96), .B(n_98), .C(n_99), .Y(n_699) );
OAI21xp5_ASAP7_75t_L g700 ( .A1(n_629), .A2(n_100), .B(n_102), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_661), .B(n_667), .C(n_664), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_642), .B(n_648), .C(n_662), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_655), .A2(n_627), .B(n_666), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_657), .A2(n_650), .B1(n_641), .B2(n_635), .C(n_653), .Y(n_704) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_658), .A2(n_633), .B(n_634), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_672), .B(n_702), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_688), .B(n_695), .C(n_672), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_678), .B(n_704), .C(n_671), .Y(n_708) );
AND2x4_ASAP7_75t_L g709 ( .A(n_668), .B(n_675), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_676), .B(n_691), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_L g711 ( .A1(n_681), .A2(n_679), .B(n_674), .C(n_705), .Y(n_711) );
AO221x1_ASAP7_75t_L g712 ( .A1(n_670), .A2(n_685), .B1(n_686), .B2(n_682), .C(n_684), .Y(n_712) );
AO221x2_ASAP7_75t_L g713 ( .A1(n_708), .A2(n_703), .B1(n_700), .B2(n_669), .C(n_683), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_706), .B(n_701), .C(n_690), .D(n_692), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_707), .B(n_696), .C(n_694), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_711), .B(n_697), .C(n_698), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_714), .B(n_709), .Y(n_717) );
AND2x4_ASAP7_75t_L g718 ( .A(n_715), .B(n_673), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_716), .B(n_710), .Y(n_719) );
INVx1_ASAP7_75t_SL g720 ( .A(n_717), .Y(n_720) );
INVx4_ASAP7_75t_L g721 ( .A(n_718), .Y(n_721) );
XOR2xp5_ASAP7_75t_L g722 ( .A(n_720), .B(n_719), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_721), .A2(n_713), .B1(n_718), .B2(n_712), .Y(n_723) );
AOI21x1_ASAP7_75t_L g724 ( .A1(n_722), .A2(n_677), .B(n_687), .Y(n_724) );
AO21x2_ASAP7_75t_L g725 ( .A1(n_724), .A2(n_723), .B(n_680), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_725), .B(n_699), .Y(n_726) );
OR2x6_ASAP7_75t_L g727 ( .A(n_726), .B(n_659), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_727), .A2(n_689), .B(n_693), .Y(n_728) );
endmodule