module fake_jpeg_3347_n_177 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx8_ASAP7_75t_SL g58 ( 
.A(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_2),
.B(n_19),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_57),
.Y(n_61)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

HAxp5_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_0),
.CON(n_66),
.SN(n_66)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_1),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_65),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_80),
.Y(n_82)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_55),
.B1(n_45),
.B2(n_43),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_41),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_65),
.B1(n_62),
.B2(n_55),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_95),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_41),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_92),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_49),
.B1(n_53),
.B2(n_45),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_91),
.B1(n_96),
.B2(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_42),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_66),
.B(n_43),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_77),
.B1(n_75),
.B2(n_42),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_74),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_54),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_109),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_105),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_48),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_46),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_59),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_3),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_4),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_119),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_84),
.C(n_52),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_134),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_20),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_100),
.B1(n_98),
.B2(n_112),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_128),
.B1(n_9),
.B2(n_10),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_125),
.B(n_126),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_4),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_52),
.B1(n_44),
.B2(n_7),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_5),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_132),
.B(n_9),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_44),
.B(n_6),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_135),
.A2(n_5),
.B(n_8),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_40),
.B(n_21),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_143),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_145),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_39),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_141),
.C(n_128),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_118),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_11),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_152),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_134),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_131),
.B1(n_127),
.B2(n_120),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_149),
.B1(n_136),
.B2(n_148),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_160),
.C(n_138),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_24),
.C(n_37),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_159),
.B1(n_154),
.B2(n_12),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_137),
.C(n_144),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_158),
.B(n_161),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_166),
.C(n_157),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_140),
.C(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_168),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_163),
.C(n_25),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_23),
.B(n_36),
.Y(n_173)
);

AOI21x1_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_172),
.B(n_18),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_17),
.B(n_34),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_16),
.B1(n_27),
.B2(n_13),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_14),
.Y(n_177)
);


endmodule