module real_jpeg_32342_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_641, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_641;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_578;
wire n_332;
wire n_366;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_0),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_0),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_0),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_0),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_54),
.B1(n_58),
.B2(n_61),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_1),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_1),
.A2(n_61),
.B1(n_132),
.B2(n_135),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_1),
.A2(n_61),
.B1(n_341),
.B2(n_343),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_1),
.A2(n_61),
.B1(n_578),
.B2(n_582),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_2),
.A2(n_144),
.B(n_149),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_2),
.B(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_2),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_2),
.B(n_206),
.Y(n_488)
);

OAI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_2),
.A2(n_125),
.B1(n_499),
.B2(n_516),
.Y(n_515)
);

OAI32xp33_ASAP7_75t_L g536 ( 
.A1(n_2),
.A2(n_181),
.A3(n_432),
.B1(n_537),
.B2(n_538),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_2),
.A2(n_177),
.B1(n_285),
.B2(n_335),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_4),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_4),
.B(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_4),
.A2(n_85),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_4),
.A2(n_85),
.B1(n_328),
.B2(n_332),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_SL g566 ( 
.A1(n_4),
.A2(n_85),
.B1(n_567),
.B2(n_568),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_5),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_5),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_167),
.B1(n_214),
.B2(n_217),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_5),
.A2(n_167),
.B1(n_232),
.B2(n_316),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_5),
.A2(n_167),
.B1(n_425),
.B2(n_427),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_6),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_6),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_6),
.A2(n_199),
.B1(n_319),
.B2(n_322),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_6),
.A2(n_164),
.B1(n_199),
.B2(n_417),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_6),
.A2(n_199),
.B1(n_479),
.B2(n_482),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_7),
.A2(n_98),
.B1(n_101),
.B2(n_106),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_7),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_7),
.A2(n_106),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_7),
.A2(n_106),
.B1(n_248),
.B2(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_7),
.A2(n_106),
.B1(n_231),
.B2(n_384),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_10),
.Y(n_120)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_11),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_11),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_11),
.A2(n_158),
.B1(n_241),
.B2(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_11),
.A2(n_158),
.B1(n_457),
.B2(n_461),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_11),
.A2(n_158),
.B1(n_500),
.B2(n_505),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_12),
.A2(n_170),
.B1(n_171),
.B2(n_177),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_12),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_12),
.A2(n_170),
.B1(n_228),
.B2(n_231),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_12),
.A2(n_170),
.B1(n_367),
.B2(n_492),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_12),
.A2(n_170),
.B1(n_295),
.B2(n_509),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_13),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_13),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_13),
.A2(n_121),
.B1(n_304),
.B2(n_309),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_13),
.A2(n_121),
.B1(n_373),
.B2(n_375),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_13),
.A2(n_121),
.B1(n_567),
.B2(n_598),
.Y(n_597)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_14),
.Y(n_81)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_14),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_15),
.A2(n_54),
.B1(n_58),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_15),
.A2(n_64),
.B1(n_295),
.B2(n_298),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_15),
.A2(n_64),
.B1(n_101),
.B2(n_366),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_15),
.A2(n_64),
.B1(n_578),
.B2(n_604),
.Y(n_603)
);

CKINVDCx11_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_17),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_17),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_18),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_18),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_21),
.B(n_24),
.Y(n_20)
);

BUFx12f_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_629),
.B(n_637),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_66),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_26),
.B(n_638),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_65),
.Y(n_27)
);

INVxp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_29),
.B(n_622),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_29),
.B(n_622),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_29),
.B(n_639),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_SL g65 ( 
.A1(n_30),
.A2(n_62),
.B(n_63),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_30),
.A2(n_62),
.B1(n_143),
.B2(n_154),
.Y(n_142)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_30),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_30),
.A2(n_62),
.B1(n_314),
.B2(n_318),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_30),
.A2(n_62),
.B1(n_227),
.B2(n_318),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_L g392 ( 
.A1(n_30),
.A2(n_62),
.B1(n_227),
.B2(n_318),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_30),
.A2(n_62),
.B1(n_596),
.B2(n_597),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_30),
.A2(n_53),
.B1(n_62),
.B2(n_597),
.Y(n_620)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_31),
.A2(n_225),
.B1(n_315),
.B2(n_383),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_44),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_36),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_36),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_36),
.Y(n_321)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_36),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_38),
.Y(n_240)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_39),
.Y(n_157)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_39),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_40),
.Y(n_153)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

AOI22x1_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_48),
.Y(n_182)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_48),
.Y(n_204)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_48),
.Y(n_243)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_48),
.Y(n_439)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_49),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_51),
.Y(n_190)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_57),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_60),
.Y(n_386)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_62),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_62),
.B(n_285),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g639 ( 
.A(n_65),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_559),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_405),
.B(n_554),
.Y(n_67)
);

NAND4xp25_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_286),
.C(n_387),
.D(n_398),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_262),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_70),
.B(n_262),
.Y(n_556)
);

XNOR2x1_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_208),
.Y(n_70)
);

XNOR2x1_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_140),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_72),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_117),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_73),
.B(n_117),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_84),
.B1(n_97),
.B2(n_107),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_74),
.A2(n_97),
.B1(n_107),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_74),
.A2(n_107),
.B1(n_163),
.B2(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_74),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_74),
.A2(n_107),
.B1(n_490),
.B2(n_491),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_74),
.B(n_285),
.Y(n_513)
);

AO21x1_ASAP7_75t_L g573 ( 
.A1(n_74),
.A2(n_107),
.B(n_365),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_75),
.Y(n_302)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AO21x2_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_108),
.B(n_113),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_76)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_77),
.Y(n_299)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_78),
.Y(n_279)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_79),
.Y(n_259)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_84),
.A2(n_107),
.B1(n_301),
.B2(n_303),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_91),
.Y(n_84)
);

BUFx2_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_88),
.Y(n_455)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_96),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_96),
.Y(n_419)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_96),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_100),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_104),
.Y(n_342)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_104),
.Y(n_368)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_105),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_107),
.A2(n_301),
.B1(n_303),
.B2(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_107),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_112),
.Y(n_308)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_112),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_113),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_125),
.B1(n_131),
.B2(n_137),
.Y(n_117)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_118),
.Y(n_251)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_119),
.Y(n_466)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_120),
.Y(n_260)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_120),
.Y(n_504)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_125),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_125),
.A2(n_131),
.B1(n_292),
.B2(n_294),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_125),
.A2(n_478),
.B1(n_484),
.B2(n_486),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_125),
.A2(n_499),
.B1(n_508),
.B2(n_512),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

BUFx4f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_128),
.Y(n_428)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_130),
.Y(n_282)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_130),
.Y(n_297)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_130),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_130),
.Y(n_483)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_130),
.Y(n_507)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_138),
.Y(n_283)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g430 ( 
.A(n_139),
.Y(n_430)
);

INVx8_ASAP7_75t_L g512 ( 
.A(n_139),
.Y(n_512)
);

INVxp33_ASAP7_75t_L g401 ( 
.A(n_140),
.Y(n_401)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_161),
.C(n_168),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_142),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_144),
.Y(n_246)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_148),
.Y(n_599)
);

AO21x1_ASAP7_75t_L g235 ( 
.A1(n_149),
.A2(n_236),
.B(n_244),
.Y(n_235)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_152),
.Y(n_570)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_154),
.Y(n_223)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_161),
.A2(n_162),
.B1(n_168),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_168),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_180),
.B1(n_198),
.B2(n_205),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_169),
.A2(n_180),
.B1(n_205),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_175),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_176),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_176),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_179),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_198),
.B1(n_213),
.B2(n_219),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_180),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_180),
.A2(n_213),
.B1(n_219),
.B2(n_334),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_180),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_180),
.A2(n_219),
.B1(n_270),
.B2(n_541),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_180),
.A2(n_219),
.B1(n_576),
.B2(n_577),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_180),
.A2(n_219),
.B1(n_577),
.B2(n_603),
.Y(n_602)
);

AO21x2_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_186),
.B(n_191),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g431 ( 
.A1(n_181),
.A2(n_432),
.B(n_438),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_182),
.Y(n_332)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_190),
.Y(n_331)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_190),
.Y(n_374)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.Y(n_191)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_SL g584 ( 
.A(n_201),
.Y(n_584)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AO22x2_ASAP7_75t_L g326 ( 
.A1(n_206),
.A2(n_327),
.B1(n_333),
.B2(n_336),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_206),
.A2(n_327),
.B1(n_372),
.B2(n_377),
.Y(n_371)
);

OAI21xp33_ASAP7_75t_SL g618 ( 
.A1(n_206),
.A2(n_377),
.B(n_619),
.Y(n_618)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_208),
.B(n_400),
.C(n_401),
.Y(n_399)
);

XNOR2x1_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_234),
.Y(n_208)
);

OAI21x1_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_220),
.B(n_233),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_211),
.B(n_234),
.C(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_222),
.Y(n_233)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_216),
.Y(n_335)
);

INVx3_ASAP7_75t_SL g248 ( 
.A(n_217),
.Y(n_248)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_222),
.Y(n_394)
);

AOI22x1_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_224),
.A2(n_225),
.B1(n_383),
.B2(n_566),
.Y(n_565)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_249),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_235),
.A2(n_249),
.B1(n_250),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_235),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_238),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_245),
.C(n_247),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_257),
.B2(n_261),
.Y(n_250)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_253),
.B(n_285),
.Y(n_518)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_255),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_256),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_261),
.B1(n_277),
.B2(n_283),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OA21x2_ASAP7_75t_L g346 ( 
.A1(n_261),
.A2(n_347),
.B(n_348),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_261),
.A2(n_277),
.B1(n_424),
.B2(n_429),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_261),
.A2(n_523),
.B1(n_524),
.B2(n_525),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.C(n_268),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_263),
.B(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_266),
.B(n_268),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_275),
.C(n_284),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_269),
.B(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_275),
.A2(n_276),
.B1(n_284),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_284),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_285),
.B(n_433),
.Y(n_432)
);

NAND3xp33_ASAP7_75t_L g438 ( 
.A(n_285),
.B(n_439),
.C(n_440),
.Y(n_438)
);

OAI21xp33_ASAP7_75t_SL g450 ( 
.A1(n_285),
.A2(n_451),
.B(n_453),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_285),
.B(n_454),
.Y(n_453)
);

A2O1A1O1Ixp25_ASAP7_75t_L g554 ( 
.A1(n_286),
.A2(n_387),
.B(n_555),
.C(n_557),
.D(n_558),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_357),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_287),
.B(n_357),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_337),
.C(n_349),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_289),
.B(n_338),
.Y(n_397)
);

XNOR2x1_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_312),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_290),
.B(n_359),
.C(n_360),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_300),
.Y(n_290)
);

XOR2x2_ASAP7_75t_L g395 ( 
.A(n_291),
.B(n_300),
.Y(n_395)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_296),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_298),
.Y(n_519)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_302),
.A2(n_364),
.B1(n_369),
.B2(n_370),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_302),
.A2(n_369),
.B1(n_416),
.B2(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_311),
.Y(n_452)
);

XNOR2x1_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_326),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_319),
.Y(n_567)
);

INVx11_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx12f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_326),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_345),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_346),
.Y(n_379)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_340),
.Y(n_370)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_344),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_345),
.A2(n_346),
.B1(n_381),
.B2(n_382),
.Y(n_380)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_346),
.A2(n_587),
.B1(n_588),
.B2(n_641),
.Y(n_586)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_347),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.C(n_354),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_391),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_352),
.A2(n_355),
.B1(n_356),
.B2(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_358),
.B(n_625),
.C(n_626),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_378),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_362),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_371),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_363),
.B(n_371),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_369),
.A2(n_450),
.B1(n_456),
.B2(n_462),
.Y(n_449)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_372),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_378),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_379),
.Y(n_587)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_382),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_396),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_388),
.B(n_396),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_393),
.C(n_395),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_390),
.B(n_404),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_395),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_399),
.B(n_402),
.C(n_556),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_443),
.B(n_553),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_407),
.B(n_409),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_414),
.C(n_420),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_410),
.A2(n_411),
.B1(n_547),
.B2(n_548),
.Y(n_546)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_414),
.A2(n_420),
.B1(n_421),
.B2(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_414),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_419),
.Y(n_492)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_431),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_422),
.A2(n_423),
.B1(n_431),
.B2(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_424),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_426),
.Y(n_474)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_439),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_440),
.Y(n_538)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_545),
.B(n_552),
.Y(n_443)
);

AOI21x1_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_531),
.B(n_544),
.Y(n_444)
);

OAI21x1_ASAP7_75t_SL g445 ( 
.A1(n_446),
.A2(n_495),
.B(n_530),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_476),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_447),
.B(n_476),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_463),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_448),
.A2(n_449),
.B1(n_463),
.B2(n_464),
.Y(n_528)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_453),
.Y(n_471)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_456),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx3_ASAP7_75t_SL g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_465),
.A2(n_471),
.B1(n_472),
.B2(n_475),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_487),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_477),
.B(n_489),
.C(n_493),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_478),
.Y(n_524)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_483),
.Y(n_511)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_489),
.B1(n_493),
.B2(n_494),
.Y(n_487)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_488),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_489),
.Y(n_494)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_491),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_496),
.A2(n_521),
.B(n_529),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_497),
.A2(n_514),
.B(n_520),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_513),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_498),
.B(n_513),
.Y(n_520)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_508),
.Y(n_523)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_515),
.B(n_517),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_518),
.B(n_519),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_528),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_528),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_533),
.Y(n_531)
);

NOR2x1_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_533),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_539),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_542),
.C(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_542),
.Y(n_539)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_540),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_550),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_546),
.B(n_550),
.Y(n_552)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

NOR3xp33_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_607),
.C(n_623),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_561),
.A2(n_633),
.B(n_634),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_562),
.B(n_589),
.Y(n_561)
);

NOR2xp67_ASAP7_75t_L g634 ( 
.A(n_562),
.B(n_589),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_585),
.C(n_586),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g628 ( 
.A(n_564),
.B(n_585),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_571),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_565),
.B(n_572),
.C(n_575),
.Y(n_590)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_565),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_566),
.Y(n_596)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx3_ASAP7_75t_SL g569 ( 
.A(n_570),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_572),
.A2(n_573),
.B1(n_574),
.B2(n_575),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_572),
.A2(n_573),
.B1(n_601),
.B2(n_602),
.Y(n_600)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_573),
.B(n_595),
.C(n_602),
.Y(n_615)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_586),
.B(n_628),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_590),
.B(n_591),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_590),
.B(n_592),
.C(n_594),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_592),
.B(n_594),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_SL g594 ( 
.A(n_595),
.B(n_600),
.Y(n_594)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_603),
.Y(n_619)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx8_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_608),
.B(n_621),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_609),
.A2(n_632),
.B(n_635),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_610),
.B(n_612),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_611),
.B(n_613),
.Y(n_635)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_614),
.A2(n_615),
.B1(n_616),
.B2(n_617),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_614),
.B(n_618),
.C(n_620),
.Y(n_622)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_618),
.B(n_620),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_621),
.A2(n_631),
.B(n_636),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_624),
.B(n_627),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_624),
.B(n_627),
.Y(n_633)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);


endmodule