module fake_aes_1865_n_20 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_20);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_20;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
NAND2xp5_ASAP7_75t_L g12 ( .A(n_11), .B(n_3), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_5), .B(n_1), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_2), .B(n_7), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_6), .B(n_8), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
NAND3xp33_ASAP7_75t_SL g18 ( .A(n_17), .B(n_12), .C(n_13), .Y(n_18) );
AOI22xp5_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_16), .B1(n_15), .B2(n_0), .Y(n_19) );
AOI221x1_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_0), .B1(n_4), .B2(n_9), .C(n_10), .Y(n_20) );
endmodule