module real_jpeg_6350_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_1),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_1),
.A2(n_28),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_1),
.A2(n_28),
.B1(n_171),
.B2(n_174),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_1),
.B(n_92),
.Y(n_225)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_1),
.A2(n_201),
.B(n_249),
.C(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_1),
.B(n_274),
.C(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_1),
.B(n_129),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_1),
.B(n_22),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_1),
.B(n_48),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_2),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_2),
.A2(n_104),
.B1(n_209),
.B2(n_212),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_2),
.A2(n_104),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_2),
.A2(n_104),
.B1(n_284),
.B2(n_286),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_4),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_5),
.Y(n_152)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_5),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_6),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_6),
.A2(n_44),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_6),
.A2(n_44),
.B1(n_123),
.B2(n_126),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_6),
.A2(n_44),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_7),
.Y(n_117)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_9),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_9),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_9),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_9),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_10),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_10),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_10),
.A2(n_61),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_10),
.A2(n_61),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_11),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_352),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_216),
.B(n_350),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_185),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_15),
.B(n_185),
.Y(n_351)
);

BUFx24_ASAP7_75t_SL g380 ( 
.A(n_15),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_149),
.CI(n_158),
.CON(n_15),
.SN(n_15)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_16),
.B(n_149),
.C(n_158),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_82),
.B2(n_83),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_17),
.B(n_84),
.C(n_120),
.Y(n_378)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_19),
.B(n_46),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_20),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_21),
.A2(n_33),
.B(n_161),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_24),
.A2(n_34),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_24),
.B(n_34),
.Y(n_227)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_27),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_28),
.A2(n_87),
.B(n_89),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_28),
.B(n_90),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_28),
.A2(n_251),
.B(n_254),
.Y(n_250)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_32),
.B(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_40),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_34),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_34),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_37),
.Y(n_163)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_40),
.B(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_41),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_42),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_43),
.Y(n_285)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_45),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_55),
.B(n_64),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_47),
.A2(n_155),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_47),
.B(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_48),
.B(n_65),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_48),
.B(n_262),
.Y(n_278)
);

AO22x1_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_55),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_60),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_64),
.B(n_278),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_64),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_71),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_67),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_67),
.B(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_70),
.Y(n_256)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_71),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_71),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_80),
.A2(n_131),
.B1(n_134),
.B2(n_136),
.Y(n_130)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_80),
.Y(n_264)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_120),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_101),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_92),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_86),
.B(n_109),
.Y(n_232)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_86),
.Y(n_367)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_89),
.Y(n_198)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_92),
.B(n_102),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_92),
.B(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_92),
.Y(n_366)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_98),
.B2(n_100),
.Y(n_92)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_93),
.Y(n_197)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx8_ASAP7_75t_L g372 ( 
.A(n_95),
.Y(n_372)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_97),
.Y(n_201)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_97),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_97),
.Y(n_214)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_99),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_101),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_109),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI32xp33_ASAP7_75t_L g194 ( 
.A1(n_106),
.A2(n_195),
.A3(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_109),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_109),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_118),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_138),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_121),
.B(n_207),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_129),
.Y(n_121)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_122),
.Y(n_237)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_128),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_139),
.B(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_129),
.B(n_208),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_129),
.A2(n_236),
.B(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_130),
.B(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_132),
.Y(n_253)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_133),
.Y(n_249)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_138),
.B(n_238),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_139),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_140),
.B(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_145),
.Y(n_206)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_153),
.B1(n_154),
.B2(n_157),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_150),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_150),
.A2(n_157),
.B1(n_248),
.B2(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_150),
.B(n_154),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_150),
.A2(n_157),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_156),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_156),
.B(n_261),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_175),
.C(n_177),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_160),
.B(n_168),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_165),
.B(n_166),
.Y(n_160)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_166),
.B(n_282),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_169),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_170),
.Y(n_241)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_184),
.B(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_215),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_186),
.B(n_215),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_189),
.B(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_203),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_190),
.B(n_203),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_192),
.B(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_194),
.Y(n_229)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

INVx6_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_334),
.B(n_347),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_266),
.B(n_333),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_243),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_219),
.B(n_243),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_228),
.B2(n_229),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_222),
.B(n_228),
.C(n_230),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.C(n_226),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_245),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_226),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_227),
.B(n_298),
.Y(n_310)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_231),
.B(n_234),
.C(n_240),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_239),
.B1(n_240),
.B2(n_242),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.C(n_257),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_244),
.B(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_247),
.A2(n_257),
.B1(n_258),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_247),
.Y(n_330)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_248),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_260),
.B(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_327),
.B(n_332),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_317),
.B(n_326),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_292),
.B(n_316),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_279),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_279),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_277),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_272),
.B1(n_277),
.B2(n_295),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_287),
.Y(n_279)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_288),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_290),
.C(n_319),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_303),
.B(n_315),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_296),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_311),
.B(n_314),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_310),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_320),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_323),
.C(n_324),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_331),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_331),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_343),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_337),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_341),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_340),
.C(n_341),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_343),
.A2(n_348),
.B(n_349),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_344),
.B(n_346),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_379),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_355),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_378),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_368),
.B2(n_369),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_361),
.B2(n_362),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_366),
.B(n_367),
.Y(n_364)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_375),
.B(n_377),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_370),
.B(n_375),
.Y(n_377)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);


endmodule