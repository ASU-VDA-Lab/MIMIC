module real_jpeg_3222_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_0),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_26),
.B1(n_60),
.B2(n_61),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_1),
.A2(n_26),
.B1(n_32),
.B2(n_37),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_1),
.A2(n_26),
.B1(n_76),
.B2(n_78),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_4),
.A2(n_27),
.B1(n_29),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_4),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_4),
.A2(n_32),
.B1(n_37),
.B2(n_85),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_85),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_4),
.A2(n_76),
.B1(n_78),
.B2(n_85),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_5),
.A2(n_41),
.B1(n_60),
.B2(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_5),
.A2(n_41),
.B1(n_76),
.B2(n_78),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_5),
.A2(n_32),
.B1(n_37),
.B2(n_41),
.Y(n_150)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_6),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_7),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_7),
.A2(n_32),
.B1(n_37),
.B2(n_115),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_7),
.A2(n_60),
.B1(n_61),
.B2(n_115),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_7),
.A2(n_76),
.B1(n_78),
.B2(n_115),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_9),
.A2(n_27),
.B1(n_29),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_9),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_9),
.A2(n_32),
.B1(n_37),
.B2(n_177),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_177),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_9),
.A2(n_76),
.B1(n_78),
.B2(n_177),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_20),
.B(n_344),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_12),
.B(n_345),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_13),
.A2(n_32),
.B1(n_37),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_68),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_68),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_13),
.A2(n_68),
.B1(n_76),
.B2(n_78),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_14),
.A2(n_32),
.B1(n_37),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_14),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_65),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_65),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_14),
.A2(n_65),
.B1(n_76),
.B2(n_78),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_15),
.A2(n_27),
.B1(n_29),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_15),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_15),
.A2(n_32),
.B1(n_37),
.B2(n_137),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_137),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_15),
.A2(n_76),
.B1(n_78),
.B2(n_137),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_17),
.B(n_29),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_17),
.B(n_42),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_17),
.A2(n_37),
.B(n_57),
.C(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_17),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_17),
.B(n_59),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_17),
.A2(n_32),
.B1(n_37),
.B2(n_227),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_17),
.B(n_73),
.C(n_76),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_17),
.A2(n_60),
.B1(n_61),
.B2(n_227),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_17),
.B(n_105),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_17),
.B(n_94),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_46),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_44),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_43),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_23),
.B(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_24),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_24),
.B(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_40),
.B2(n_42),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_25),
.A2(n_30),
.B1(n_42),
.B2(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g197 ( 
.A1(n_27),
.A2(n_35),
.A3(n_37),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_27),
.A2(n_86),
.B(n_227),
.C(n_236),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_40),
.B(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_30),
.B(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_30),
.A2(n_42),
.B1(n_136),
.B2(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_31),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_31),
.A2(n_84),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_31),
.B(n_114),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_31),
.A2(n_86),
.B1(n_87),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_31),
.A2(n_112),
.B(n_191),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_31)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_32),
.B(n_38),
.Y(n_199)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_57),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

OAI21x1_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_339),
.B(n_341),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_327),
.B(n_338),
.Y(n_47)
);

AO21x1_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_153),
.B(n_324),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_140),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_116),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_51),
.B(n_116),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_97),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_81),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_53),
.A2(n_54),
.B(n_69),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_53),
.B(n_81),
.C(n_97),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_69),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_66),
.B1(n_67),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_55),
.A2(n_64),
.B1(n_66),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_55),
.A2(n_66),
.B1(n_91),
.B2(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_55),
.A2(n_193),
.B(n_195),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_55),
.A2(n_195),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_56),
.B(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_56),
.A2(n_59),
.B1(n_194),
.B2(n_211),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_56),
.A2(n_59),
.B(n_331),
.Y(n_330)
);

AO22x1_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_59),
.B(n_174),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_61),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_60),
.A2(n_63),
.B(n_227),
.Y(n_226)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_61),
.B(n_272),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_66),
.A2(n_133),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_66),
.A2(n_173),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_75),
.B1(n_79),
.B2(n_80),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_75),
.B1(n_79),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_70),
.A2(n_75),
.B1(n_220),
.B2(n_254),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_70),
.A2(n_222),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_71),
.A2(n_94),
.B1(n_110),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_71),
.A2(n_94),
.B1(n_131),
.B2(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_71),
.A2(n_219),
.B(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_71),
.B(n_223),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_75),
.A2(n_242),
.B(n_243),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_75),
.A2(n_243),
.B(n_254),
.Y(n_253)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_76),
.B(n_283),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_96),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_82),
.A2(n_83),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g151 ( 
.A(n_83),
.B(n_89),
.C(n_93),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_83),
.B(n_144),
.C(n_151),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_86),
.A2(n_135),
.B(n_138),
.Y(n_134)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_92),
.A2(n_93),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_93),
.B(n_145),
.C(n_149),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_94),
.B(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B(n_111),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_99),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_108),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_101),
.B1(n_111),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_100),
.A2(n_101),
.B1(n_108),
.B2(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_105),
.B(n_106),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_102),
.A2(n_105),
.B1(n_128),
.B2(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_102),
.A2(n_227),
.B(n_260),
.Y(n_284)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_103),
.A2(n_104),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_103),
.A2(n_104),
.B1(n_202),
.B2(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_103),
.B(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_103),
.A2(n_258),
.B(n_259),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_103),
.A2(n_104),
.B1(n_258),
.B2(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_104),
.A2(n_217),
.B(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_104),
.B(n_231),
.Y(n_260)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_105),
.A2(n_230),
.B(n_287),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_108),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.C(n_123),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_132),
.C(n_134),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_125),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_126),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_134),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_139),
.B(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_140),
.A2(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_152),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_141),
.B(n_152),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_151),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_146),
.Y(n_333)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_150),
.Y(n_331)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_178),
.B(n_323),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_155),
.B(n_158),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.C(n_175),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_166),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_167),
.B(n_169),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_168),
.Y(n_242)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

OAI21x1_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_204),
.B(n_322),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_180),
.B(n_182),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.C(n_189),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_183),
.B(n_187),
.Y(n_307)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_189),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_196),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_190),
.B(n_192),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_196),
.B(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_197),
.A2(n_200),
.B1(n_201),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI31xp33_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_304),
.A3(n_314),
.B(n_319),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_248),
.B(n_303),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_232),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_207),
.B(n_232),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.C(n_224),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_208),
.B(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_213),
.C(n_216),
.Y(n_247)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_218),
.B(n_224),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_228),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_244),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_233),
.B(n_245),
.C(n_247),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_234),
.B(n_239),
.C(n_240),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_298),
.B(n_302),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_267),
.B(n_297),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_261),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_261),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.C(n_256),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_257),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_265),
.C(n_266),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_279),
.B(n_296),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_275),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_275),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_270),
.A2(n_271),
.B1(n_273),
.B2(n_294),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_290),
.B(n_295),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_285),
.B(n_289),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_288),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_287),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_293),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_301),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_305),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_308),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.C(n_312),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_316),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_311),
.A2(n_312),
.B1(n_313),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_311),
.Y(n_317)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_318),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_337),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_337),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_336),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_334),
.C(n_336),
.Y(n_340)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_340),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);


endmodule