module fake_jpeg_2382_n_159 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_13),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_60),
.Y(n_63)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_41),
.B1(n_43),
.B2(n_40),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_62),
.B1(n_58),
.B2(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_49),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_52),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_60),
.C(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_63),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_78),
.Y(n_92)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_77),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_80),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_58),
.B1(n_56),
.B2(n_54),
.Y(n_81)
);

AOI22x1_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_84),
.B1(n_69),
.B2(n_60),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_83),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_49),
.C(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_85),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_44),
.B1(n_65),
.B2(n_70),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_60),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_101),
.B1(n_1),
.B2(n_2),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_77),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_53),
.B(n_50),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_101),
.B(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_102),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_53),
.B1(n_51),
.B2(n_39),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_45),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_5),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_119),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_107),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_0),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_115),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_1),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_121),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_2),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_11),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_93),
.B1(n_87),
.B2(n_88),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_3),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_120),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_21),
.C(n_37),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_4),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_10),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_6),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_121)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_116),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_116),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_30),
.B(n_20),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_14),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_23),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_131),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_120),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_134),
.A2(n_135),
.B1(n_132),
.B2(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_146),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_124),
.B(n_133),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_118),
.B(n_123),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_141),
.A2(n_135),
.B1(n_127),
.B2(n_134),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_147),
.A2(n_141),
.B1(n_136),
.B2(n_142),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_146),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_151),
.B(n_152),
.Y(n_153)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_137),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_150),
.B(n_144),
.Y(n_155)
);

NOR2xp67_ASAP7_75t_SL g156 ( 
.A(n_155),
.B(n_126),
.Y(n_156)
);

AOI21x1_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_126),
.B(n_32),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_31),
.B(n_35),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_36),
.Y(n_159)
);


endmodule