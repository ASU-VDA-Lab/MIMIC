module real_jpeg_23442_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_0),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_2),
.A2(n_25),
.B1(n_31),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_2),
.A2(n_52),
.B1(n_53),
.B2(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_3),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_3),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_3),
.B(n_53),
.C(n_55),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_3),
.B(n_78),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_3),
.A2(n_52),
.B1(n_53),
.B2(n_100),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_3),
.B(n_25),
.C(n_86),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_24),
.B(n_152),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_59),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_59),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_6),
.A2(n_25),
.B1(n_31),
.B2(n_59),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_8),
.A2(n_25),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_41),
.B1(n_62),
.B2(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_10),
.A2(n_25),
.B1(n_31),
.B2(n_62),
.Y(n_124)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_12),
.A2(n_37),
.B1(n_38),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_80),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_12),
.A2(n_25),
.B1(n_31),
.B2(n_80),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_14),
.Y(n_154)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_14),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_127),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_105),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_18),
.B(n_105),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_73),
.B2(n_74),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_49),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_23),
.A2(n_165),
.B1(n_167),
.B2(n_169),
.Y(n_164)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_24),
.A2(n_30),
.B1(n_70),
.B2(n_72),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_24),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_24),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_25),
.A2(n_31),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_31),
.B(n_179),
.Y(n_178)
);

AOI32xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.A3(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_38),
.B1(n_55),
.B2(n_56),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_68)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_38),
.B(n_118),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_94),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_66),
.C(n_69),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_57),
.B(n_60),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_53),
.B1(n_85),
.B2(n_86),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_53),
.B(n_161),
.Y(n_160)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_63),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_61),
.B(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_64),
.A2(n_136),
.B(n_137),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_72),
.A2(n_166),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_91),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_87),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_84),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_84),
.A2(n_87),
.B(n_133),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_84),
.B(n_100),
.Y(n_174)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_88),
.A2(n_113),
.B1(n_115),
.B2(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_96),
.B(n_102),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_103),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_100),
.B(n_101),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_100),
.B(n_154),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_116),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_107),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_116),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B(n_114),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_111),
.A2(n_114),
.B(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_119),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_123),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_141),
.B(n_190),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_138),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_129),
.B(n_138),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.C(n_134),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_184),
.B(n_189),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_162),
.B(n_183),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_156),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_156),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_149),
.C(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_160),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_172),
.B(n_182),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_170),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_177),
.B(n_181),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_175),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_188),
.Y(n_189)
);


endmodule