module fake_jpeg_27155_n_102 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx9p33_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_24),
.B(n_30),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_32),
.B1(n_11),
.B2(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_33),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_15),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_7),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_11),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_38),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_14),
.B1(n_18),
.B2(n_28),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_50),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_52),
.B1(n_54),
.B2(n_60),
.Y(n_64)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_28),
.B1(n_14),
.B2(n_20),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_56),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_20),
.B1(n_21),
.B2(n_29),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_12),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_12),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_21),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_44),
.B1(n_37),
.B2(n_39),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_55),
.B(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_41),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_44),
.B1(n_41),
.B2(n_23),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_71),
.B1(n_54),
.B2(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_70),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_44),
.B1(n_45),
.B2(n_10),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_70),
.A2(n_56),
.B1(n_57),
.B2(n_55),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_50),
.B(n_45),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_77),
.B(n_80),
.Y(n_82)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_79),
.C(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_67),
.Y(n_80)
);

AOI221xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_67),
.B1(n_71),
.B2(n_64),
.C(n_59),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_83),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_59),
.C(n_45),
.Y(n_83)
);

AOI21x1_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_76),
.B(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_91),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_77),
.B(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_94),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_90),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_97),
.B(n_98),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_96),
.B(n_27),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_99),
.Y(n_102)
);


endmodule