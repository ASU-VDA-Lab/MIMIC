module fake_jpeg_93_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_52),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_36),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_60),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_43),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_65),
.C(n_34),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_46),
.B1(n_45),
.B2(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_42),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_71),
.Y(n_79)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_76),
.Y(n_81)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_56),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_33),
.C(n_14),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_41),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_59),
.B1(n_45),
.B2(n_3),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_91),
.B1(n_67),
.B2(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_1),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_59),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_97),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_100),
.B1(n_106),
.B2(n_9),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_70),
.B1(n_76),
.B2(n_3),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_1),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_18),
.B1(n_32),
.B2(n_31),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_87),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_16),
.B1(n_30),
.B2(n_28),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_20),
.B(n_26),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_2),
.C(n_6),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_118),
.C(n_107),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_7),
.B(n_8),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_117),
.Y(n_129)
);

HAxp5_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_7),
.CON(n_113),
.SN(n_113)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_116),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_10),
.B(n_11),
.Y(n_118)
);

OA21x2_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_13),
.B(n_21),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_127),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_120),
.B(n_24),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_111),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_108),
.C(n_133),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_125),
.A2(n_111),
.B1(n_117),
.B2(n_115),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_130),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_126),
.C(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_112),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_129),
.B(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_136),
.B(n_126),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_105),
.B(n_113),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_25),
.Y(n_145)
);


endmodule