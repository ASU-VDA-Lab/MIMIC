module fake_netlist_5_2167_n_1650 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1650);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1650;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx2_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_112),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_0),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_13),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_81),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_36),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_106),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_25),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_7),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_130),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_132),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_11),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_95),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_110),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_57),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_78),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_60),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_54),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_59),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_68),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_111),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_10),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_32),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_88),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_93),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_145),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_79),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_87),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_32),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_0),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_46),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_21),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_43),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_61),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_143),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_84),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_39),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_33),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_75),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_42),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_43),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_28),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_49),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_67),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_116),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_105),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_149),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_9),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_73),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_80),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_58),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_7),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_63),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_18),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_118),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_115),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_91),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_135),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_18),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_14),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_131),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_50),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_9),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_62),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_97),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_121),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_24),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_65),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_5),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_141),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_52),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_11),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_109),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_13),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_17),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_113),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_83),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_144),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_3),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_69),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_101),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_140),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_152),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_1),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_15),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_98),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_129),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_74),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_146),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_27),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_72),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_12),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_26),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_86),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_5),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_82),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_92),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_21),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_45),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_3),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_8),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_134),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_45),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_56),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_137),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_94),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_147),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_4),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_122),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_12),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_128),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_36),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_37),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_77),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_34),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_123),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_24),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_124),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_108),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_16),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_138),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_64),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_40),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_41),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_27),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_41),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_42),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_22),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_76),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_37),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_40),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_30),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_266),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_177),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_180),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_230),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_227),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_272),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_154),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_230),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_182),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_230),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_230),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_177),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_153),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_155),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_230),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_210),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_187),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_265),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_187),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_293),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_244),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_155),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_183),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_236),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_156),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_228),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_265),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_168),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_189),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_250),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_196),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_265),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_161),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_207),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_208),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_215),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_242),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_162),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_246),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_232),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_178),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_184),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_251),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_159),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_252),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_262),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_185),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_276),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_280),
.Y(n_354)
);

INVxp33_ASAP7_75t_SL g355 ( 
.A(n_162),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_163),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_175),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_188),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_285),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_169),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_190),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_192),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_265),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_294),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_277),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_260),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_193),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_165),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_194),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_327),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_305),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_305),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_305),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_223),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_320),
.Y(n_379)
);

NOR2x1_ASAP7_75t_L g380 ( 
.A(n_304),
.B(n_173),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_310),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_316),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_310),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_357),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_346),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_352),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_305),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_175),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_305),
.Y(n_391)
);

INVxp33_ASAP7_75t_SL g392 ( 
.A(n_370),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_302),
.B(n_220),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_312),
.B(n_313),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_313),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_317),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_331),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_307),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_331),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_307),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_307),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_307),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_357),
.B(n_220),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_307),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_307),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_301),
.B(n_160),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_357),
.B(n_222),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_315),
.B(n_222),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_357),
.B(n_174),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_363),
.Y(n_414)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_357),
.B(n_176),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_329),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_302),
.B(n_260),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_363),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g420 ( 
.A(n_357),
.B(n_179),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_308),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_358),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_302),
.B(n_181),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_348),
.B(n_191),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_316),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_335),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_335),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_348),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_348),
.B(n_157),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_314),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_337),
.B(n_186),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_361),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_314),
.B(n_197),
.Y(n_434)
);

AND3x2_ASAP7_75t_L g435 ( 
.A(n_412),
.B(n_198),
.C(n_303),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_373),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_394),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_L g439 ( 
.A(n_390),
.B(n_362),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_383),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_372),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_394),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_404),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_394),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_394),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_432),
.B(n_301),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_373),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_385),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_408),
.Y(n_449)
);

OAI22xp33_ASAP7_75t_L g450 ( 
.A1(n_390),
.A2(n_309),
.B1(n_334),
.B2(n_323),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_408),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_425),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_408),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_371),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_368),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_371),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_425),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_371),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_392),
.B(n_345),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_373),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_392),
.B(n_345),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_355),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_386),
.B(n_306),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_379),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_379),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_377),
.B(n_157),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_373),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_323),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_378),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_387),
.B(n_306),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_378),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_L g474 ( 
.A(n_377),
.B(n_424),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_422),
.B(n_160),
.Y(n_475)
);

AOI21x1_ASAP7_75t_L g476 ( 
.A1(n_410),
.A2(n_202),
.B(n_200),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_412),
.B(n_325),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_414),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_423),
.B(n_325),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_433),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_383),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_383),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_407),
.B(n_311),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_377),
.B(n_160),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_379),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_381),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_421),
.Y(n_488)
);

OAI22xp33_ASAP7_75t_L g489 ( 
.A1(n_411),
.A2(n_234),
.B1(n_219),
.B2(n_221),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_407),
.B(n_237),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_385),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_382),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_411),
.B(n_237),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_417),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_397),
.Y(n_495)
);

AO21x2_ASAP7_75t_L g496 ( 
.A1(n_410),
.A2(n_216),
.B(n_205),
.Y(n_496)
);

AOI21x1_ASAP7_75t_L g497 ( 
.A1(n_399),
.A2(n_229),
.B(n_225),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_417),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_397),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_417),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_384),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_373),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_381),
.B(n_430),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_384),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_431),
.B(n_237),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_431),
.B(n_158),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_373),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_389),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_389),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_400),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_400),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_400),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_419),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_431),
.B(n_158),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_421),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_430),
.B(n_393),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_395),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_395),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_396),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_396),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_415),
.B(n_164),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_373),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_398),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_398),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_373),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_393),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_385),
.Y(n_530)
);

NAND3xp33_ASAP7_75t_L g531 ( 
.A(n_415),
.B(n_333),
.C(n_332),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_414),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_414),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_419),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_419),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_415),
.B(n_253),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_414),
.Y(n_537)
);

AND3x2_ASAP7_75t_L g538 ( 
.A(n_393),
.B(n_233),
.C(n_231),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_419),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_409),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_414),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_409),
.Y(n_542)
);

NAND3xp33_ASAP7_75t_L g543 ( 
.A(n_423),
.B(n_434),
.C(n_380),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_409),
.Y(n_544)
);

AND2x2_ASAP7_75t_SL g545 ( 
.A(n_404),
.B(n_238),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_409),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_414),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_409),
.Y(n_548)
);

AO22x2_ASAP7_75t_L g549 ( 
.A1(n_434),
.A2(n_248),
.B1(n_255),
.B2(n_256),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_413),
.Y(n_550)
);

INVx5_ASAP7_75t_L g551 ( 
.A(n_424),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_414),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_413),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_423),
.B(n_201),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_374),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_374),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_434),
.B(n_166),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_434),
.B(n_166),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_374),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_413),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_414),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_416),
.B(n_326),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_375),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_413),
.A2(n_226),
.B1(n_263),
.B2(n_283),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_427),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_404),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_375),
.Y(n_567)
);

AND3x2_ASAP7_75t_L g568 ( 
.A(n_404),
.B(n_275),
.C(n_273),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_385),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_427),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_413),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_416),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_375),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_380),
.B(n_343),
.C(n_365),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_391),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_399),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_418),
.A2(n_239),
.B1(n_241),
.B2(n_209),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_376),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_519),
.B(n_401),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_529),
.B(n_401),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_463),
.B(n_167),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_443),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_488),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_443),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_529),
.B(n_402),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_545),
.B(n_427),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_545),
.B(n_427),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_494),
.B(n_167),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_494),
.B(n_290),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_491),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_436),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_452),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_436),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_L g594 ( 
.A(n_460),
.B(n_418),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_498),
.B(n_402),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_449),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_498),
.B(n_500),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_500),
.B(n_406),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_536),
.B(n_478),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_545),
.B(n_406),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_449),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_438),
.B(n_376),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_438),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_458),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_458),
.B(n_318),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_451),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_524),
.A2(n_531),
.B1(n_496),
.B2(n_549),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_442),
.B(n_376),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_566),
.A2(n_531),
.B1(n_439),
.B2(n_572),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_442),
.B(n_376),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_444),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_444),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_483),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_445),
.B(n_376),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_451),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_496),
.A2(n_424),
.B1(n_265),
.B2(n_297),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_445),
.B(n_388),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_550),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_491),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_550),
.B(n_388),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_504),
.B(n_170),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g622 ( 
.A(n_450),
.B(n_328),
.C(n_326),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_553),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_553),
.B(n_560),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_560),
.B(n_571),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_491),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_453),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_453),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_543),
.A2(n_429),
.B(n_428),
.C(n_426),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_566),
.B(n_427),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_471),
.B(n_388),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_551),
.B(n_427),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_483),
.B(n_328),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_471),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_504),
.B(n_572),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_440),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_473),
.B(n_388),
.Y(n_637)
);

INVx8_ASAP7_75t_L g638 ( 
.A(n_441),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_440),
.B(n_330),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_441),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_473),
.B(n_388),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_480),
.B(n_426),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_446),
.B(n_171),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_542),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_477),
.B(n_403),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_542),
.Y(n_646)
);

NOR3xp33_ASAP7_75t_L g647 ( 
.A(n_490),
.B(n_468),
.C(n_485),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_482),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_477),
.B(n_403),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_481),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_493),
.B(n_171),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_481),
.Y(n_652)
);

AND2x6_ASAP7_75t_L g653 ( 
.A(n_480),
.B(n_391),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_564),
.A2(n_269),
.B1(n_172),
.B2(n_169),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_543),
.A2(n_344),
.B1(n_351),
.B2(n_366),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_492),
.B(n_403),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_551),
.B(n_427),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_470),
.B(n_270),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_482),
.B(n_465),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_489),
.B(n_270),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_554),
.B(n_274),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_568),
.B(n_428),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_501),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_487),
.B(n_367),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_544),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_505),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_505),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_551),
.B(n_427),
.Y(n_668)
);

NAND3xp33_ASAP7_75t_SL g669 ( 
.A(n_564),
.B(n_271),
.C(n_296),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_546),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_511),
.B(n_405),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_511),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_488),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_551),
.B(n_265),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_551),
.B(n_265),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_546),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_577),
.B(n_268),
.C(n_257),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_512),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_475),
.B(n_279),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_462),
.B(n_367),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_454),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_570),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_520),
.B(n_521),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_520),
.B(n_405),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_570),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_456),
.B(n_279),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_435),
.B(n_282),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_521),
.B(n_405),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_SL g689 ( 
.A(n_484),
.B(n_172),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_522),
.B(n_391),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_551),
.B(n_265),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_454),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_570),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_538),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_578),
.B(n_429),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_562),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_557),
.B(n_282),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_522),
.B(n_424),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_523),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_523),
.B(n_424),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_526),
.B(n_424),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_526),
.B(n_527),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_472),
.B(n_338),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_527),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_518),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_448),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_530),
.B(n_424),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_576),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_L g709 ( 
.A(n_570),
.B(n_424),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_558),
.B(n_284),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_576),
.B(n_424),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_455),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_569),
.B(n_424),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_455),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_484),
.B(n_261),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_574),
.B(n_338),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_569),
.B(n_578),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_569),
.B(n_429),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_532),
.B(n_420),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_532),
.B(n_420),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_541),
.B(n_206),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_508),
.B(n_286),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_474),
.A2(n_212),
.B1(n_211),
.B2(n_213),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_517),
.A2(n_214),
.B1(n_217),
.B2(n_218),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_507),
.B(n_287),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_457),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_532),
.B(n_420),
.Y(n_727)
);

NOR2xp67_ASAP7_75t_L g728 ( 
.A(n_574),
.B(n_224),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_555),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_457),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_537),
.B(n_420),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_549),
.A2(n_235),
.B1(n_240),
.B2(n_243),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_518),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_540),
.B(n_289),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_555),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_459),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_556),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_537),
.B(n_420),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_591),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_640),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_599),
.A2(n_607),
.B1(n_581),
.B2(n_609),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_593),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_696),
.B(n_548),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_603),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_696),
.B(n_579),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_611),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_636),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_612),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_618),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_623),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_636),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_635),
.B(n_648),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_604),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_683),
.B(n_534),
.Y(n_754)
);

AND2x6_ASAP7_75t_L g755 ( 
.A(n_716),
.B(n_707),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_635),
.B(n_479),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_594),
.B(n_613),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_588),
.B(n_479),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_642),
.B(n_339),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_590),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_702),
.B(n_534),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_596),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_642),
.B(n_339),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_592),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_634),
.B(n_539),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_682),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_708),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_662),
.B(n_340),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_663),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_666),
.B(n_539),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_667),
.B(n_496),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_672),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_664),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_662),
.B(n_340),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_678),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_601),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_699),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_704),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_605),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_633),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_606),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_597),
.B(n_537),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_682),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_R g784 ( 
.A(n_639),
.B(n_289),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_582),
.B(n_341),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_607),
.A2(n_549),
.B1(n_288),
.B2(n_296),
.Y(n_786)
);

XNOR2x2_ASAP7_75t_L g787 ( 
.A(n_669),
.B(n_549),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_624),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_588),
.B(n_479),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_633),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_659),
.A2(n_283),
.B1(n_299),
.B2(n_298),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_615),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_625),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_682),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_584),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_694),
.B(n_341),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_690),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_716),
.B(n_547),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_580),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_650),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_627),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_628),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_600),
.A2(n_533),
.B(n_552),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_585),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_590),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_619),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_644),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_586),
.A2(n_533),
.B(n_552),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_703),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_629),
.B(n_547),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_583),
.Y(n_811)
);

CKINVDCx14_ASAP7_75t_R g812 ( 
.A(n_652),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_622),
.A2(n_514),
.B(n_486),
.C(n_495),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_661),
.B(n_647),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_589),
.B(n_459),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_589),
.B(n_464),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_633),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_595),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_647),
.B(n_541),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_646),
.Y(n_820)
);

BUFx8_ASAP7_75t_L g821 ( 
.A(n_673),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_589),
.B(n_464),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_621),
.B(n_479),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_622),
.A2(n_486),
.B(n_466),
.C(n_467),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_598),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_586),
.A2(n_514),
.B(n_506),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_705),
.Y(n_827)
);

NOR2x2_ASAP7_75t_L g828 ( 
.A(n_654),
.B(n_261),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_638),
.B(n_343),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_619),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_638),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_638),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_631),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_637),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_589),
.A2(n_533),
.B1(n_552),
.B2(n_525),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_641),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_680),
.B(n_541),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_589),
.B(n_466),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_665),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_670),
.Y(n_840)
);

AO22x1_ASAP7_75t_L g841 ( 
.A1(n_660),
.A2(n_288),
.B1(n_269),
.B2(n_271),
.Y(n_841)
);

AND3x2_ASAP7_75t_SL g842 ( 
.A(n_654),
.B(n_278),
.C(n_281),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_733),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_706),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_626),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_655),
.B(n_347),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_722),
.A2(n_447),
.B1(n_502),
.B2(n_525),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_626),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_621),
.B(n_467),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_677),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_643),
.B(n_347),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_643),
.B(n_349),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_697),
.A2(n_447),
.B1(n_565),
.B2(n_567),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_689),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_645),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_587),
.A2(n_575),
.B(n_573),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_660),
.A2(n_575),
.B1(n_573),
.B2(n_567),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_682),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_728),
.B(n_349),
.Y(n_859)
);

CKINVDCx11_ASAP7_75t_R g860 ( 
.A(n_715),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_649),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_630),
.B(n_350),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_679),
.B(n_565),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_697),
.A2(n_563),
.B1(n_556),
.B2(n_559),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_676),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_681),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_653),
.B(n_495),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_630),
.B(n_350),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_653),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_692),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_712),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_587),
.B(n_353),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_653),
.B(n_499),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_714),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_602),
.A2(n_515),
.B(n_535),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_R g876 ( 
.A(n_687),
.B(n_476),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_653),
.A2(n_515),
.B1(n_535),
.B2(n_509),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_653),
.B(n_658),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_651),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_687),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_726),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_710),
.B(n_561),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_679),
.B(n_195),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_656),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_730),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_658),
.B(n_503),
.Y(n_886)
);

OAI21xp33_ASAP7_75t_L g887 ( 
.A1(n_710),
.A2(n_299),
.B(n_278),
.Y(n_887)
);

AND2x6_ASAP7_75t_SL g888 ( 
.A(n_734),
.B(n_353),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_686),
.B(n_199),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_671),
.Y(n_890)
);

AND2x6_ASAP7_75t_L g891 ( 
.A(n_732),
.B(n_561),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_736),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_723),
.B(n_561),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_725),
.B(n_354),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_717),
.B(n_503),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_718),
.B(n_506),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_729),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_685),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_721),
.A2(n_264),
.B1(n_249),
.B2(n_254),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_608),
.A2(n_617),
.B(n_610),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_735),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_685),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_684),
.B(n_513),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_688),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_721),
.A2(n_258),
.B1(n_245),
.B2(n_247),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_685),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_614),
.B(n_513),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_620),
.A2(n_516),
.B(n_528),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_745),
.A2(n_616),
.B1(n_701),
.B2(n_698),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_759),
.B(n_695),
.Y(n_910)
);

AO32x1_ASAP7_75t_L g911 ( 
.A1(n_741),
.A2(n_737),
.A3(n_365),
.B1(n_354),
.B2(n_359),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_893),
.A2(n_693),
.B(n_713),
.Y(n_912)
);

INVxp67_ASAP7_75t_SL g913 ( 
.A(n_760),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_766),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_747),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_742),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_766),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_741),
.A2(n_734),
.B1(n_616),
.B2(n_700),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_883),
.A2(n_711),
.B(n_724),
.C(n_727),
.Y(n_919)
);

OAI21xp33_ASAP7_75t_L g920 ( 
.A1(n_887),
.A2(n_292),
.B(n_298),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_803),
.A2(n_693),
.B(n_709),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_745),
.A2(n_693),
.B1(n_731),
.B2(n_720),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_788),
.B(n_516),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_793),
.B(n_719),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_751),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_811),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_752),
.B(n_738),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_809),
.B(n_359),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_750),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_809),
.A2(n_814),
.B1(n_804),
.B2(n_799),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_818),
.B(n_825),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_759),
.B(n_632),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_827),
.B(n_657),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_763),
.B(n_668),
.Y(n_934)
);

OAI22x1_ASAP7_75t_L g935 ( 
.A1(n_879),
.A2(n_292),
.B1(n_291),
.B2(n_281),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_764),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_749),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_844),
.A2(n_675),
.B1(n_674),
.B2(n_691),
.Y(n_938)
);

AOI21x1_ASAP7_75t_L g939 ( 
.A1(n_882),
.A2(n_476),
.B(n_497),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_743),
.A2(n_291),
.B1(n_203),
.B2(n_204),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_766),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_767),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_783),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_889),
.A2(n_691),
.B(n_674),
.C(n_267),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_743),
.A2(n_761),
.B1(n_754),
.B2(n_872),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_769),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_851),
.B(n_528),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_SL g948 ( 
.A1(n_819),
.A2(n_364),
.B(n_319),
.C(n_324),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_773),
.B(n_528),
.Y(n_949)
);

NOR3xp33_ASAP7_75t_SL g950 ( 
.A(n_784),
.B(n_364),
.C(n_321),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_800),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_783),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_852),
.B(n_528),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_772),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_763),
.B(n_319),
.Y(n_955)
);

BUFx12f_ASAP7_75t_L g956 ( 
.A(n_821),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_775),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_739),
.Y(n_958)
);

NOR2x1_ASAP7_75t_L g959 ( 
.A(n_832),
.B(n_528),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_797),
.B(n_510),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_821),
.Y(n_961)
);

AOI21x1_ASAP7_75t_L g962 ( 
.A1(n_771),
.A2(n_324),
.B(n_322),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_812),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_758),
.B(n_510),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_SL g965 ( 
.A1(n_878),
.A2(n_133),
.B(n_126),
.C(n_119),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_810),
.A2(n_420),
.B(n_469),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_779),
.B(n_796),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_789),
.B(n_756),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_810),
.A2(n_420),
.B(n_469),
.Y(n_969)
);

NOR3xp33_ASAP7_75t_L g970 ( 
.A(n_841),
.B(n_1),
.C(n_2),
.Y(n_970)
);

AND2x2_ASAP7_75t_SL g971 ( 
.A(n_842),
.B(n_4),
.Y(n_971)
);

O2A1O1Ixp5_ASAP7_75t_L g972 ( 
.A1(n_823),
.A2(n_510),
.B(n_469),
.C(n_461),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_777),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_754),
.A2(n_510),
.B1(n_469),
.B2(n_461),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_863),
.B(n_461),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_850),
.B(n_461),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_786),
.A2(n_6),
.B(n_8),
.C(n_14),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_778),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_817),
.B(n_461),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_753),
.B(n_437),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_794),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_862),
.B(n_437),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_831),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_796),
.B(n_6),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_768),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_856),
.A2(n_437),
.B(n_420),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_862),
.B(n_437),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_744),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_805),
.A2(n_437),
.B(n_420),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_746),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_748),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_868),
.B(n_420),
.Y(n_992)
);

AOI21xp33_ASAP7_75t_L g993 ( 
.A1(n_846),
.A2(n_15),
.B(n_16),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_761),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_859),
.B(n_117),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_868),
.A2(n_19),
.B1(n_20),
.B2(n_23),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_785),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_880),
.B(n_23),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_805),
.A2(n_47),
.B(n_102),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_780),
.B(n_25),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_849),
.B(n_48),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_859),
.B(n_107),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_790),
.B(n_26),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_849),
.B(n_28),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_833),
.B(n_51),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_886),
.A2(n_100),
.B(n_99),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_774),
.B(n_29),
.Y(n_1007)
);

INVxp67_ASAP7_75t_SL g1008 ( 
.A(n_794),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_786),
.A2(n_29),
.B(n_31),
.C(n_33),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_R g1010 ( 
.A(n_854),
.B(n_89),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_794),
.Y(n_1011)
);

OR2x6_ASAP7_75t_L g1012 ( 
.A(n_843),
.B(n_71),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_834),
.B(n_31),
.Y(n_1013)
);

OR2x6_ASAP7_75t_L g1014 ( 
.A(n_829),
.B(n_70),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_886),
.A2(n_53),
.B(n_55),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_808),
.A2(n_44),
.B(n_35),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_791),
.B(n_34),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_878),
.A2(n_35),
.B(n_38),
.C(n_39),
.Y(n_1018)
);

BUFx10_ASAP7_75t_L g1019 ( 
.A(n_888),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_872),
.A2(n_38),
.B1(n_44),
.B2(n_798),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_872),
.A2(n_798),
.B1(n_771),
.B2(n_765),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_757),
.A2(n_837),
.B(n_894),
.C(n_795),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_836),
.B(n_855),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_829),
.B(n_774),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_898),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_897),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_808),
.A2(n_848),
.B(n_782),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_829),
.B(n_861),
.Y(n_1028)
);

AO22x1_ASAP7_75t_L g1029 ( 
.A1(n_842),
.A2(n_891),
.B1(n_755),
.B2(n_869),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_876),
.B(n_898),
.Y(n_1030)
);

CKINVDCx10_ASAP7_75t_R g1031 ( 
.A(n_860),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_901),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_898),
.B(n_906),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_765),
.A2(n_770),
.B1(n_830),
.B2(n_806),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_L g1035 ( 
.A(n_899),
.B(n_905),
.C(n_822),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_906),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_866),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_782),
.A2(n_900),
.B(n_895),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_906),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_806),
.B(n_830),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_884),
.A2(n_904),
.B(n_890),
.C(n_900),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1023),
.B(n_755),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1022),
.A2(n_824),
.B(n_813),
.C(n_815),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_921),
.A2(n_908),
.B(n_875),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_931),
.B(n_927),
.Y(n_1045)
);

CKINVDCx6p67_ASAP7_75t_R g1046 ( 
.A(n_1031),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_918),
.A2(n_857),
.B1(n_845),
.B2(n_877),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_964),
.A2(n_896),
.B(n_895),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_1014),
.B(n_858),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_929),
.Y(n_1050)
);

AO31x2_ASAP7_75t_L g1051 ( 
.A1(n_1021),
.A2(n_838),
.A3(n_816),
.B(n_867),
.Y(n_1051)
);

O2A1O1Ixp5_ASAP7_75t_L g1052 ( 
.A1(n_1029),
.A2(n_826),
.B(n_875),
.C(n_903),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_915),
.Y(n_1053)
);

AOI221x1_ASAP7_75t_L g1054 ( 
.A1(n_1016),
.A2(n_826),
.B1(n_787),
.B2(n_903),
.C(n_907),
.Y(n_1054)
);

OA21x2_ASAP7_75t_L g1055 ( 
.A1(n_972),
.A2(n_864),
.B(n_907),
.Y(n_1055)
);

NAND3x1_ASAP7_75t_L g1056 ( 
.A(n_1017),
.B(n_828),
.C(n_902),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_997),
.B(n_762),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_930),
.A2(n_776),
.B(n_781),
.C(n_792),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_SL g1059 ( 
.A1(n_1005),
.A2(n_873),
.B(n_867),
.C(n_835),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_926),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_SL g1061 ( 
.A1(n_945),
.A2(n_853),
.B(n_847),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_930),
.B(n_807),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_955),
.B(n_984),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_936),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_919),
.A2(n_891),
.B(n_865),
.Y(n_1065)
);

AO31x2_ASAP7_75t_L g1066 ( 
.A1(n_1021),
.A2(n_874),
.A3(n_892),
.B(n_885),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_983),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_924),
.B(n_801),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_951),
.B(n_820),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_942),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_925),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_1035),
.A2(n_802),
.B(n_839),
.C(n_840),
.Y(n_1072)
);

AND2x6_ASAP7_75t_L g1073 ( 
.A(n_932),
.B(n_902),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_946),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_947),
.B(n_870),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_SL g1076 ( 
.A(n_920),
.B(n_891),
.C(n_871),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_SL g1077 ( 
.A(n_971),
.B(n_891),
.Y(n_1077)
);

AOI211x1_ASAP7_75t_L g1078 ( 
.A1(n_993),
.A2(n_881),
.B(n_1020),
.C(n_994),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_SL g1079 ( 
.A1(n_996),
.A2(n_993),
.B(n_1009),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_917),
.Y(n_1080)
);

AO31x2_ASAP7_75t_L g1081 ( 
.A1(n_974),
.A2(n_1034),
.A3(n_1001),
.B(n_909),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1001),
.A2(n_909),
.B(n_966),
.Y(n_1082)
);

OA21x2_ASAP7_75t_L g1083 ( 
.A1(n_966),
.A2(n_969),
.B(n_1004),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_988),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_963),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_954),
.A2(n_957),
.B1(n_973),
.B2(n_978),
.Y(n_1086)
);

NAND2xp33_ASAP7_75t_L g1087 ( 
.A(n_1013),
.B(n_990),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1028),
.B(n_910),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_969),
.A2(n_922),
.B(n_1034),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_953),
.B(n_923),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_974),
.A2(n_989),
.B(n_922),
.Y(n_1091)
);

AO21x2_ASAP7_75t_L g1092 ( 
.A1(n_976),
.A2(n_1005),
.B(n_1030),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_913),
.A2(n_960),
.B(n_987),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_951),
.B(n_950),
.Y(n_1094)
);

AO21x1_ASAP7_75t_L g1095 ( 
.A1(n_977),
.A2(n_1020),
.B(n_994),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_SL g1096 ( 
.A1(n_944),
.A2(n_982),
.B(n_1014),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_938),
.A2(n_1015),
.B(n_1006),
.Y(n_1097)
);

AOI221x1_ASAP7_75t_L g1098 ( 
.A1(n_970),
.A2(n_1018),
.B1(n_935),
.B2(n_1003),
.C(n_1000),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_914),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_999),
.A2(n_992),
.B(n_1040),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_910),
.A2(n_932),
.B(n_934),
.C(n_937),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_995),
.A2(n_1002),
.B(n_980),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_985),
.B(n_934),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_991),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_933),
.B(n_1026),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_949),
.A2(n_959),
.B(n_1033),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_916),
.A2(n_1032),
.B(n_1037),
.Y(n_1107)
);

AOI21x1_ASAP7_75t_L g1108 ( 
.A1(n_979),
.A2(n_928),
.B(n_933),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1008),
.A2(n_965),
.B(n_911),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_948),
.A2(n_940),
.B(n_979),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_998),
.B(n_1007),
.Y(n_1111)
);

OA21x2_ASAP7_75t_L g1112 ( 
.A1(n_911),
.A2(n_1024),
.B(n_940),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_911),
.A2(n_933),
.B(n_1014),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_941),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_952),
.B(n_1036),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_943),
.A2(n_1025),
.B(n_981),
.Y(n_1116)
);

OAI21xp33_ASAP7_75t_L g1117 ( 
.A1(n_1010),
.A2(n_1012),
.B(n_961),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1012),
.A2(n_914),
.B(n_1011),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1012),
.B(n_1019),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_SL g1120 ( 
.A1(n_914),
.A2(n_1011),
.B(n_1039),
.C(n_1019),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_956),
.Y(n_1121)
);

NAND2xp33_ASAP7_75t_L g1122 ( 
.A(n_968),
.B(n_640),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_931),
.B(n_745),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_915),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_921),
.A2(n_912),
.B(n_986),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_931),
.B(n_745),
.Y(n_1126)
);

NOR2xp67_ASAP7_75t_L g1127 ( 
.A(n_983),
.B(n_740),
.Y(n_1127)
);

NAND3x1_ASAP7_75t_L g1128 ( 
.A(n_1017),
.B(n_970),
.C(n_883),
.Y(n_1128)
);

AO32x2_ASAP7_75t_L g1129 ( 
.A1(n_1021),
.A2(n_741),
.A3(n_945),
.B1(n_994),
.B2(n_930),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_967),
.B(n_635),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_1021),
.A2(n_741),
.A3(n_945),
.B(n_1038),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_997),
.B(n_967),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_921),
.A2(n_912),
.B(n_986),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_921),
.A2(n_912),
.B(n_986),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_931),
.B(n_504),
.Y(n_1135)
);

NAND3x1_ASAP7_75t_L g1136 ( 
.A(n_1017),
.B(n_970),
.C(n_883),
.Y(n_1136)
);

AOI21x1_ASAP7_75t_L g1137 ( 
.A1(n_962),
.A2(n_939),
.B(n_975),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1031),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1017),
.A2(n_883),
.B(n_581),
.C(n_463),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_921),
.A2(n_912),
.B(n_986),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_968),
.A2(n_741),
.B(n_1041),
.Y(n_1141)
);

AO21x1_ASAP7_75t_L g1142 ( 
.A1(n_968),
.A2(n_741),
.B(n_814),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_921),
.A2(n_912),
.B(n_986),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_968),
.B(n_745),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_914),
.Y(n_1145)
);

AOI21x1_ASAP7_75t_L g1146 ( 
.A1(n_962),
.A2(n_939),
.B(n_975),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_967),
.B(n_635),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1038),
.A2(n_968),
.B(n_975),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_926),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_968),
.B(n_745),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_958),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_968),
.A2(n_741),
.B(n_1041),
.Y(n_1152)
);

AOI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_968),
.A2(n_741),
.B(n_883),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_929),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_968),
.B(n_745),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_968),
.B(n_745),
.Y(n_1156)
);

OA21x2_ASAP7_75t_L g1157 ( 
.A1(n_972),
.A2(n_1038),
.B(n_1027),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_931),
.B(n_308),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_968),
.B(n_745),
.Y(n_1159)
);

CKINVDCx11_ASAP7_75t_R g1160 ( 
.A(n_956),
.Y(n_1160)
);

AOI211x1_ASAP7_75t_L g1161 ( 
.A1(n_993),
.A2(n_654),
.B(n_669),
.C(n_930),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1139),
.B(n_1144),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_1105),
.B(n_1108),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1044),
.A2(n_1133),
.B(n_1125),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1130),
.B(n_1147),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1134),
.A2(n_1143),
.B(n_1140),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_SL g1167 ( 
.A(n_1138),
.B(n_1067),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_1098),
.B(n_1153),
.C(n_1161),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1153),
.A2(n_1095),
.B1(n_1077),
.B2(n_1152),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1103),
.B(n_1132),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1141),
.A2(n_1152),
.B(n_1082),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_1062),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1050),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1144),
.B(n_1150),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_SL g1175 ( 
.A1(n_1102),
.A2(n_1113),
.B(n_1110),
.Y(n_1175)
);

AND2x4_ASAP7_75t_SL g1176 ( 
.A(n_1053),
.B(n_1124),
.Y(n_1176)
);

INVx8_ASAP7_75t_L g1177 ( 
.A(n_1073),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1063),
.B(n_1111),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1141),
.A2(n_1077),
.B(n_1079),
.C(n_1045),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1045),
.A2(n_1150),
.B1(n_1155),
.B2(n_1159),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1079),
.A2(n_1156),
.B(n_1155),
.C(n_1159),
.Y(n_1181)
);

AOI222xp33_ASAP7_75t_L g1182 ( 
.A1(n_1158),
.A2(n_1122),
.B1(n_1126),
.B2(n_1123),
.C1(n_1156),
.C2(n_1094),
.Y(n_1182)
);

OR2x6_ASAP7_75t_L g1183 ( 
.A(n_1049),
.B(n_1096),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_1135),
.B(n_1088),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1084),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_SL g1186 ( 
.A(n_1046),
.B(n_1127),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1151),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_SL g1188 ( 
.A1(n_1110),
.A2(n_1042),
.B(n_1100),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1148),
.A2(n_1097),
.B(n_1065),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1137),
.A2(n_1146),
.B(n_1048),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1128),
.A2(n_1136),
.B1(n_1117),
.B2(n_1056),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1052),
.A2(n_1100),
.B(n_1093),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1071),
.B(n_1069),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1090),
.B(n_1068),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1090),
.B(n_1068),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_1105),
.B(n_1080),
.Y(n_1196)
);

OA21x2_ASAP7_75t_L g1197 ( 
.A1(n_1089),
.A2(n_1043),
.B(n_1072),
.Y(n_1197)
);

NAND2x1p5_ASAP7_75t_L g1198 ( 
.A(n_1080),
.B(n_1116),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1049),
.B(n_1101),
.Y(n_1199)
);

INVx2_ASAP7_75t_SL g1200 ( 
.A(n_1060),
.Y(n_1200)
);

AOI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1055),
.A2(n_1157),
.B(n_1089),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1157),
.A2(n_1106),
.B(n_1058),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1149),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1087),
.A2(n_1112),
.B1(n_1047),
.B2(n_1049),
.Y(n_1204)
);

OAI221xp5_ASAP7_75t_L g1205 ( 
.A1(n_1061),
.A2(n_1086),
.B1(n_1076),
.B2(n_1104),
.C(n_1154),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1066),
.Y(n_1206)
);

AOI221xp5_ASAP7_75t_L g1207 ( 
.A1(n_1078),
.A2(n_1086),
.B1(n_1047),
.B2(n_1074),
.C(n_1070),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1066),
.Y(n_1208)
);

AOI222xp33_ASAP7_75t_L g1209 ( 
.A1(n_1119),
.A2(n_1121),
.B1(n_1064),
.B2(n_1057),
.C1(n_1160),
.C2(n_1075),
.Y(n_1209)
);

AO21x2_ASAP7_75t_L g1210 ( 
.A1(n_1059),
.A2(n_1092),
.B(n_1075),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1107),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1057),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1083),
.A2(n_1112),
.B(n_1118),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1114),
.B(n_1115),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1099),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1099),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1066),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1131),
.A2(n_1129),
.B(n_1081),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1129),
.A2(n_1131),
.B(n_1081),
.C(n_1051),
.Y(n_1219)
);

BUFx4_ASAP7_75t_SL g1220 ( 
.A(n_1085),
.Y(n_1220)
);

INVx6_ASAP7_75t_L g1221 ( 
.A(n_1145),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1129),
.A2(n_1051),
.B(n_1120),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1073),
.B(n_1139),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1073),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1128),
.A2(n_883),
.B1(n_1136),
.B2(n_311),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1064),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1064),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1044),
.A2(n_1133),
.B(n_1125),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1050),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1139),
.A2(n_1153),
.B(n_968),
.C(n_1152),
.Y(n_1230)
);

INVxp33_ASAP7_75t_SL g1231 ( 
.A(n_1067),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1044),
.A2(n_1133),
.B(n_1125),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1064),
.Y(n_1233)
);

INVx5_ASAP7_75t_L g1234 ( 
.A(n_1073),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1139),
.B(n_883),
.C(n_581),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_SL g1236 ( 
.A1(n_1153),
.A2(n_1139),
.B(n_814),
.C(n_968),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_SL g1237 ( 
.A1(n_1139),
.A2(n_1045),
.B(n_968),
.Y(n_1237)
);

OA21x2_ASAP7_75t_L g1238 ( 
.A1(n_1054),
.A2(n_1091),
.B(n_1044),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1067),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1139),
.B(n_581),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1139),
.A2(n_1153),
.B(n_1152),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1044),
.A2(n_1133),
.B(n_1125),
.Y(n_1242)
);

OR2x6_ASAP7_75t_L g1243 ( 
.A(n_1049),
.B(n_1096),
.Y(n_1243)
);

INVxp67_ASAP7_75t_SL g1244 ( 
.A(n_1062),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1050),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1153),
.A2(n_971),
.B1(n_1095),
.B2(n_1017),
.Y(n_1246)
);

AO21x2_ASAP7_75t_L g1247 ( 
.A1(n_1141),
.A2(n_1152),
.B(n_1153),
.Y(n_1247)
);

AO21x2_ASAP7_75t_L g1248 ( 
.A1(n_1141),
.A2(n_1152),
.B(n_1153),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1135),
.B(n_1088),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1044),
.A2(n_1133),
.B(n_1125),
.Y(n_1250)
);

CKINVDCx11_ASAP7_75t_R g1251 ( 
.A(n_1046),
.Y(n_1251)
);

INVx5_ASAP7_75t_L g1252 ( 
.A(n_1073),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1073),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1144),
.B(n_1150),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1099),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1144),
.B(n_1150),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1050),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1142),
.A2(n_1054),
.A3(n_1095),
.B(n_1109),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1064),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1142),
.A2(n_1054),
.A3(n_1095),
.B(n_1109),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1044),
.A2(n_1133),
.B(n_1125),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1139),
.B(n_1153),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1046),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1044),
.A2(n_1133),
.B(n_1125),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1099),
.Y(n_1265)
);

OAI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1077),
.A2(n_968),
.B1(n_1045),
.B2(n_1144),
.Y(n_1266)
);

CKINVDCx11_ASAP7_75t_R g1267 ( 
.A(n_1046),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1060),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1173),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1162),
.B(n_1181),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1268),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1240),
.A2(n_1235),
.B(n_1262),
.C(n_1230),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1215),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1162),
.B(n_1181),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1240),
.A2(n_1262),
.B(n_1230),
.C(n_1236),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1178),
.B(n_1165),
.Y(n_1276)
);

NAND3xp33_ASAP7_75t_L g1277 ( 
.A(n_1246),
.B(n_1182),
.C(n_1225),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_SL g1278 ( 
.A1(n_1179),
.A2(n_1172),
.B(n_1244),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1184),
.B(n_1249),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1215),
.Y(n_1280)
);

NOR2xp67_ASAP7_75t_L g1281 ( 
.A(n_1239),
.B(n_1193),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1213),
.A2(n_1202),
.B(n_1189),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1191),
.A2(n_1246),
.B1(n_1223),
.B2(n_1169),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1241),
.A2(n_1223),
.B(n_1171),
.C(n_1179),
.Y(n_1284)
);

NOR2xp67_ASAP7_75t_L g1285 ( 
.A(n_1193),
.B(n_1200),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_1251),
.Y(n_1286)
);

NOR2xp67_ASAP7_75t_L g1287 ( 
.A(n_1185),
.B(n_1187),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1215),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1214),
.B(n_1212),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1176),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1236),
.A2(n_1241),
.B(n_1266),
.C(n_1168),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1231),
.B(n_1259),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1180),
.A2(n_1169),
.B1(n_1256),
.B2(n_1254),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1180),
.B(n_1174),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1229),
.B(n_1245),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1203),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1257),
.B(n_1194),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1194),
.B(n_1195),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1195),
.A2(n_1237),
.B1(n_1197),
.B2(n_1234),
.Y(n_1299)
);

O2A1O1Ixp5_ASAP7_75t_L g1300 ( 
.A1(n_1222),
.A2(n_1218),
.B(n_1219),
.C(n_1201),
.Y(n_1300)
);

AOI21x1_ASAP7_75t_SL g1301 ( 
.A1(n_1206),
.A2(n_1208),
.B(n_1217),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1183),
.A2(n_1243),
.B(n_1199),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1205),
.A2(n_1209),
.B(n_1175),
.C(n_1188),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1205),
.A2(n_1247),
.B(n_1248),
.C(n_1163),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1207),
.B(n_1248),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1197),
.A2(n_1252),
.B1(n_1234),
.B2(n_1207),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1183),
.A2(n_1243),
.B(n_1199),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1226),
.B(n_1233),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1227),
.B(n_1196),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1163),
.B(n_1216),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1199),
.A2(n_1219),
.B(n_1183),
.C(n_1243),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1234),
.A2(n_1252),
.B1(n_1204),
.B2(n_1218),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1204),
.A2(n_1253),
.B(n_1186),
.C(n_1211),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1167),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1252),
.A2(n_1210),
.B(n_1177),
.Y(n_1315)
);

INVxp67_ASAP7_75t_L g1316 ( 
.A(n_1255),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1258),
.B(n_1260),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1177),
.A2(n_1221),
.B1(n_1265),
.B2(n_1255),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1164),
.A2(n_1242),
.B(n_1264),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1198),
.A2(n_1238),
.B(n_1263),
.C(n_1220),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1228),
.A2(n_1261),
.B(n_1250),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1255),
.B(n_1221),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1232),
.B(n_1166),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1238),
.B(n_1198),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1221),
.A2(n_1246),
.B1(n_971),
.B2(n_968),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1220),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1267),
.B(n_308),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1162),
.B(n_1181),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1224),
.B(n_1170),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1184),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1213),
.A2(n_1190),
.B(n_1192),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1162),
.B(n_1180),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1162),
.B(n_1180),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1203),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1178),
.B(n_1165),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1240),
.A2(n_1139),
.B(n_968),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1178),
.B(n_1165),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1240),
.A2(n_1139),
.B(n_1235),
.C(n_883),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_SL g1339 ( 
.A1(n_1240),
.A2(n_1139),
.B(n_968),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1162),
.B(n_1181),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1178),
.B(n_1165),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1246),
.A2(n_971),
.B1(n_968),
.B2(n_1180),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1213),
.A2(n_1190),
.B(n_1192),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1162),
.B(n_1181),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1323),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1269),
.Y(n_1346)
);

AO21x1_ASAP7_75t_SL g1347 ( 
.A1(n_1317),
.A2(n_1270),
.B(n_1340),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1324),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1277),
.B(n_1332),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1270),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1300),
.B(n_1282),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1323),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1274),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1274),
.B(n_1328),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1305),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1305),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1328),
.B(n_1340),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1284),
.B(n_1331),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1343),
.B(n_1312),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1319),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1295),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1315),
.A2(n_1301),
.B(n_1307),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1312),
.B(n_1344),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1344),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1333),
.B(n_1294),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1283),
.A2(n_1325),
.B1(n_1342),
.B2(n_1293),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1297),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1279),
.B(n_1304),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1321),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1330),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1321),
.Y(n_1371)
);

BUFx12f_ASAP7_75t_L g1372 ( 
.A(n_1326),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1299),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1299),
.Y(n_1374)
);

INVx5_ASAP7_75t_L g1375 ( 
.A(n_1302),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1278),
.B(n_1289),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1306),
.B(n_1275),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1294),
.B(n_1293),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1338),
.A2(n_1339),
.B(n_1336),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1272),
.B(n_1342),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1291),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1311),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1310),
.Y(n_1383)
);

AO21x2_ASAP7_75t_L g1384 ( 
.A1(n_1306),
.A2(n_1325),
.B(n_1303),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1276),
.B(n_1341),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1335),
.B(n_1337),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1298),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1346),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1348),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1360),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1355),
.B(n_1309),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1358),
.B(n_1320),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1358),
.B(n_1351),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1349),
.A2(n_1314),
.B1(n_1281),
.B2(n_1329),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1360),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1347),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1358),
.B(n_1313),
.Y(n_1397)
);

CKINVDCx14_ASAP7_75t_R g1398 ( 
.A(n_1372),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1351),
.B(n_1287),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1351),
.B(n_1334),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1350),
.Y(n_1401)
);

NOR2x1_ASAP7_75t_L g1402 ( 
.A(n_1379),
.B(n_1285),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1369),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1359),
.B(n_1308),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1350),
.B(n_1316),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1355),
.B(n_1322),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1369),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1353),
.B(n_1290),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1371),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1345),
.B(n_1352),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1353),
.B(n_1296),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1371),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1347),
.B(n_1288),
.Y(n_1413)
);

AOI221xp5_ASAP7_75t_L g1414 ( 
.A1(n_1397),
.A2(n_1349),
.B1(n_1381),
.B2(n_1380),
.C(n_1354),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1393),
.B(n_1368),
.Y(n_1415)
);

AOI33xp33_ASAP7_75t_L g1416 ( 
.A1(n_1392),
.A2(n_1381),
.A3(n_1366),
.B1(n_1377),
.B2(n_1368),
.B3(n_1363),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1405),
.B(n_1364),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1401),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1401),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1394),
.A2(n_1366),
.B1(n_1380),
.B2(n_1381),
.Y(n_1420)
);

AOI221xp5_ASAP7_75t_L g1421 ( 
.A1(n_1397),
.A2(n_1354),
.B1(n_1365),
.B2(n_1368),
.C(n_1370),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1405),
.B(n_1364),
.Y(n_1422)
);

OAI321xp33_ASAP7_75t_L g1423 ( 
.A1(n_1392),
.A2(n_1377),
.A3(n_1382),
.B1(n_1374),
.B2(n_1373),
.C(n_1378),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1410),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1402),
.A2(n_1379),
.B(n_1384),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1389),
.B(n_1348),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1393),
.B(n_1348),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1409),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1410),
.B(n_1352),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_1389),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1392),
.A2(n_1379),
.B1(n_1384),
.B2(n_1377),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1388),
.Y(n_1432)
);

NAND3xp33_ASAP7_75t_L g1433 ( 
.A(n_1402),
.B(n_1357),
.C(n_1378),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1388),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1393),
.B(n_1347),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1404),
.B(n_1364),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1411),
.Y(n_1437)
);

AOI33xp33_ASAP7_75t_L g1438 ( 
.A1(n_1392),
.A2(n_1363),
.A3(n_1356),
.B1(n_1387),
.B2(n_1373),
.B3(n_1374),
.Y(n_1438)
);

INVx5_ASAP7_75t_L g1439 ( 
.A(n_1396),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1397),
.A2(n_1379),
.B1(n_1384),
.B2(n_1382),
.Y(n_1440)
);

BUFx2_ASAP7_75t_SL g1441 ( 
.A(n_1413),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1397),
.A2(n_1384),
.B1(n_1382),
.B2(n_1364),
.Y(n_1442)
);

AOI221xp5_ASAP7_75t_L g1443 ( 
.A1(n_1408),
.A2(n_1365),
.B1(n_1370),
.B2(n_1357),
.C(n_1363),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1388),
.Y(n_1444)
);

OAI33xp33_ASAP7_75t_L g1445 ( 
.A1(n_1391),
.A2(n_1357),
.A3(n_1356),
.B1(n_1378),
.B2(n_1387),
.B3(n_1361),
.Y(n_1445)
);

AOI21xp33_ASAP7_75t_L g1446 ( 
.A1(n_1394),
.A2(n_1356),
.B(n_1376),
.Y(n_1446)
);

AOI31xp33_ASAP7_75t_L g1447 ( 
.A1(n_1398),
.A2(n_1376),
.A3(n_1327),
.B(n_1367),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1404),
.B(n_1383),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1409),
.Y(n_1449)
);

A2O1A1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1398),
.A2(n_1376),
.B(n_1362),
.C(n_1375),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1411),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1426),
.B(n_1393),
.Y(n_1452)
);

INVx4_ASAP7_75t_SL g1453 ( 
.A(n_1435),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1432),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1418),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1432),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1426),
.B(n_1436),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1434),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1434),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1439),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1444),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1419),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1428),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1433),
.A2(n_1390),
.B(n_1395),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1444),
.Y(n_1465)
);

AND2x6_ASAP7_75t_L g1466 ( 
.A(n_1435),
.B(n_1396),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1430),
.Y(n_1467)
);

AOI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1425),
.A2(n_1409),
.B(n_1412),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1448),
.B(n_1406),
.Y(n_1469)
);

INVx4_ASAP7_75t_SL g1470 ( 
.A(n_1429),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1433),
.A2(n_1390),
.B(n_1395),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1439),
.Y(n_1472)
);

OA21x2_ASAP7_75t_L g1473 ( 
.A1(n_1450),
.A2(n_1403),
.B(n_1407),
.Y(n_1473)
);

INVx4_ASAP7_75t_SL g1474 ( 
.A(n_1429),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1451),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1449),
.Y(n_1476)
);

NOR2x1p5_ASAP7_75t_L g1477 ( 
.A(n_1451),
.B(n_1372),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1414),
.A2(n_1403),
.B(n_1407),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1439),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1417),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1422),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1454),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1468),
.Y(n_1483)
);

NOR3xp33_ASAP7_75t_L g1484 ( 
.A(n_1460),
.B(n_1420),
.C(n_1447),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1460),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1475),
.B(n_1286),
.Y(n_1486)
);

XOR2xp5_ASAP7_75t_L g1487 ( 
.A(n_1462),
.B(n_1271),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1453),
.B(n_1439),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_1479),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1455),
.B(n_1421),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1479),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1481),
.B(n_1416),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1457),
.B(n_1415),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1456),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1480),
.B(n_1443),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1453),
.B(n_1415),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1453),
.B(n_1441),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1458),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1459),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1461),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1453),
.B(n_1441),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1470),
.B(n_1429),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1472),
.Y(n_1503)
);

OAI31xp33_ASAP7_75t_L g1504 ( 
.A1(n_1477),
.A2(n_1431),
.A3(n_1440),
.B(n_1442),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1467),
.B(n_1438),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1457),
.B(n_1437),
.Y(n_1506)
);

AND2x4_ASAP7_75t_SL g1507 ( 
.A(n_1472),
.B(n_1396),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1469),
.B(n_1372),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1470),
.B(n_1424),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1465),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1452),
.B(n_1406),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1470),
.B(n_1439),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1474),
.B(n_1427),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1466),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1474),
.B(n_1427),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1474),
.B(n_1466),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1474),
.B(n_1400),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1466),
.B(n_1400),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1463),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1489),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1482),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1488),
.B(n_1478),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1485),
.Y(n_1523)
);

AND2x4_ASAP7_75t_SL g1524 ( 
.A(n_1488),
.B(n_1396),
.Y(n_1524)
);

OAI21xp33_ASAP7_75t_L g1525 ( 
.A1(n_1490),
.A2(n_1446),
.B(n_1404),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1492),
.A2(n_1478),
.B(n_1423),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1482),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1485),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1493),
.B(n_1478),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1494),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1484),
.Y(n_1531)
);

NOR2x1_ASAP7_75t_L g1532 ( 
.A(n_1503),
.B(n_1464),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1505),
.B(n_1385),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1489),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1488),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1487),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1503),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1516),
.B(n_1466),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1503),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1494),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1495),
.B(n_1385),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1491),
.B(n_1385),
.Y(n_1542)
);

NAND3xp33_ASAP7_75t_L g1543 ( 
.A(n_1504),
.B(n_1473),
.C(n_1471),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1516),
.B(n_1466),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1508),
.B(n_1386),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1507),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1493),
.B(n_1463),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1506),
.B(n_1386),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1498),
.Y(n_1549)
);

OAI21xp33_ASAP7_75t_L g1550 ( 
.A1(n_1506),
.A2(n_1399),
.B(n_1391),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1496),
.B(n_1466),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1498),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1511),
.B(n_1476),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1499),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1551),
.B(n_1497),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1521),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1521),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1527),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1527),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1536),
.B(n_1486),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1520),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1530),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1530),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1534),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1535),
.B(n_1512),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1540),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1531),
.A2(n_1487),
.B1(n_1496),
.B2(n_1517),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1524),
.Y(n_1568)
);

NAND2xp33_ASAP7_75t_L g1569 ( 
.A(n_1543),
.B(n_1497),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1533),
.B(n_1499),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1523),
.B(n_1513),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1540),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1523),
.B(n_1513),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_L g1574 ( 
.A(n_1537),
.B(n_1512),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_1528),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1534),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1551),
.B(n_1538),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1537),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1549),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1565),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1565),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1569),
.A2(n_1526),
.B(n_1525),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_SL g1583 ( 
.A1(n_1575),
.A2(n_1528),
.B1(n_1372),
.B2(n_1535),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1561),
.A2(n_1532),
.B1(n_1529),
.B2(n_1541),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1565),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1574),
.Y(n_1586)
);

INVxp67_ASAP7_75t_SL g1587 ( 
.A(n_1568),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1569),
.A2(n_1512),
.B(n_1539),
.Y(n_1588)
);

OAI21xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1577),
.A2(n_1544),
.B(n_1538),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1568),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1571),
.B(n_1548),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1578),
.B(n_1549),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1564),
.B(n_1552),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1576),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1560),
.B(n_1556),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1562),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1568),
.Y(n_1597)
);

AOI21xp33_ASAP7_75t_SL g1598 ( 
.A1(n_1567),
.A2(n_1539),
.B(n_1546),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1594),
.Y(n_1599)
);

AOI222xp33_ASAP7_75t_L g1600 ( 
.A1(n_1586),
.A2(n_1560),
.B1(n_1573),
.B2(n_1563),
.C1(n_1579),
.C2(n_1572),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1593),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1582),
.A2(n_1577),
.B1(n_1566),
.B2(n_1557),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1580),
.B(n_1555),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1587),
.B(n_1555),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1581),
.B(n_1544),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1585),
.B(n_1558),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1590),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1597),
.B(n_1559),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1598),
.B(n_1546),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_SL g1610 ( 
.A1(n_1595),
.A2(n_1524),
.B(n_1514),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1609),
.B(n_1595),
.Y(n_1611)
);

NOR3xp33_ASAP7_75t_L g1612 ( 
.A(n_1604),
.B(n_1583),
.C(n_1589),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1600),
.A2(n_1584),
.B(n_1588),
.Y(n_1613)
);

AOI211xp5_ASAP7_75t_L g1614 ( 
.A1(n_1610),
.A2(n_1584),
.B(n_1592),
.C(n_1593),
.Y(n_1614)
);

AOI32xp33_ASAP7_75t_L g1615 ( 
.A1(n_1605),
.A2(n_1592),
.A3(n_1596),
.B1(n_1522),
.B2(n_1562),
.Y(n_1615)
);

A2O1A1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1602),
.A2(n_1591),
.B(n_1514),
.C(n_1522),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1602),
.B(n_1603),
.Y(n_1617)
);

AOI222xp33_ASAP7_75t_L g1618 ( 
.A1(n_1601),
.A2(n_1554),
.B1(n_1552),
.B2(n_1483),
.C1(n_1550),
.C2(n_1445),
.Y(n_1618)
);

NAND3xp33_ASAP7_75t_L g1619 ( 
.A(n_1599),
.B(n_1554),
.C(n_1570),
.Y(n_1619)
);

NOR3xp33_ASAP7_75t_SL g1620 ( 
.A(n_1606),
.B(n_1545),
.C(n_1292),
.Y(n_1620)
);

OAI221xp5_ASAP7_75t_L g1621 ( 
.A1(n_1613),
.A2(n_1607),
.B1(n_1608),
.B2(n_1570),
.C(n_1514),
.Y(n_1621)
);

OAI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1611),
.A2(n_1529),
.B1(n_1501),
.B2(n_1483),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1615),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1619),
.Y(n_1624)
);

XNOR2x1_ASAP7_75t_L g1625 ( 
.A(n_1612),
.B(n_1501),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1624),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1625),
.A2(n_1617),
.B(n_1614),
.Y(n_1627)
);

NAND3xp33_ASAP7_75t_L g1628 ( 
.A(n_1623),
.B(n_1616),
.C(n_1621),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1622),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1623),
.B(n_1620),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1625),
.B(n_1502),
.Y(n_1631)
);

XNOR2x1_ASAP7_75t_L g1632 ( 
.A(n_1628),
.B(n_1517),
.Y(n_1632)
);

AOI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1627),
.A2(n_1618),
.B1(n_1507),
.B2(n_1542),
.C(n_1500),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1631),
.B(n_1547),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1626),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1630),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1632),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1634),
.B(n_1629),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1636),
.A2(n_1633),
.B(n_1635),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1638),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1640),
.A2(n_1637),
.B1(n_1639),
.B2(n_1517),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1641),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1642),
.Y(n_1643)
);

OAI22xp33_ASAP7_75t_SL g1644 ( 
.A1(n_1643),
.A2(n_1547),
.B1(n_1553),
.B2(n_1500),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1644),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1645),
.A2(n_1502),
.B(n_1519),
.Y(n_1646)
);

AO22x2_ASAP7_75t_L g1647 ( 
.A1(n_1646),
.A2(n_1519),
.B1(n_1510),
.B2(n_1509),
.Y(n_1647)
);

XNOR2xp5_ASAP7_75t_L g1648 ( 
.A(n_1647),
.B(n_1515),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_SL g1649 ( 
.A1(n_1648),
.A2(n_1518),
.B1(n_1280),
.B2(n_1288),
.Y(n_1649)
);

AOI211xp5_ASAP7_75t_L g1650 ( 
.A1(n_1649),
.A2(n_1318),
.B(n_1280),
.C(n_1273),
.Y(n_1650)
);


endmodule