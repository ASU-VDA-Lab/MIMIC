module fake_jpeg_8591_n_170 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_5),
.B(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_1),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_14),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_22),
.Y(n_40)
);

AOI32xp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_33),
.A3(n_24),
.B1(n_32),
.B2(n_34),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_41),
.B(n_32),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_23),
.B1(n_28),
.B2(n_21),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_47),
.B1(n_54),
.B2(n_15),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_55),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_23),
.B1(n_27),
.B2(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_19),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_22),
.C(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_35),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_20),
.B1(n_27),
.B2(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_40),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_68),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_63),
.B(n_66),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_55),
.A2(n_24),
.B1(n_20),
.B2(n_16),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_46),
.Y(n_87)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_15),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_77),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_48),
.B1(n_42),
.B2(n_41),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_82),
.B1(n_54),
.B2(n_56),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_48),
.B1(n_42),
.B2(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_46),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_57),
.B1(n_60),
.B2(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_73),
.Y(n_101)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_100),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_61),
.B1(n_72),
.B2(n_58),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_106),
.B(n_107),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_40),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_78),
.C(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_30),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_89),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_69),
.B1(n_36),
.B2(n_34),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_79),
.A2(n_69),
.B1(n_36),
.B2(n_34),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_114),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_30),
.B(n_29),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_74),
.B(n_75),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_99),
.B(n_96),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_74),
.C(n_53),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_30),
.C(n_29),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_14),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_1),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_122),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_124),
.Y(n_139)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_99),
.B(n_97),
.C(n_103),
.D(n_107),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_111),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_122),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_132),
.C(n_113),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_117),
.B(n_120),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_3),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_133),
.B(n_2),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_127),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_141),
.C(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_140),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_144),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_109),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_30),
.C(n_12),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_12),
.C(n_10),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_134),
.B(n_2),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_144),
.C(n_130),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_126),
.B1(n_124),
.B2(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_149),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_125),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_152),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_123),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_148),
.A2(n_4),
.B(n_5),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_155),
.B1(n_9),
.B2(n_156),
.Y(n_161)
);

OAI31xp33_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_8),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_9),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_157),
.B(n_147),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_161),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_165),
.B(n_163),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_168),
.B(n_164),
.Y(n_169)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_166),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_165),
.Y(n_170)
);


endmodule