module real_jpeg_26194_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;
wire n_16;

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_0),
.B(n_32),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_0),
.B(n_29),
.Y(n_76)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_3),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_3),
.B(n_32),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_5),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_5),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_6),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_6),
.B(n_23),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_8),
.B(n_11),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_10),
.B(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_10),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_10),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_10),
.B(n_65),
.Y(n_78)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_70),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_48),
.C(n_49),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_34),
.C(n_39),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_26),
.B2(n_27),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_28),
.C(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.C(n_43),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_60),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_54),
.C(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_59),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_69),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_68),
.C(n_69),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_83),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);


endmodule