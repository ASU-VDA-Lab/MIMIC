module fake_aes_1378_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_5), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_9), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_12), .B(n_0), .Y(n_18) );
NOR2x1p5_ASAP7_75t_L g19 ( .A(n_15), .B(n_0), .Y(n_19) );
AOI221xp5_ASAP7_75t_L g20 ( .A1(n_16), .A2(n_1), .B1(n_2), .B2(n_8), .C(n_10), .Y(n_20) );
INVx2_ASAP7_75t_SL g21 ( .A(n_13), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx4_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_21), .Y(n_25) );
OAI21x1_ASAP7_75t_L g26 ( .A1(n_18), .A2(n_11), .B(n_14), .Y(n_26) );
BUFx3_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
AOI21xp5_ASAP7_75t_L g29 ( .A1(n_23), .A2(n_20), .B(n_11), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_23), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
NOR2x1_ASAP7_75t_L g32 ( .A(n_31), .B(n_19), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_30), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_29), .B1(n_24), .B2(n_26), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_32), .B(n_29), .Y(n_35) );
NAND2xp5_ASAP7_75t_L g36 ( .A(n_33), .B(n_25), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
AOI211xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_14), .B(n_30), .C(n_1), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
OAI221xp5_ASAP7_75t_R g41 ( .A1(n_40), .A2(n_2), .B1(n_24), .B2(n_34), .C(n_39), .Y(n_41) );
endmodule