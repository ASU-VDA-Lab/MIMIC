module fake_jpeg_28528_n_324 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_6),
.B(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_45),
.B(n_60),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_42),
.Y(n_47)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_0),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_24),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_17),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_52),
.Y(n_108)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_23),
.B(n_1),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_33),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_69),
.Y(n_85)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_25),
.B1(n_22),
.B2(n_37),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_72),
.A2(n_57),
.B1(n_69),
.B2(n_61),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_73),
.B(n_96),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_29),
.B(n_28),
.C(n_21),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_78),
.B(n_98),
.Y(n_134)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_90),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_60),
.Y(n_90)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_39),
.B1(n_26),
.B2(n_20),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_32),
.B1(n_26),
.B2(n_36),
.Y(n_136)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_24),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_40),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_24),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_40),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_35),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

CKINVDCx12_ASAP7_75t_R g103 ( 
.A(n_48),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_103),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_52),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_52),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_38),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_46),
.Y(n_144)
);

CKINVDCx9p33_ASAP7_75t_R g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_116),
.A2(n_129),
.B1(n_133),
.B2(n_125),
.Y(n_186)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_78),
.B(n_26),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_135),
.B(n_112),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_120),
.B(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_27),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_82),
.B(n_27),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_140),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_79),
.A2(n_25),
.B1(n_64),
.B2(n_68),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_46),
.C(n_54),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_151),
.C(n_71),
.Y(n_158)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_86),
.A2(n_30),
.B1(n_32),
.B2(n_36),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_83),
.B(n_35),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_136),
.A2(n_72),
.B1(n_87),
.B2(n_75),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_107),
.Y(n_162)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_144),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_96),
.A2(n_32),
.B1(n_31),
.B2(n_36),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_147),
.B1(n_34),
.B2(n_31),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_91),
.B(n_38),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_148),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_105),
.A2(n_34),
.B1(n_31),
.B2(n_20),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_88),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_34),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_152),
.A2(n_154),
.B1(n_159),
.B2(n_166),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_75),
.B1(n_84),
.B2(n_100),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_84),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_156),
.B(n_167),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_183),
.C(n_137),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_123),
.B(n_150),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_162),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_136),
.A2(n_107),
.B1(n_74),
.B2(n_20),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_23),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_109),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_170),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_77),
.B1(n_109),
.B2(n_71),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_169),
.A2(n_173),
.B1(n_179),
.B2(n_180),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_102),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_93),
.B1(n_81),
.B2(n_77),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_122),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_177),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_119),
.A2(n_81),
.B1(n_102),
.B2(n_69),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_76),
.B1(n_108),
.B2(n_85),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_176),
.A2(n_181),
.B1(n_125),
.B2(n_114),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_120),
.B(n_108),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_104),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_139),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_132),
.A2(n_69),
.B1(n_76),
.B2(n_85),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_151),
.A2(n_121),
.B1(n_124),
.B2(n_127),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_88),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_182),
.B(n_184),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_115),
.B(n_88),
.C(n_4),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_16),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_115),
.B(n_16),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_3),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_186),
.A2(n_150),
.B1(n_114),
.B2(n_125),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_142),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_187),
.B(n_207),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_208),
.Y(n_222)
);

XNOR2x1_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_183),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_191),
.B(n_181),
.Y(n_227)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_199),
.B1(n_202),
.B2(n_152),
.Y(n_228)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_156),
.A2(n_127),
.B1(n_143),
.B2(n_138),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_167),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_200),
.B(n_157),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_159),
.A2(n_138),
.B1(n_150),
.B2(n_118),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_205),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_204),
.A2(n_206),
.B1(n_176),
.B2(n_197),
.Y(n_235)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_118),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_131),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_216),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_153),
.A2(n_114),
.B(n_140),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_214),
.B(n_215),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_153),
.A2(n_3),
.B(n_6),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_153),
.A2(n_7),
.B(n_8),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_8),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_217),
.B(n_218),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_213),
.B(n_180),
.CI(n_158),
.CON(n_219),
.SN(n_219)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_193),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_239),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_182),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_226),
.C(n_242),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_169),
.Y(n_226)
);

AOI21x1_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_214),
.B(n_215),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_239),
.B1(n_240),
.B2(n_220),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_229),
.B(n_240),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_161),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_232),
.B(n_234),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_186),
.B(n_175),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_199),
.B(n_162),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_185),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_237),
.B1(n_211),
.B2(n_210),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_206),
.A2(n_187),
.B1(n_210),
.B2(n_201),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_173),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_208),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_188),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_252),
.C(n_260),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_248),
.A2(n_249),
.B1(n_227),
.B2(n_223),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_211),
.B1(n_195),
.B2(n_202),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_224),
.Y(n_280)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_201),
.C(n_212),
.Y(n_252)
);

AOI32xp33_ASAP7_75t_L g253 ( 
.A1(n_220),
.A2(n_193),
.A3(n_209),
.B1(n_200),
.B2(n_216),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_262),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_241),
.B(n_223),
.Y(n_276)
);

A2O1A1O1Ixp25_ASAP7_75t_L g258 ( 
.A1(n_222),
.A2(n_189),
.B(n_192),
.C(n_194),
.D(n_217),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_222),
.Y(n_265)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_175),
.A3(n_205),
.B1(n_218),
.B2(n_166),
.Y(n_259)
);

AO21x1_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_236),
.B(n_230),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_164),
.C(n_175),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_179),
.C(n_203),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_241),
.C(n_224),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_228),
.A2(n_196),
.B1(n_12),
.B2(n_14),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_229),
.B(n_9),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_263),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_279),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_233),
.B1(n_221),
.B2(n_235),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_269),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_236),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_280),
.Y(n_283)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_273),
.Y(n_286)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_249),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_276),
.A2(n_261),
.B(n_245),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_281),
.A2(n_276),
.B(n_277),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_264),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_285),
.Y(n_298)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_271),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_287),
.B(n_293),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_247),
.C(n_244),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_290),
.C(n_272),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_252),
.C(n_260),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_292),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_255),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_300),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_279),
.C(n_265),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_302),
.Y(n_310)
);

AOI31xp67_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_270),
.A3(n_258),
.B(n_278),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_269),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_267),
.B1(n_275),
.B2(n_266),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_284),
.B1(n_291),
.B2(n_245),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_280),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_284),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_277),
.C(n_251),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_238),
.B(n_243),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_292),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_309),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_238),
.B1(n_298),
.B2(n_243),
.Y(n_312)
);

NOR2x1_ASAP7_75t_SL g315 ( 
.A(n_308),
.B(n_294),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_273),
.A3(n_293),
.B1(n_269),
.B2(n_288),
.C1(n_259),
.C2(n_250),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_273),
.B1(n_283),
.B2(n_288),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_295),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_313),
.C(n_317),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_315),
.B(n_316),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_9),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_305),
.B(n_14),
.Y(n_319)
);

OAI221xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_311),
.B1(n_15),
.B2(n_16),
.C(n_12),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g321 ( 
.A(n_320),
.B(n_307),
.CI(n_312),
.CON(n_321),
.SN(n_321)
);

AOI211xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_322),
.B(n_318),
.C(n_15),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_307),
.Y(n_324)
);


endmodule