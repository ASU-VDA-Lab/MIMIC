module fake_aes_6366_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g11 ( .A(n_3), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_7), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_9), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_10), .B(n_9), .Y(n_17) );
NAND3xp33_ASAP7_75t_L g18 ( .A(n_16), .B(n_0), .C(n_8), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_14), .B(n_0), .Y(n_19) );
NOR2xp33_ASAP7_75t_SL g20 ( .A(n_16), .B(n_1), .Y(n_20) );
O2A1O1Ixp33_ASAP7_75t_L g21 ( .A1(n_16), .A2(n_2), .B(n_3), .C(n_4), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_11), .B(n_2), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
OAI22xp5_ASAP7_75t_L g24 ( .A1(n_18), .A2(n_11), .B1(n_15), .B2(n_13), .Y(n_24) );
AOI22xp5_ASAP7_75t_L g25 ( .A1(n_19), .A2(n_15), .B1(n_12), .B2(n_17), .Y(n_25) );
INVx1_ASAP7_75t_SL g26 ( .A(n_20), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
OAI222xp33_ASAP7_75t_L g28 ( .A1(n_24), .A2(n_21), .B1(n_18), .B2(n_6), .C1(n_7), .C2(n_8), .Y(n_28) );
BUFx2_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
AOI21xp5_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_23), .B(n_25), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_27), .Y(n_31) );
OR2x6_ASAP7_75t_L g32 ( .A(n_30), .B(n_29), .Y(n_32) );
OAI22xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_27), .B1(n_29), .B2(n_28), .Y(n_33) );
OAI21xp5_ASAP7_75t_SL g34 ( .A1(n_33), .A2(n_28), .B(n_29), .Y(n_34) );
INVx1_ASAP7_75t_SL g35 ( .A(n_32), .Y(n_35) );
INVx1_ASAP7_75t_SL g36 ( .A(n_35), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
AOI22xp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_4), .B1(n_5), .B2(n_36), .Y(n_38) );
endmodule