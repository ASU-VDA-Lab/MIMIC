module real_jpeg_2483_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_51),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_51),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_4),
.A2(n_31),
.B1(n_39),
.B2(n_40),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_4),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_5),
.A2(n_7),
.B(n_33),
.C(n_39),
.Y(n_32)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_5),
.A2(n_39),
.B(n_57),
.C(n_58),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_5),
.B(n_39),
.Y(n_57)
);

AO22x2_ASAP7_75t_L g58 ( 
.A1(n_5),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_7),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_7),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_7),
.B(n_58),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_7),
.B(n_24),
.C(n_47),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_7),
.B(n_21),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_7),
.B(n_68),
.Y(n_126)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_53),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_11),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_90),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_89),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_62),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_17),
.B(n_62),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_43),
.C(n_54),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_18),
.B(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_32),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_32),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B(n_27),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_24),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_20),
.A2(n_22),
.B1(n_29),
.B2(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_20),
.B(n_30),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_20),
.A2(n_29),
.B1(n_99),
.B2(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_21),
.A2(n_28),
.B(n_125),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_23),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_49)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_24),
.B(n_120),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_29),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B(n_36),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_35),
.A2(n_101),
.B(n_122),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_37),
.B(n_109),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_39),
.A2(n_40),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_43),
.B(n_54),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_44),
.A2(n_67),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_65),
.B(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_45),
.B(n_69),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_49),
.A2(n_50),
.B(n_95),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_59),
.B(n_60),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_71),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_85),
.B2(n_86),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_104),
.B(n_135),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_102),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.C(n_97),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_98),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_116),
.B(n_134),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_132),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_128),
.B(n_133),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_123),
.B(n_127),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_126),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_131),
.Y(n_133)
);


endmodule