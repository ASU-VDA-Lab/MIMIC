module real_aes_7669_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g511 ( .A1(n_0), .A2(n_154), .B(n_512), .C(n_513), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_1), .B(n_173), .Y(n_515) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_3), .A2(n_140), .B(n_145), .C(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_4), .A2(n_135), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_5), .B(n_210), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_6), .A2(n_102), .B1(n_115), .B2(n_750), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_7), .A2(n_135), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_8), .B(n_173), .Y(n_239) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_9), .A2(n_158), .B(n_466), .Y(n_465) );
AND2x6_ASAP7_75t_L g140 ( .A(n_10), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_11), .A2(n_140), .B(n_145), .C(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g152 ( .A(n_12), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_13), .B(n_42), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_14), .B(n_150), .Y(n_187) );
INVx1_ASAP7_75t_L g133 ( .A(n_15), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_16), .B(n_210), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_17), .A2(n_153), .B(n_167), .C(n_171), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_18), .B(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_19), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_20), .B(n_279), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_21), .A2(n_197), .B(n_198), .C(n_200), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_22), .A2(n_145), .B(n_214), .C(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_23), .B(n_150), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_24), .B(n_150), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g221 ( .A(n_25), .Y(n_221) );
INVx1_ASAP7_75t_L g209 ( .A(n_26), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_27), .A2(n_145), .B(n_214), .C(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_28), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_29), .Y(n_180) );
INVx1_ASAP7_75t_L g275 ( .A(n_30), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_31), .A2(n_135), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g138 ( .A(n_32), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_33), .A2(n_226), .B(n_447), .C(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_34), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_35), .A2(n_197), .B(n_235), .C(n_237), .Y(n_234) );
INVxp67_ASAP7_75t_L g276 ( .A(n_36), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_37), .B(n_471), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_38), .A2(n_145), .B(n_208), .C(n_214), .Y(n_207) );
CKINVDCx14_ASAP7_75t_R g233 ( .A(n_39), .Y(n_233) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_40), .A2(n_47), .B1(n_741), .B2(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_40), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_41), .A2(n_46), .B1(n_726), .B2(n_727), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_41), .Y(n_727) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_43), .A2(n_149), .B(n_151), .C(n_154), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_44), .B(n_270), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_45), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_46), .Y(n_726) );
INVx1_ASAP7_75t_L g742 ( .A(n_47), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_48), .B(n_210), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_49), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_50), .B(n_135), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_51), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_52), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_53), .A2(n_226), .B(n_447), .C(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g514 ( .A(n_54), .Y(n_514) );
INVx1_ASAP7_75t_L g449 ( .A(n_55), .Y(n_449) );
INVx1_ASAP7_75t_L g195 ( .A(n_56), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_57), .B(n_135), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_58), .Y(n_495) );
CKINVDCx14_ASAP7_75t_R g143 ( .A(n_59), .Y(n_143) );
INVx1_ASAP7_75t_L g141 ( .A(n_60), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_61), .B(n_135), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_62), .B(n_173), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_63), .A2(n_213), .B(n_460), .C(n_461), .Y(n_459) );
INVx1_ASAP7_75t_L g132 ( .A(n_64), .Y(n_132) );
INVx1_ASAP7_75t_SL g236 ( .A(n_65), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_66), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_67), .B(n_210), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_68), .B(n_173), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_69), .B(n_153), .Y(n_524) );
INVx1_ASAP7_75t_L g224 ( .A(n_70), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g510 ( .A(n_71), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_72), .B(n_186), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_73), .A2(n_145), .B(n_226), .C(n_500), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_74), .Y(n_458) );
INVx1_ASAP7_75t_L g108 ( .A(n_75), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_76), .A2(n_135), .B(n_142), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_77), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_78), .A2(n_135), .B(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_79), .A2(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g165 ( .A(n_80), .Y(n_165) );
CKINVDCx16_ASAP7_75t_R g206 ( .A(n_81), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_82), .B(n_185), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_83), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_84), .A2(n_135), .B(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g168 ( .A(n_85), .Y(n_168) );
INVx2_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
INVx1_ASAP7_75t_L g184 ( .A(n_87), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_88), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_89), .B(n_150), .Y(n_525) );
OR2x2_ASAP7_75t_L g110 ( .A(n_90), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g122 ( .A(n_90), .Y(n_122) );
OR2x2_ASAP7_75t_L g438 ( .A(n_90), .B(n_112), .Y(n_438) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_91), .A2(n_145), .B(n_223), .C(n_226), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_92), .B(n_135), .Y(n_479) );
INVx1_ASAP7_75t_L g482 ( .A(n_93), .Y(n_482) );
INVxp67_ASAP7_75t_L g462 ( .A(n_94), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_95), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_96), .B(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g199 ( .A(n_97), .Y(n_199) );
INVx1_ASAP7_75t_L g501 ( .A(n_98), .Y(n_501) );
INVx1_ASAP7_75t_L g521 ( .A(n_99), .Y(n_521) );
AND2x2_ASAP7_75t_L g452 ( .A(n_100), .B(n_129), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g751 ( .A(n_105), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g743 ( .A(n_110), .Y(n_743) );
INVx2_ASAP7_75t_L g749 ( .A(n_110), .Y(n_749) );
NOR2x2_ASAP7_75t_L g732 ( .A(n_111), .B(n_122), .Y(n_732) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g121 ( .A(n_112), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AO221x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_734), .B1(n_737), .B2(n_744), .C(n_746), .Y(n_115) );
OAI222xp33_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_724), .B1(n_725), .B2(n_728), .C1(n_731), .C2(n_733), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B1(n_435), .B2(n_439), .Y(n_117) );
AOI22x1_ASAP7_75t_SL g728 ( .A1(n_118), .A2(n_435), .B1(n_729), .B2(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g729 ( .A(n_123), .Y(n_729) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_365), .Y(n_123) );
NAND5xp2_ASAP7_75t_L g124 ( .A(n_125), .B(n_280), .C(n_312), .D(n_329), .E(n_352), .Y(n_124) );
AOI221xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_203), .B1(n_240), .B2(n_244), .C(n_248), .Y(n_125) );
INVx1_ASAP7_75t_L g392 ( .A(n_126), .Y(n_392) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_175), .Y(n_126) );
AND3x2_ASAP7_75t_L g367 ( .A(n_127), .B(n_177), .C(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_160), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_128), .B(n_246), .Y(n_245) );
BUFx3_ASAP7_75t_L g255 ( .A(n_128), .Y(n_255) );
AND2x2_ASAP7_75t_L g259 ( .A(n_128), .B(n_191), .Y(n_259) );
INVx2_ASAP7_75t_L g289 ( .A(n_128), .Y(n_289) );
OR2x2_ASAP7_75t_L g300 ( .A(n_128), .B(n_192), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_128), .B(n_176), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_128), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g379 ( .A(n_128), .B(n_192), .Y(n_379) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_134), .B(n_157), .Y(n_128) );
INVx1_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_129), .A2(n_181), .B(n_206), .C(n_207), .Y(n_205) );
INVx2_ASAP7_75t_L g229 ( .A(n_129), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_129), .A2(n_445), .B(n_446), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_129), .A2(n_479), .B(n_480), .Y(n_478) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_L g159 ( .A(n_130), .B(n_131), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
BUFx2_ASAP7_75t_L g270 ( .A(n_135), .Y(n_270) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g181 ( .A(n_136), .B(n_140), .Y(n_181) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g213 ( .A(n_137), .Y(n_213) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
INVx1_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
INVx1_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
INVx3_ASAP7_75t_L g153 ( .A(n_139), .Y(n_153) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
INVx1_ASAP7_75t_L g471 ( .A(n_139), .Y(n_471) );
INVx4_ASAP7_75t_SL g156 ( .A(n_140), .Y(n_156) );
BUFx3_ASAP7_75t_L g214 ( .A(n_140), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_SL g142 ( .A1(n_143), .A2(n_144), .B(n_148), .C(n_156), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_SL g164 ( .A1(n_144), .A2(n_156), .B(n_165), .C(n_166), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_SL g194 ( .A1(n_144), .A2(n_156), .B(n_195), .C(n_196), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_144), .A2(n_156), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g271 ( .A1(n_144), .A2(n_156), .B(n_272), .C(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g447 ( .A(n_144), .Y(n_447) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_144), .A2(n_156), .B(n_458), .C(n_459), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_SL g509 ( .A1(n_144), .A2(n_156), .B(n_510), .C(n_511), .Y(n_509) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx3_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_146), .Y(n_238) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g197 ( .A(n_150), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
INVx5_ASAP7_75t_L g210 ( .A(n_153), .Y(n_210) );
INVx2_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g171 ( .A(n_155), .Y(n_171) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_155), .Y(n_451) );
INVx1_ASAP7_75t_L g226 ( .A(n_156), .Y(n_226) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_158), .Y(n_162) );
INVx4_ASAP7_75t_L g174 ( .A(n_158), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_158), .A2(n_467), .B(n_468), .Y(n_466) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g267 ( .A(n_159), .Y(n_267) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_160), .Y(n_258) );
AND2x2_ASAP7_75t_L g320 ( .A(n_160), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_160), .B(n_176), .Y(n_339) );
INVx1_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
OR2x2_ASAP7_75t_L g247 ( .A(n_161), .B(n_176), .Y(n_247) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_161), .Y(n_254) );
AND2x2_ASAP7_75t_L g306 ( .A(n_161), .B(n_192), .Y(n_306) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_161), .B(n_175), .C(n_289), .Y(n_331) );
AND2x2_ASAP7_75t_L g396 ( .A(n_161), .B(n_177), .Y(n_396) );
AND2x2_ASAP7_75t_L g430 ( .A(n_161), .B(n_176), .Y(n_430) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_172), .Y(n_161) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_162), .A2(n_193), .B(n_202), .Y(n_192) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_162), .A2(n_231), .B(n_239), .Y(n_230) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_162), .A2(n_456), .B(n_463), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_169), .B(n_199), .Y(n_198) );
OAI22xp33_ASAP7_75t_L g274 ( .A1(n_169), .A2(n_210), .B1(n_275), .B2(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g460 ( .A(n_169), .Y(n_460) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g186 ( .A(n_170), .Y(n_186) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_173), .A2(n_508), .B(n_515), .Y(n_507) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_174), .B(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_174), .B(n_216), .Y(n_215) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_174), .A2(n_220), .B(n_227), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_174), .B(n_485), .Y(n_484) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_174), .A2(n_498), .B(n_505), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_174), .B(n_506), .Y(n_505) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_174), .A2(n_520), .B(n_526), .Y(n_519) );
INVxp67_ASAP7_75t_L g256 ( .A(n_175), .Y(n_256) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_191), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_176), .B(n_289), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_176), .B(n_320), .Y(n_328) );
AND2x2_ASAP7_75t_L g378 ( .A(n_176), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g406 ( .A(n_176), .Y(n_406) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g313 ( .A(n_177), .B(n_306), .Y(n_313) );
BUFx3_ASAP7_75t_L g345 ( .A(n_177), .Y(n_345) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_189), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_178), .B(n_495), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_181), .A2(n_221), .B(n_222), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_181), .A2(n_521), .B(n_522), .Y(n_520) );
O2A1O1Ixp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_187), .C(n_188), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_185), .A2(n_188), .B(n_224), .C(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_185), .A2(n_449), .B(n_450), .C(n_451), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_185), .A2(n_451), .B(n_482), .C(n_483), .Y(n_481) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g321 ( .A(n_191), .Y(n_321) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_192), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_197), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_197), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g473 ( .A(n_200), .Y(n_473) );
INVx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_203), .A2(n_381), .B1(n_383), .B2(n_384), .Y(n_380) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_217), .Y(n_203) );
AND2x2_ASAP7_75t_L g240 ( .A(n_204), .B(n_241), .Y(n_240) );
INVx3_ASAP7_75t_SL g251 ( .A(n_204), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_204), .B(n_284), .Y(n_316) );
OR2x2_ASAP7_75t_L g335 ( .A(n_204), .B(n_218), .Y(n_335) );
AND2x2_ASAP7_75t_L g340 ( .A(n_204), .B(n_292), .Y(n_340) );
AND2x2_ASAP7_75t_L g343 ( .A(n_204), .B(n_285), .Y(n_343) );
AND2x2_ASAP7_75t_L g355 ( .A(n_204), .B(n_230), .Y(n_355) );
AND2x2_ASAP7_75t_L g371 ( .A(n_204), .B(n_219), .Y(n_371) );
AND2x4_ASAP7_75t_L g374 ( .A(n_204), .B(n_242), .Y(n_374) );
OR2x2_ASAP7_75t_L g391 ( .A(n_204), .B(n_327), .Y(n_391) );
OR2x2_ASAP7_75t_L g422 ( .A(n_204), .B(n_264), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_204), .B(n_350), .Y(n_424) );
OR2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_215), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .C(n_212), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_210), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g512 ( .A(n_210), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_212), .A2(n_492), .B(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_213), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g298 ( .A(n_217), .B(n_262), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_217), .B(n_285), .Y(n_417) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_230), .Y(n_217) );
AND2x2_ASAP7_75t_L g250 ( .A(n_218), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g284 ( .A(n_218), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g292 ( .A(n_218), .B(n_264), .Y(n_292) );
AND2x2_ASAP7_75t_L g310 ( .A(n_218), .B(n_242), .Y(n_310) );
OR2x2_ASAP7_75t_L g327 ( .A(n_218), .B(n_285), .Y(n_327) );
INVx2_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
BUFx2_ASAP7_75t_L g243 ( .A(n_219), .Y(n_243) );
AND2x2_ASAP7_75t_L g350 ( .A(n_219), .B(n_230), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g279 ( .A(n_229), .Y(n_279) );
INVx2_ASAP7_75t_L g242 ( .A(n_230), .Y(n_242) );
INVx1_ASAP7_75t_L g362 ( .A(n_230), .Y(n_362) );
AND2x2_ASAP7_75t_L g412 ( .A(n_230), .B(n_251), .Y(n_412) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_238), .Y(n_503) );
AND2x2_ASAP7_75t_L g261 ( .A(n_241), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g296 ( .A(n_241), .B(n_251), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_241), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
AND2x2_ASAP7_75t_L g283 ( .A(n_242), .B(n_251), .Y(n_283) );
OR2x2_ASAP7_75t_L g399 ( .A(n_243), .B(n_373), .Y(n_399) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_246), .B(n_379), .Y(n_385) );
INVx2_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OAI32xp33_ASAP7_75t_L g341 ( .A1(n_247), .A2(n_342), .A3(n_344), .B1(n_346), .B2(n_347), .Y(n_341) );
OR2x2_ASAP7_75t_L g358 ( .A(n_247), .B(n_300), .Y(n_358) );
OAI21xp33_ASAP7_75t_SL g383 ( .A1(n_247), .A2(n_257), .B(n_288), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_252), .B1(n_257), .B2(n_260), .Y(n_248) );
INVxp33_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_250), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_251), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g309 ( .A(n_251), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g409 ( .A(n_251), .B(n_350), .Y(n_409) );
OR2x2_ASAP7_75t_L g433 ( .A(n_251), .B(n_327), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g416 ( .A1(n_252), .A2(n_315), .B(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_256), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g293 ( .A(n_254), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_254), .B(n_259), .Y(n_311) );
AND2x2_ASAP7_75t_L g333 ( .A(n_255), .B(n_306), .Y(n_333) );
INVx1_ASAP7_75t_L g346 ( .A(n_255), .Y(n_346) );
OR2x2_ASAP7_75t_L g351 ( .A(n_255), .B(n_285), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_258), .B(n_300), .Y(n_299) );
OAI22xp33_ASAP7_75t_L g281 ( .A1(n_259), .A2(n_282), .B1(n_287), .B2(n_291), .Y(n_281) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_262), .A2(n_324), .B1(n_331), .B2(n_332), .Y(n_330) );
AND2x2_ASAP7_75t_L g408 ( .A(n_262), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_264), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g427 ( .A(n_264), .B(n_310), .Y(n_427) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_268), .B(n_277), .Y(n_264) );
INVx1_ASAP7_75t_L g286 ( .A(n_265), .Y(n_286) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_267), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_269), .A2(n_278), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI21xp5_ASAP7_75t_SL g488 ( .A1(n_279), .A2(n_489), .B(n_490), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_293), .B1(n_294), .B2(n_299), .C(n_301), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_283), .B(n_285), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_283), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g302 ( .A(n_284), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g389 ( .A1(n_284), .A2(n_390), .B(n_391), .C(n_392), .Y(n_389) );
AND2x2_ASAP7_75t_L g394 ( .A(n_284), .B(n_374), .Y(n_394) );
O2A1O1Ixp33_ASAP7_75t_SL g432 ( .A1(n_284), .A2(n_373), .B(n_433), .C(n_434), .Y(n_432) );
BUFx3_ASAP7_75t_L g324 ( .A(n_285), .Y(n_324) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_288), .B(n_345), .Y(n_388) );
AOI211xp5_ASAP7_75t_L g407 ( .A1(n_288), .A2(n_408), .B(n_410), .C(n_416), .Y(n_407) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVxp67_ASAP7_75t_L g368 ( .A(n_290), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_292), .B(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AOI211xp5_ASAP7_75t_L g312 ( .A1(n_296), .A2(n_313), .B(n_314), .C(n_322), .Y(n_312) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g397 ( .A(n_300), .Y(n_397) );
OR2x2_ASAP7_75t_L g414 ( .A(n_300), .B(n_344), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_308), .B2(n_311), .Y(n_301) );
OAI22xp33_ASAP7_75t_L g314 ( .A1(n_303), .A2(n_315), .B1(n_316), .B2(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
OR2x2_ASAP7_75t_L g401 ( .A(n_305), .B(n_345), .Y(n_401) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g356 ( .A(n_306), .B(n_346), .Y(n_356) );
INVx1_ASAP7_75t_L g364 ( .A(n_307), .Y(n_364) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_310), .B(n_324), .Y(n_372) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_320), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g429 ( .A(n_321), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_325), .B(n_328), .Y(n_322) );
INVx1_ASAP7_75t_L g359 ( .A(n_323), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_324), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_324), .B(n_355), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g375 ( .A(n_324), .B(n_350), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_324), .B(n_371), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g386 ( .A1(n_324), .A2(n_334), .B(n_374), .C(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
AOI221xp5_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_334), .B1(n_336), .B2(n_340), .C(n_341), .Y(n_329) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVxp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_338), .B(n_346), .Y(n_420) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_L g431 ( .A1(n_340), .A2(n_355), .B(n_357), .C(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_343), .B(n_350), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_344), .B(n_397), .Y(n_434) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_345), .Y(n_344) );
INVxp33_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
AOI21xp33_ASAP7_75t_SL g360 ( .A1(n_349), .A2(n_361), .B(n_363), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_349), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_350), .B(n_404), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_356), .B1(n_357), .B2(n_359), .C(n_360), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_356), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g390 ( .A(n_362), .Y(n_390) );
NAND5xp2_ASAP7_75t_L g365 ( .A(n_366), .B(n_393), .C(n_407), .D(n_418), .E(n_431), .Y(n_365) );
AOI211xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B(n_376), .C(n_389), .Y(n_366) );
INVx2_ASAP7_75t_SL g413 ( .A(n_367), .Y(n_413) );
NAND4xp25_ASAP7_75t_SL g369 ( .A(n_370), .B(n_372), .C(n_373), .D(n_375), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI211xp5_ASAP7_75t_SL g376 ( .A1(n_375), .A2(n_377), .B(n_380), .C(n_386), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_378), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_378), .A2(n_419), .B1(n_421), .B2(n_423), .C(n_425), .Y(n_418) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI221xp5_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_395), .B1(n_398), .B2(n_400), .C(n_402), .Y(n_393) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_401), .A2(n_424), .B1(n_426), .B2(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx4_ASAP7_75t_L g730 ( .A(n_439), .Y(n_730) );
XOR2xp5_ASAP7_75t_L g739 ( .A(n_439), .B(n_740), .Y(n_739) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR5x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_597), .C(n_675), .D(n_699), .E(n_716), .Y(n_440) );
OAI211xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_474), .B(n_516), .C(n_574), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_453), .Y(n_442) );
AND2x2_ASAP7_75t_L g528 ( .A(n_443), .B(n_455), .Y(n_528) );
INVx5_ASAP7_75t_SL g556 ( .A(n_443), .Y(n_556) );
AND2x2_ASAP7_75t_L g592 ( .A(n_443), .B(n_577), .Y(n_592) );
OR2x2_ASAP7_75t_L g631 ( .A(n_443), .B(n_454), .Y(n_631) );
OR2x2_ASAP7_75t_L g662 ( .A(n_443), .B(n_553), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_443), .B(n_566), .Y(n_698) );
AND2x2_ASAP7_75t_L g710 ( .A(n_443), .B(n_553), .Y(n_710) );
OR2x6_ASAP7_75t_L g443 ( .A(n_444), .B(n_452), .Y(n_443) );
AND2x2_ASAP7_75t_L g709 ( .A(n_453), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g572 ( .A(n_454), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_464), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_455), .B(n_553), .Y(n_552) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_455), .Y(n_565) );
INVx3_ASAP7_75t_L g580 ( .A(n_455), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_455), .B(n_464), .Y(n_604) );
OR2x2_ASAP7_75t_L g613 ( .A(n_455), .B(n_556), .Y(n_613) );
AND2x2_ASAP7_75t_L g617 ( .A(n_455), .B(n_577), .Y(n_617) );
AND2x2_ASAP7_75t_L g623 ( .A(n_455), .B(n_624), .Y(n_623) );
INVxp67_ASAP7_75t_L g660 ( .A(n_455), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_455), .B(n_519), .Y(n_674) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_460), .A2(n_501), .B(n_502), .C(n_503), .Y(n_500) );
OR2x2_ASAP7_75t_L g566 ( .A(n_464), .B(n_519), .Y(n_566) );
AND2x2_ASAP7_75t_L g577 ( .A(n_464), .B(n_553), .Y(n_577) );
AND2x2_ASAP7_75t_L g589 ( .A(n_464), .B(n_580), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_464), .B(n_519), .Y(n_612) );
INVx1_ASAP7_75t_SL g624 ( .A(n_464), .Y(n_624) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g518 ( .A(n_465), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_465), .B(n_556), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_472), .B(n_473), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_473), .A2(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
AND2x2_ASAP7_75t_L g537 ( .A(n_476), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_476), .B(n_496), .Y(n_541) );
AND2x2_ASAP7_75t_L g544 ( .A(n_476), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_476), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g569 ( .A(n_476), .B(n_560), .Y(n_569) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_476), .Y(n_588) );
AND2x2_ASAP7_75t_L g609 ( .A(n_476), .B(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g619 ( .A(n_476), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g665 ( .A(n_476), .B(n_548), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_476), .B(n_571), .Y(n_692) );
INVx5_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g562 ( .A(n_477), .Y(n_562) );
AND2x2_ASAP7_75t_L g628 ( .A(n_477), .B(n_560), .Y(n_628) );
AND2x2_ASAP7_75t_L g712 ( .A(n_477), .B(n_580), .Y(n_712) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_484), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_486), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_486), .Y(n_701) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_496), .Y(n_486) );
AND2x2_ASAP7_75t_L g531 ( .A(n_487), .B(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g540 ( .A(n_487), .B(n_538), .Y(n_540) );
INVx5_ASAP7_75t_L g548 ( .A(n_487), .Y(n_548) );
AND2x2_ASAP7_75t_L g571 ( .A(n_487), .B(n_507), .Y(n_571) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_487), .Y(n_608) );
OR2x6_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .Y(n_487) );
INVx1_ASAP7_75t_L g649 ( .A(n_496), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_496), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g682 ( .A(n_496), .B(n_548), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g711 ( .A1(n_496), .A2(n_605), .B(n_712), .C(n_713), .Y(n_711) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_507), .Y(n_496) );
BUFx2_ASAP7_75t_L g532 ( .A(n_497), .Y(n_532) );
INVx2_ASAP7_75t_L g536 ( .A(n_497), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_504), .Y(n_498) );
INVx2_ASAP7_75t_L g538 ( .A(n_507), .Y(n_538) );
AND2x2_ASAP7_75t_L g545 ( .A(n_507), .B(n_536), .Y(n_545) );
AND2x2_ASAP7_75t_L g636 ( .A(n_507), .B(n_548), .Y(n_636) );
AOI211x1_ASAP7_75t_SL g516 ( .A1(n_517), .A2(n_529), .B(n_542), .C(n_567), .Y(n_516) );
INVx1_ASAP7_75t_L g633 ( .A(n_517), .Y(n_633) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_528), .Y(n_517) );
INVx5_ASAP7_75t_SL g553 ( .A(n_519), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_519), .B(n_623), .Y(n_622) );
AOI311xp33_ASAP7_75t_L g641 ( .A1(n_519), .A2(n_642), .A3(n_644), .B(n_645), .C(n_651), .Y(n_641) );
A2O1A1Ixp33_ASAP7_75t_L g676 ( .A1(n_519), .A2(n_589), .B(n_677), .C(n_680), .Y(n_676) );
INVxp67_ASAP7_75t_L g596 ( .A(n_528), .Y(n_596) );
NAND4xp25_ASAP7_75t_SL g529 ( .A(n_530), .B(n_533), .C(n_539), .D(n_541), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_530), .B(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g587 ( .A(n_531), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_537), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_534), .B(n_540), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_534), .B(n_547), .Y(n_667) );
BUFx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_535), .B(n_548), .Y(n_685) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g560 ( .A(n_536), .Y(n_560) );
INVxp67_ASAP7_75t_L g595 ( .A(n_537), .Y(n_595) );
AND2x4_ASAP7_75t_L g547 ( .A(n_538), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g621 ( .A(n_538), .B(n_560), .Y(n_621) );
INVx1_ASAP7_75t_L g648 ( .A(n_538), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_538), .B(n_635), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_539), .B(n_609), .Y(n_629) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_540), .B(n_562), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_540), .B(n_609), .Y(n_708) );
INVx1_ASAP7_75t_L g719 ( .A(n_541), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_546), .B(n_549), .C(n_557), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g561 ( .A(n_545), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g599 ( .A(n_545), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g581 ( .A(n_546), .Y(n_581) );
AND2x2_ASAP7_75t_L g558 ( .A(n_547), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_547), .B(n_609), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_547), .B(n_628), .Y(n_652) );
OR2x2_ASAP7_75t_L g568 ( .A(n_548), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g600 ( .A(n_548), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_548), .B(n_560), .Y(n_615) );
AND2x2_ASAP7_75t_L g672 ( .A(n_548), .B(n_628), .Y(n_672) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_548), .Y(n_679) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_550), .A2(n_562), .B1(n_684), .B2(n_686), .C(n_689), .Y(n_683) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g573 ( .A(n_553), .B(n_556), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_553), .B(n_623), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_553), .B(n_580), .Y(n_688) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g673 ( .A(n_555), .B(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g687 ( .A(n_555), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_556), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g584 ( .A(n_556), .B(n_577), .Y(n_584) );
AND2x2_ASAP7_75t_L g654 ( .A(n_556), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_556), .B(n_603), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_556), .B(n_704), .Y(n_703) );
OAI21xp5_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_561), .B(n_563), .Y(n_557) );
INVx2_ASAP7_75t_L g590 ( .A(n_558), .Y(n_590) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g610 ( .A(n_560), .Y(n_610) );
OR2x2_ASAP7_75t_L g614 ( .A(n_562), .B(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g717 ( .A(n_562), .B(n_685), .Y(n_717) );
INVx1_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AOI21xp33_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_570), .B(n_572), .Y(n_567) );
INVx1_ASAP7_75t_L g721 ( .A(n_568), .Y(n_721) );
INVx2_ASAP7_75t_SL g635 ( .A(n_569), .Y(n_635) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_572), .A2(n_653), .B(n_717), .C(n_718), .Y(n_716) );
OAI322xp33_ASAP7_75t_SL g585 ( .A1(n_573), .A2(n_586), .A3(n_589), .B1(n_590), .B2(n_591), .C1(n_593), .C2(n_596), .Y(n_585) );
INVx2_ASAP7_75t_L g605 ( .A(n_573), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_581), .B1(n_582), .B2(n_584), .C(n_585), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI22xp33_ASAP7_75t_SL g651 ( .A1(n_576), .A2(n_652), .B1(n_653), .B2(n_656), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_577), .B(n_580), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_577), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g650 ( .A(n_579), .B(n_612), .Y(n_650) );
INVx1_ASAP7_75t_L g640 ( .A(n_580), .Y(n_640) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_584), .A2(n_694), .B(n_696), .Y(n_693) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_586), .A2(n_619), .B(n_622), .Y(n_618) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NOR2xp67_ASAP7_75t_SL g647 ( .A(n_588), .B(n_648), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_588), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g704 ( .A(n_589), .Y(n_704) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND4xp25_ASAP7_75t_L g597 ( .A(n_598), .B(n_625), .C(n_641), .D(n_657), .Y(n_597) );
AOI211xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .B(n_606), .C(n_618), .Y(n_598) );
INVx1_ASAP7_75t_L g690 ( .A(n_599), .Y(n_690) );
AND2x2_ASAP7_75t_L g638 ( .A(n_600), .B(n_621), .Y(n_638) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_605), .B(n_640), .Y(n_639) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_611), .B1(n_614), .B2(n_616), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_608), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g656 ( .A(n_609), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_609), .A2(n_648), .B(n_671), .C(n_673), .Y(n_670) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g655 ( .A(n_612), .Y(n_655) );
INVx1_ASAP7_75t_L g715 ( .A(n_613), .Y(n_715) );
NAND2xp33_ASAP7_75t_SL g705 ( .A(n_614), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g644 ( .A(n_623), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_629), .B(n_630), .C(n_632), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_637), .B2(n_639), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_635), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_640), .B(n_661), .Y(n_723) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI21xp33_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_649), .B(n_650), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_663), .B1(n_666), .B2(n_668), .C(n_670), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_673), .A2(n_690), .B1(n_691), .B2(n_692), .Y(n_689) );
NAND3xp33_ASAP7_75t_SL g675 ( .A(n_676), .B(n_683), .C(n_693), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
CKINVDCx16_ASAP7_75t_R g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI211xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B(n_702), .C(n_711), .Y(n_699) );
INVx1_ASAP7_75t_L g720 ( .A(n_700), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .B1(n_707), .B2(n_709), .Y(n_702) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_718) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
CKINVDCx16_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g745 ( .A(n_736), .Y(n_745) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_743), .Y(n_738) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
endmodule