module fake_jpeg_29674_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_43;
wire n_37;
wire n_50;
wire n_29;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

OR2x2_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_5),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_0),
.Y(n_21)
);

OAI32xp33_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_17),
.A3(n_18),
.B1(n_10),
.B2(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_17),
.B1(n_13),
.B2(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_16),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

AND2x6_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_21),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

AND2x6_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_27),
.C(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.C(n_27),
.Y(n_44)
);

AND2x6_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_10),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_20),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_19),
.Y(n_50)
);

AOI321xp33_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_26),
.A3(n_19),
.B1(n_23),
.B2(n_28),
.C(n_29),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_39),
.B(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_50),
.B(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_56),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_57),
.C(n_28),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_1),
.B(n_2),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_62),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_28),
.C(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_47),
.B(n_29),
.C(n_26),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_26),
.B(n_29),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

AOI322xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_69),
.A3(n_66),
.B1(n_15),
.B2(n_64),
.C1(n_8),
.C2(n_9),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_6),
.B(n_7),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_65),
.B(n_2),
.Y(n_71)
);


endmodule