module fake_jpeg_29603_n_184 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_184);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_19),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_81),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_61),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_97),
.Y(n_111)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_92),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_60),
.B1(n_73),
.B2(n_72),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_96),
.B1(n_77),
.B2(n_65),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_55),
.C(n_66),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_74),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_58),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_98)
);

OR2x2_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_7),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_98),
.A2(n_75),
.B1(n_56),
.B2(n_71),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_118),
.Y(n_122)
);

BUFx2_ASAP7_75t_SL g103 ( 
.A(n_95),
.Y(n_103)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_57),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_109),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_68),
.B1(n_62),
.B2(n_52),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_9),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_70),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_1),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_5),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_5),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_8),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_6),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_8),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_62),
.B1(n_52),
.B2(n_68),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_34),
.B1(n_49),
.B2(n_47),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_6),
.B(n_7),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_119),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_127)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_124),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_127),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_33),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_20),
.C(n_22),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_134),
.B1(n_13),
.B2(n_14),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_133),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_32),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_135),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_137),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_108),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_119),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_41),
.C(n_43),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_154),
.B1(n_156),
.B2(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_148),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_125),
.B(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_147),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_24),
.B(n_28),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_157),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_29),
.B1(n_35),
.B2(n_37),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_128),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_159),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_123),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_120),
.B1(n_132),
.B2(n_45),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.C(n_144),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_172),
.B(n_167),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_164),
.C(n_170),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_176),
.B(n_162),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_173),
.C(n_166),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_178),
.A2(n_165),
.B(n_171),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_179),
.A2(n_155),
.B(n_160),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_181),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_145),
.A3(n_153),
.B1(n_169),
.B2(n_50),
.C1(n_150),
.C2(n_142),
.Y(n_183)
);

BUFx24_ASAP7_75t_SL g184 ( 
.A(n_183),
.Y(n_184)
);


endmodule