module fake_jpeg_12761_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_48),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx6p67_ASAP7_75t_R g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_20),
.B(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_58),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_39),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_7),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_59),
.A2(n_75),
.B(n_5),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_63),
.B(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_11),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_71),
.Y(n_99)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_74),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_76),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_78),
.Y(n_122)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_80),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_33),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_24),
.A2(n_11),
.B1(n_13),
.B2(n_2),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_42),
.B1(n_38),
.B2(n_37),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_85),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_28),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_60),
.A2(n_24),
.B1(n_29),
.B2(n_34),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_87),
.A2(n_89),
.B1(n_95),
.B2(n_100),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_29),
.B1(n_34),
.B2(n_40),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_40),
.C(n_28),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_93),
.B(n_117),
.CI(n_94),
.CON(n_170),
.SN(n_170)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_96),
.B(n_120),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_46),
.A2(n_29),
.B1(n_27),
.B2(n_37),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_18),
.B1(n_16),
.B2(n_21),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_110),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_45),
.A2(n_18),
.B1(n_16),
.B2(n_21),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_49),
.A2(n_42),
.B1(n_38),
.B2(n_0),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_132),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_53),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_54),
.A2(n_1),
.B1(n_12),
.B2(n_13),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_51),
.A2(n_12),
.B(n_13),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_116),
.B(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_55),
.B(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_65),
.B(n_14),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_1),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_14),
.B1(n_77),
.B2(n_75),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_127),
.B1(n_114),
.B2(n_119),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_43),
.B(n_52),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_43),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_132),
.B(n_124),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_52),
.B(n_57),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_57),
.B(n_44),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_138),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_122),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_136),
.B(n_162),
.Y(n_208)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_85),
.A2(n_96),
.B(n_119),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_141),
.A2(n_133),
.B(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_115),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_142),
.B(n_145),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_90),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_147),
.B(n_152),
.Y(n_179)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_83),
.A2(n_120),
.B(n_93),
.C(n_99),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_151),
.A2(n_165),
.A3(n_146),
.B1(n_153),
.B2(n_170),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_123),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_154),
.B(n_161),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_101),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_155),
.B(n_156),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_113),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

BUFx4f_ASAP7_75t_SL g181 ( 
.A(n_157),
.Y(n_181)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_82),
.B(n_104),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_106),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_106),
.B(n_104),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_164),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_113),
.B(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_126),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_127),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_170),
.Y(n_185)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_171),
.Y(n_186)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_174),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

BUFx8_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_108),
.B(n_130),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_162),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_166),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_133),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_198),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_141),
.A2(n_170),
.B1(n_139),
.B2(n_154),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_172),
.B1(n_158),
.B2(n_168),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_139),
.A2(n_165),
.B1(n_134),
.B2(n_136),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_SL g233 ( 
.A(n_195),
.B(n_188),
.C(n_207),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_196),
.B(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_149),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_161),
.B(n_153),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_138),
.B(n_137),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_202),
.B(n_183),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_159),
.A2(n_144),
.B1(n_171),
.B2(n_169),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_180),
.B1(n_208),
.B2(n_177),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_148),
.B(n_174),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_207),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_176),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_219),
.C(n_228),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_157),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_181),
.B1(n_189),
.B2(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_215),
.A2(n_216),
.B1(n_223),
.B2(n_224),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_193),
.A2(n_204),
.B1(n_178),
.B2(n_197),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_185),
.A2(n_205),
.B1(n_187),
.B2(n_201),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_221),
.B1(n_230),
.B2(n_211),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_142),
.C(n_173),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_191),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_222),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_143),
.B1(n_150),
.B2(n_180),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_203),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_199),
.B1(n_203),
.B2(n_200),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_199),
.B1(n_200),
.B2(n_194),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_186),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_183),
.B1(n_188),
.B2(n_194),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_190),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_190),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_181),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_233),
.A2(n_184),
.B(n_182),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_234),
.A2(n_243),
.B(n_223),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_236),
.A2(n_245),
.B1(n_247),
.B2(n_224),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_237),
.B(n_211),
.Y(n_255)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_242),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_221),
.B(n_218),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_215),
.A2(n_184),
.B1(n_189),
.B2(n_181),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_249),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_250),
.C(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_181),
.C(n_189),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_257),
.Y(n_271)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_244),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_253),
.B1(n_235),
.B2(n_240),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g261 ( 
.A(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_244),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_266),
.B1(n_238),
.B2(n_241),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_227),
.A3(n_225),
.B1(n_233),
.B2(n_226),
.C1(n_217),
.C2(n_229),
.Y(n_263)
);

AOI321xp33_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_238),
.A3(n_235),
.B1(n_237),
.B2(n_239),
.C(n_243),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_246),
.B(n_225),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_267),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_252),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_220),
.C(n_209),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_257),
.CI(n_250),
.CON(n_279),
.SN(n_279)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_189),
.Y(n_269)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_265),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_271),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_253),
.B1(n_236),
.B2(n_239),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_280),
.A2(n_266),
.B1(n_262),
.B2(n_267),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_286),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_278),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_287),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_264),
.B1(n_268),
.B2(n_259),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_255),
.B1(n_234),
.B2(n_254),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_289),
.C(n_291),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_293),
.B(n_294),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_279),
.C(n_272),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_275),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_290),
.B(n_282),
.Y(n_299)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_300),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_296),
.A2(n_282),
.B1(n_287),
.B2(n_286),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_295),
.A2(n_292),
.B1(n_294),
.B2(n_276),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_270),
.C(n_277),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_302),
.A2(n_297),
.B(n_279),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_304),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_305),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_310),
.C(n_301),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_300),
.C(n_299),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_303),
.Y(n_313)
);


endmodule