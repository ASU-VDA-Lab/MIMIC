module fake_jpeg_32197_n_138 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_138);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_0),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_58),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_55),
.Y(n_61)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_20),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_46),
.Y(n_70)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_71),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_46),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_57),
.B1(n_45),
.B2(n_51),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_1),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_94),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_59),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_90),
.Y(n_95)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_49),
.B(n_2),
.C(n_3),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_10),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_56),
.B1(n_44),
.B2(n_47),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_47),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_4),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_5),
.B(n_6),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_97),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_6),
.B(n_8),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_104),
.C(n_106),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_101),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_12),
.Y(n_101)
);

XOR2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_13),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_18),
.B(n_21),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g107 ( 
.A(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_109),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_22),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_24),
.C(n_26),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_28),
.C(n_29),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_32),
.Y(n_122)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_119),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_30),
.C(n_31),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_123),
.B(n_124),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_33),
.C(n_38),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_103),
.B(n_100),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_127),
.B(n_103),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_115),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_131),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_99),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_117),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_128),
.C(n_132),
.Y(n_136)
);

NAND2x1_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_126),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_114),
.Y(n_138)
);


endmodule