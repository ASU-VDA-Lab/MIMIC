module real_aes_9092_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_266;
wire n_183;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g167 ( .A1(n_0), .A2(n_168), .B(n_169), .C(n_173), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_1), .B(n_162), .Y(n_175) );
INVx1_ASAP7_75t_L g106 ( .A(n_2), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_3), .B(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_4), .A2(n_156), .B(n_465), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_5), .A2(n_136), .B(n_153), .C(n_509), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_6), .A2(n_156), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_7), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_8), .B(n_162), .Y(n_471) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_9), .A2(n_128), .B(n_250), .Y(n_249) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_10), .A2(n_441), .B1(n_711), .B2(n_714), .C1(n_718), .C2(n_719), .Y(n_440) );
AND2x6_ASAP7_75t_L g153 ( .A(n_11), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_12), .A2(n_136), .B(n_153), .C(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g562 ( .A(n_13), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_14), .B(n_40), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_14), .B(n_40), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_15), .B(n_172), .Y(n_511) );
INVx1_ASAP7_75t_L g133 ( .A(n_16), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_17), .B(n_147), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_18), .A2(n_148), .B(n_520), .C(n_522), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_19), .B(n_162), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_20), .B(n_190), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_21), .A2(n_136), .B(n_182), .C(n_189), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_22), .A2(n_171), .B(n_224), .C(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_23), .B(n_172), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_24), .B(n_172), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_25), .Y(n_489) );
INVx1_ASAP7_75t_L g459 ( .A(n_26), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_27), .A2(n_136), .B(n_189), .C(n_253), .Y(n_252) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_28), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_29), .Y(n_507) );
INVx1_ASAP7_75t_L g483 ( .A(n_30), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_31), .A2(n_156), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g138 ( .A(n_32), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_33), .A2(n_151), .B(n_205), .C(n_206), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_34), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_35), .A2(n_171), .B(n_468), .C(n_470), .Y(n_467) );
INVxp67_ASAP7_75t_L g484 ( .A(n_36), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_37), .B(n_255), .Y(n_254) );
CKINVDCx14_ASAP7_75t_R g466 ( .A(n_38), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_39), .A2(n_136), .B(n_189), .C(n_458), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_41), .A2(n_173), .B(n_560), .C(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_42), .B(n_180), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_43), .A2(n_102), .B1(n_110), .B2(n_724), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_44), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_45), .B(n_147), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_46), .B(n_156), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_47), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_48), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_49), .A2(n_151), .B(n_205), .C(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g170 ( .A(n_50), .Y(n_170) );
INVx1_ASAP7_75t_L g234 ( .A(n_51), .Y(n_234) );
INVx1_ASAP7_75t_L g527 ( .A(n_52), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_53), .B(n_156), .Y(n_231) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_54), .A2(n_71), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_54), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_55), .Y(n_194) );
CKINVDCx14_ASAP7_75t_R g558 ( .A(n_56), .Y(n_558) );
INVx1_ASAP7_75t_L g154 ( .A(n_57), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_58), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_59), .B(n_162), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_60), .A2(n_143), .B(n_188), .C(n_245), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_61), .A2(n_70), .B1(n_712), .B2(n_713), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_61), .Y(n_712) );
INVx1_ASAP7_75t_L g132 ( .A(n_62), .Y(n_132) );
INVx1_ASAP7_75t_SL g469 ( .A(n_63), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_64), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_65), .B(n_147), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_66), .B(n_162), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_67), .B(n_148), .Y(n_221) );
INVx1_ASAP7_75t_L g492 ( .A(n_68), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_69), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_70), .Y(n_713) );
INVx1_ASAP7_75t_L g120 ( .A(n_71), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_72), .B(n_184), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_73), .A2(n_136), .B(n_141), .C(n_151), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_74), .Y(n_243) );
INVx1_ASAP7_75t_L g109 ( .A(n_75), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_76), .A2(n_156), .B(n_557), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_77), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_78), .A2(n_156), .B(n_517), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_79), .A2(n_180), .B(n_479), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g456 ( .A(n_80), .Y(n_456) );
INVx1_ASAP7_75t_L g518 ( .A(n_81), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_82), .B(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_83), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_84), .A2(n_156), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g521 ( .A(n_85), .Y(n_521) );
INVx2_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
INVx1_ASAP7_75t_L g510 ( .A(n_87), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_88), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_89), .B(n_172), .Y(n_222) );
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_90), .B(n_106), .C(n_107), .Y(n_105) );
OR2x2_ASAP7_75t_L g432 ( .A(n_90), .B(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g445 ( .A(n_90), .B(n_434), .Y(n_445) );
INVx2_ASAP7_75t_L g710 ( .A(n_90), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_91), .A2(n_136), .B(n_151), .C(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_92), .B(n_156), .Y(n_203) );
INVx1_ASAP7_75t_L g207 ( .A(n_93), .Y(n_207) );
INVxp67_ASAP7_75t_L g246 ( .A(n_94), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_95), .B(n_128), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_96), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g142 ( .A(n_97), .Y(n_142) );
INVx1_ASAP7_75t_L g217 ( .A(n_98), .Y(n_217) );
INVx2_ASAP7_75t_L g530 ( .A(n_99), .Y(n_530) );
AND2x2_ASAP7_75t_L g236 ( .A(n_100), .B(n_192), .Y(n_236) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g725 ( .A(n_103), .Y(n_725) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x2_ASAP7_75t_L g434 ( .A(n_106), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
OA21x2_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_116), .B(n_439), .Y(n_110) );
BUFx2_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_SL g723 ( .A(n_114), .Y(n_723) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_431), .B(n_436), .Y(n_116) );
XNOR2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
INVx1_ASAP7_75t_L g442 ( .A(n_121), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_121), .A2(n_447), .B1(n_715), .B2(n_716), .Y(n_714) );
OR3x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_339), .C(n_388), .Y(n_121) );
NAND5xp2_ASAP7_75t_L g122 ( .A(n_123), .B(n_273), .C(n_302), .D(n_310), .E(n_325), .Y(n_122) );
O2A1O1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_196), .B(n_212), .C(n_257), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_176), .Y(n_124) );
AND2x2_ASAP7_75t_L g268 ( .A(n_125), .B(n_265), .Y(n_268) );
AND2x2_ASAP7_75t_L g301 ( .A(n_125), .B(n_177), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_125), .B(n_200), .Y(n_394) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_161), .Y(n_125) );
INVx2_ASAP7_75t_L g199 ( .A(n_126), .Y(n_199) );
BUFx2_ASAP7_75t_L g368 ( .A(n_126), .Y(n_368) );
AO21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_134), .B(n_159), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_127), .B(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g162 ( .A(n_127), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_127), .B(n_211), .Y(n_210) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_127), .A2(n_216), .B(n_226), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_127), .B(n_462), .Y(n_461) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_127), .A2(n_488), .B(n_495), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_127), .B(n_513), .Y(n_512) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_128), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_128), .A2(n_251), .B(n_252), .Y(n_250) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g228 ( .A(n_129), .Y(n_228) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g192 ( .A(n_130), .B(n_131), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_155), .Y(n_134) );
INVx5_ASAP7_75t_L g166 ( .A(n_136), .Y(n_166) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
BUFx3_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g158 ( .A(n_138), .Y(n_158) );
INVx1_ASAP7_75t_L g225 ( .A(n_138), .Y(n_225) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_140), .Y(n_145) );
INVx3_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
AND2x2_ASAP7_75t_L g157 ( .A(n_140), .B(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
INVx1_ASAP7_75t_L g255 ( .A(n_140), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_146), .C(n_149), .Y(n_141) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g482 ( .A1(n_144), .A2(n_147), .B1(n_483), .B2(n_484), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_144), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_144), .B(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
INVx2_ASAP7_75t_L g168 ( .A(n_147), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_147), .B(n_246), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_147), .A2(n_187), .B(n_459), .C(n_460), .Y(n_458) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_148), .B(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g470 ( .A(n_150), .Y(n_470) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_SL g164 ( .A1(n_152), .A2(n_165), .B(n_166), .C(n_167), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_152), .A2(n_166), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_152), .A2(n_166), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_152), .A2(n_166), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g517 ( .A1(n_152), .A2(n_166), .B(n_518), .C(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_SL g526 ( .A1(n_152), .A2(n_166), .B(n_527), .C(n_528), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_SL g557 ( .A1(n_152), .A2(n_166), .B(n_558), .C(n_559), .Y(n_557) );
INVx4_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g156 ( .A(n_153), .B(n_157), .Y(n_156) );
BUFx3_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g218 ( .A(n_153), .B(n_157), .Y(n_218) );
BUFx2_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
INVx1_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
AND2x2_ASAP7_75t_L g176 ( .A(n_161), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g266 ( .A(n_161), .Y(n_266) );
AND2x2_ASAP7_75t_L g352 ( .A(n_161), .B(n_265), .Y(n_352) );
AND2x2_ASAP7_75t_L g407 ( .A(n_161), .B(n_199), .Y(n_407) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_175), .Y(n_161) );
INVx2_ASAP7_75t_L g205 ( .A(n_166), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_171), .B(n_469), .Y(n_468) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g560 ( .A(n_172), .Y(n_560) );
INVx2_ASAP7_75t_L g494 ( .A(n_173), .Y(n_494) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_174), .Y(n_209) );
INVx1_ASAP7_75t_L g522 ( .A(n_174), .Y(n_522) );
INVx1_ASAP7_75t_L g324 ( .A(n_176), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_176), .B(n_200), .Y(n_371) );
INVx5_ASAP7_75t_L g265 ( .A(n_177), .Y(n_265) );
AND2x4_ASAP7_75t_L g286 ( .A(n_177), .B(n_266), .Y(n_286) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_177), .Y(n_308) );
AND2x2_ASAP7_75t_L g383 ( .A(n_177), .B(n_368), .Y(n_383) );
AND2x2_ASAP7_75t_L g386 ( .A(n_177), .B(n_201), .Y(n_386) );
OR2x6_ASAP7_75t_L g177 ( .A(n_178), .B(n_193), .Y(n_177) );
AOI21xp5_ASAP7_75t_SL g178 ( .A1(n_179), .A2(n_181), .B(n_190), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_185), .B(n_187), .Y(n_182) );
INVx2_ASAP7_75t_L g186 ( .A(n_184), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_186), .A2(n_207), .B(n_208), .C(n_209), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_186), .A2(n_209), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_186), .A2(n_492), .B(n_493), .C(n_494), .Y(n_491) );
O2A1O1Ixp5_ASAP7_75t_L g509 ( .A1(n_186), .A2(n_494), .B(n_510), .C(n_511), .Y(n_509) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_188), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_191), .B(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g195 ( .A(n_192), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_192), .A2(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_192), .A2(n_231), .B(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_192), .A2(n_218), .B(n_456), .C(n_457), .Y(n_455) );
OA21x2_ASAP7_75t_L g555 ( .A1(n_192), .A2(n_556), .B(n_563), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_195), .A2(n_506), .B(n_512), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_196), .B(n_266), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_196), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_200), .Y(n_197) );
AND2x2_ASAP7_75t_L g291 ( .A(n_198), .B(n_266), .Y(n_291) );
AND2x2_ASAP7_75t_L g309 ( .A(n_198), .B(n_201), .Y(n_309) );
INVx1_ASAP7_75t_L g329 ( .A(n_198), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_198), .B(n_265), .Y(n_374) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_198), .Y(n_416) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_199), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_200), .B(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_200), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_200), .A2(n_261), .B(n_322), .C(n_324), .Y(n_321) );
AND2x2_ASAP7_75t_L g328 ( .A(n_200), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g337 ( .A(n_200), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g341 ( .A(n_200), .B(n_265), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_200), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g356 ( .A(n_200), .B(n_266), .Y(n_356) );
AND2x2_ASAP7_75t_L g406 ( .A(n_200), .B(n_407), .Y(n_406) );
INVx5_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
BUFx2_ASAP7_75t_L g270 ( .A(n_201), .Y(n_270) );
AND2x2_ASAP7_75t_L g311 ( .A(n_201), .B(n_264), .Y(n_311) );
AND2x2_ASAP7_75t_L g323 ( .A(n_201), .B(n_298), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_201), .B(n_352), .Y(n_370) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_210), .Y(n_201) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_237), .Y(n_212) );
INVx1_ASAP7_75t_L g259 ( .A(n_213), .Y(n_259) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_229), .Y(n_213) );
OR2x2_ASAP7_75t_L g261 ( .A(n_214), .B(n_229), .Y(n_261) );
NAND3xp33_ASAP7_75t_L g267 ( .A(n_214), .B(n_268), .C(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_214), .B(n_239), .Y(n_278) );
OR2x2_ASAP7_75t_L g293 ( .A(n_214), .B(n_281), .Y(n_293) );
AND2x2_ASAP7_75t_L g299 ( .A(n_214), .B(n_248), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_214), .B(n_430), .Y(n_429) );
INVx5_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_215), .B(n_239), .Y(n_296) );
AND2x2_ASAP7_75t_L g335 ( .A(n_215), .B(n_249), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_215), .B(n_248), .Y(n_363) );
OR2x2_ASAP7_75t_L g366 ( .A(n_215), .B(n_248), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_219), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_218), .A2(n_489), .B(n_490), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_218), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_223), .A2(n_254), .B(n_256), .Y(n_253) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g477 ( .A(n_228), .Y(n_477) );
INVx5_ASAP7_75t_SL g281 ( .A(n_229), .Y(n_281) );
OR2x2_ASAP7_75t_L g287 ( .A(n_229), .B(n_238), .Y(n_287) );
AND2x2_ASAP7_75t_L g303 ( .A(n_229), .B(n_304), .Y(n_303) );
AOI321xp33_ASAP7_75t_L g310 ( .A1(n_229), .A2(n_311), .A3(n_312), .B1(n_313), .B2(n_319), .C(n_321), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_229), .B(n_237), .Y(n_320) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_229), .Y(n_333) );
OR2x2_ASAP7_75t_L g380 ( .A(n_229), .B(n_278), .Y(n_380) );
AND2x2_ASAP7_75t_L g402 ( .A(n_229), .B(n_299), .Y(n_402) );
AND2x2_ASAP7_75t_L g421 ( .A(n_229), .B(n_239), .Y(n_421) );
OR2x6_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_248), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_239), .B(n_248), .Y(n_262) );
AND2x2_ASAP7_75t_L g271 ( .A(n_239), .B(n_272), .Y(n_271) );
INVx3_ASAP7_75t_L g298 ( .A(n_239), .Y(n_298) );
AND2x2_ASAP7_75t_L g304 ( .A(n_239), .B(n_299), .Y(n_304) );
INVxp67_ASAP7_75t_L g334 ( .A(n_239), .Y(n_334) );
OR2x2_ASAP7_75t_L g376 ( .A(n_239), .B(n_281), .Y(n_376) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_247), .Y(n_239) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_240), .A2(n_464), .B(n_471), .Y(n_463) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_240), .A2(n_516), .B(n_523), .Y(n_515) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_240), .A2(n_525), .B(n_531), .Y(n_524) );
OR2x2_ASAP7_75t_L g258 ( .A(n_248), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_SL g272 ( .A(n_248), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_248), .B(n_261), .Y(n_305) );
AND2x2_ASAP7_75t_L g354 ( .A(n_248), .B(n_298), .Y(n_354) );
AND2x2_ASAP7_75t_L g392 ( .A(n_248), .B(n_281), .Y(n_392) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_249), .B(n_281), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_260), .B(n_263), .C(n_267), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_258), .A2(n_260), .B1(n_385), .B2(n_387), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_260), .A2(n_283), .B1(n_338), .B2(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_SL g412 ( .A(n_261), .Y(n_412) );
INVx1_ASAP7_75t_SL g312 ( .A(n_262), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_264), .B(n_284), .Y(n_314) );
AOI222xp33_ASAP7_75t_L g325 ( .A1(n_264), .A2(n_305), .B1(n_312), .B2(n_326), .C1(n_330), .C2(n_336), .Y(n_325) );
AND2x2_ASAP7_75t_L g415 ( .A(n_264), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g290 ( .A(n_265), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_265), .B(n_285), .Y(n_360) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_265), .Y(n_397) );
AND2x2_ASAP7_75t_L g400 ( .A(n_265), .B(n_309), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_265), .B(n_416), .Y(n_426) );
INVx1_ASAP7_75t_L g317 ( .A(n_266), .Y(n_317) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_266), .Y(n_345) );
O2A1O1Ixp33_ASAP7_75t_L g408 ( .A1(n_268), .A2(n_409), .B(n_410), .C(n_413), .Y(n_408) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_270), .B(n_332), .C(n_335), .Y(n_331) );
OR2x2_ASAP7_75t_L g359 ( .A(n_270), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_270), .B(n_286), .Y(n_387) );
OR2x2_ASAP7_75t_L g292 ( .A(n_272), .B(n_293), .Y(n_292) );
AOI211xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .B(n_282), .C(n_294), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_275), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g381 ( .A(n_276), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_277), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g295 ( .A(n_280), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_281), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g349 ( .A(n_281), .B(n_299), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_281), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_281), .B(n_298), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_287), .B1(n_288), .B2(n_292), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_284), .B(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_286), .B(n_328), .Y(n_327) );
OAI221xp5_ASAP7_75t_SL g350 ( .A1(n_287), .A2(n_351), .B1(n_353), .B2(n_355), .C(n_357), .Y(n_350) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x2_ASAP7_75t_L g405 ( .A(n_290), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g418 ( .A(n_290), .B(n_407), .Y(n_418) );
INVx1_ASAP7_75t_L g338 ( .A(n_291), .Y(n_338) );
INVx1_ASAP7_75t_L g409 ( .A(n_292), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_293), .A2(n_376), .B(n_399), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_297), .B(n_300), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OAI21xp5_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_305), .B(n_306), .Y(n_302) );
INVx1_ASAP7_75t_L g342 ( .A(n_303), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_304), .A2(n_390), .B1(n_393), .B2(n_395), .C(n_398), .Y(n_389) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_312), .A2(n_402), .B1(n_403), .B2(n_405), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g378 ( .A(n_314), .Y(n_378) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp67_ASAP7_75t_SL g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g382 ( .A(n_318), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g347 ( .A(n_323), .Y(n_347) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_328), .B(n_352), .Y(n_404) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_334), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g420 ( .A(n_335), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g427 ( .A(n_335), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI211xp5_ASAP7_75t_SL g339 ( .A1(n_340), .A2(n_342), .B(n_343), .C(n_377), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .B(n_350), .C(n_369), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g430 ( .A(n_354), .Y(n_430) );
AND2x2_ASAP7_75t_L g367 ( .A(n_356), .B(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_361), .B1(n_365), .B2(n_367), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
OR2x2_ASAP7_75t_L g375 ( .A(n_363), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g428 ( .A(n_364), .Y(n_428) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI31xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .A3(n_372), .B(n_375), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI211xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B(n_381), .C(n_384), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
CKINVDCx16_ASAP7_75t_R g385 ( .A(n_386), .Y(n_385) );
NAND5xp2_ASAP7_75t_L g388 ( .A(n_389), .B(n_401), .C(n_408), .D(n_422), .E(n_425), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_400), .A2(n_426), .B1(n_427), .B2(n_429), .Y(n_425) );
INVx1_ASAP7_75t_SL g424 ( .A(n_402), .Y(n_424) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_417), .B(n_419), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_432), .Y(n_438) );
NOR2x2_ASAP7_75t_L g721 ( .A(n_433), .B(n_710), .Y(n_721) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g709 ( .A(n_434), .B(n_710), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_436), .B(n_440), .C(n_722), .Y(n_439) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
OAI22xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_443), .B1(n_446), .B2(n_709), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g715 ( .A(n_444), .Y(n_715) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR3x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_620), .C(n_667), .Y(n_447) );
NAND3xp33_ASAP7_75t_SL g448 ( .A(n_449), .B(n_566), .C(n_591), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_504), .B1(n_532), .B2(n_535), .C(n_543), .Y(n_449) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_472), .B(n_497), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_452), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_452), .B(n_548), .Y(n_664) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_463), .Y(n_452) );
AND2x2_ASAP7_75t_L g534 ( .A(n_453), .B(n_503), .Y(n_534) );
AND2x2_ASAP7_75t_L g584 ( .A(n_453), .B(n_502), .Y(n_584) );
AND2x2_ASAP7_75t_L g605 ( .A(n_453), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g610 ( .A(n_453), .B(n_577), .Y(n_610) );
OR2x2_ASAP7_75t_L g618 ( .A(n_453), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g690 ( .A(n_453), .B(n_486), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_453), .B(n_639), .Y(n_704) );
INVx3_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g549 ( .A(n_454), .B(n_463), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_454), .B(n_486), .Y(n_550) );
AND2x4_ASAP7_75t_L g572 ( .A(n_454), .B(n_503), .Y(n_572) );
AND2x2_ASAP7_75t_L g602 ( .A(n_454), .B(n_474), .Y(n_602) );
AND2x2_ASAP7_75t_L g611 ( .A(n_454), .B(n_601), .Y(n_611) );
AND2x2_ASAP7_75t_L g627 ( .A(n_454), .B(n_487), .Y(n_627) );
OR2x2_ASAP7_75t_L g636 ( .A(n_454), .B(n_619), .Y(n_636) );
AND2x2_ASAP7_75t_L g642 ( .A(n_454), .B(n_577), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_454), .B(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g656 ( .A(n_454), .B(n_499), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_454), .B(n_545), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_454), .B(n_606), .Y(n_695) );
OR2x6_ASAP7_75t_L g454 ( .A(n_455), .B(n_461), .Y(n_454) );
INVx2_ASAP7_75t_L g503 ( .A(n_463), .Y(n_503) );
AND2x2_ASAP7_75t_L g601 ( .A(n_463), .B(n_486), .Y(n_601) );
AND2x2_ASAP7_75t_L g606 ( .A(n_463), .B(n_487), .Y(n_606) );
INVx1_ASAP7_75t_L g662 ( .A(n_463), .Y(n_662) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g571 ( .A(n_473), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_486), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_474), .B(n_534), .Y(n_533) );
BUFx3_ASAP7_75t_L g548 ( .A(n_474), .Y(n_548) );
OR2x2_ASAP7_75t_L g619 ( .A(n_474), .B(n_486), .Y(n_619) );
OR2x2_ASAP7_75t_L g680 ( .A(n_474), .B(n_587), .Y(n_680) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_478), .B(n_485), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_476), .A2(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g500 ( .A(n_478), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_485), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_486), .B(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g639 ( .A(n_486), .B(n_499), .Y(n_639) );
INVx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g578 ( .A(n_487), .Y(n_578) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_498), .A2(n_684), .B1(n_688), .B2(n_691), .C(n_692), .Y(n_683) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_502), .Y(n_498) );
INVx1_ASAP7_75t_SL g546 ( .A(n_499), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_499), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g678 ( .A(n_499), .B(n_534), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_502), .B(n_548), .Y(n_670) );
AND2x2_ASAP7_75t_L g577 ( .A(n_503), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_SL g581 ( .A(n_504), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_504), .B(n_587), .Y(n_617) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_514), .Y(n_504) );
AND2x2_ASAP7_75t_L g542 ( .A(n_505), .B(n_515), .Y(n_542) );
INVx4_ASAP7_75t_L g554 ( .A(n_505), .Y(n_554) );
BUFx3_ASAP7_75t_L g597 ( .A(n_505), .Y(n_597) );
AND3x2_ASAP7_75t_L g612 ( .A(n_505), .B(n_613), .C(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g694 ( .A(n_514), .B(n_608), .Y(n_694) );
AND2x2_ASAP7_75t_L g702 ( .A(n_514), .B(n_587), .Y(n_702) );
INVx1_ASAP7_75t_SL g707 ( .A(n_514), .Y(n_707) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
INVx1_ASAP7_75t_SL g565 ( .A(n_515), .Y(n_565) );
AND2x2_ASAP7_75t_L g588 ( .A(n_515), .B(n_554), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_515), .B(n_538), .Y(n_590) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_515), .Y(n_630) );
OR2x2_ASAP7_75t_L g635 ( .A(n_515), .B(n_554), .Y(n_635) );
INVx2_ASAP7_75t_L g540 ( .A(n_524), .Y(n_540) );
AND2x2_ASAP7_75t_L g575 ( .A(n_524), .B(n_555), .Y(n_575) );
OR2x2_ASAP7_75t_L g595 ( .A(n_524), .B(n_555), .Y(n_595) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_524), .Y(n_615) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AOI21xp33_ASAP7_75t_L g665 ( .A1(n_533), .A2(n_574), .B(n_666), .Y(n_665) );
AOI322xp5_ASAP7_75t_L g701 ( .A1(n_535), .A2(n_545), .A3(n_572), .B1(n_702), .B2(n_703), .C1(n_705), .C2(n_708), .Y(n_701) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_537), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_538), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g564 ( .A(n_539), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g632 ( .A(n_540), .B(n_554), .Y(n_632) );
AND2x2_ASAP7_75t_L g699 ( .A(n_540), .B(n_555), .Y(n_699) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g640 ( .A(n_542), .B(n_594), .Y(n_640) );
AOI31xp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_547), .A3(n_550), .B(n_551), .Y(n_543) );
AND2x2_ASAP7_75t_L g599 ( .A(n_545), .B(n_577), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_545), .B(n_569), .Y(n_681) );
AND2x2_ASAP7_75t_L g700 ( .A(n_545), .B(n_605), .Y(n_700) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_548), .B(n_577), .Y(n_589) );
NAND2x1p5_ASAP7_75t_L g623 ( .A(n_548), .B(n_606), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_548), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_548), .B(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_549), .B(n_606), .Y(n_638) );
INVx1_ASAP7_75t_L g682 ( .A(n_549), .Y(n_682) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_564), .Y(n_552) );
INVxp67_ASAP7_75t_L g634 ( .A(n_553), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_554), .B(n_565), .Y(n_570) );
INVx1_ASAP7_75t_L g676 ( .A(n_554), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_554), .B(n_653), .Y(n_687) );
BUFx3_ASAP7_75t_L g587 ( .A(n_555), .Y(n_587) );
AND2x2_ASAP7_75t_L g613 ( .A(n_555), .B(n_565), .Y(n_613) );
INVx2_ASAP7_75t_L g653 ( .A(n_555), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_564), .B(n_686), .Y(n_685) );
AOI211xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_571), .B(n_573), .C(n_582), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_568), .A2(n_617), .B(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_569), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_569), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g649 ( .A(n_570), .B(n_595), .Y(n_649) );
INVx3_ASAP7_75t_L g580 ( .A(n_572), .Y(n_580) );
OAI22xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_576), .B1(n_579), .B2(n_581), .Y(n_573) );
OAI21xp5_ASAP7_75t_SL g598 ( .A1(n_575), .A2(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g624 ( .A(n_575), .B(n_588), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_575), .B(n_676), .Y(n_675) );
INVxp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g579 ( .A(n_578), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g648 ( .A(n_578), .Y(n_648) );
OAI21xp5_ASAP7_75t_SL g592 ( .A1(n_579), .A2(n_593), .B(n_598), .Y(n_592) );
OAI22xp33_ASAP7_75t_SL g582 ( .A1(n_583), .A2(n_585), .B1(n_589), .B2(n_590), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_584), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g608 ( .A(n_587), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_587), .B(n_630), .Y(n_629) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_603), .C(n_616), .Y(n_591) );
OAI22xp5_ASAP7_75t_SL g658 ( .A1(n_593), .A2(n_659), .B1(n_663), .B2(n_664), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g663 ( .A(n_595), .B(n_596), .Y(n_663) );
AND2x2_ASAP7_75t_L g671 ( .A(n_596), .B(n_652), .Y(n_671) );
CKINVDCx16_ASAP7_75t_R g596 ( .A(n_597), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_SL g679 ( .A1(n_597), .A2(n_680), .B(n_681), .C(n_682), .Y(n_679) );
OR2x2_ASAP7_75t_L g706 ( .A(n_597), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_607), .B(n_609), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_L g641 ( .A1(n_605), .A2(n_642), .B(n_643), .C(n_646), .Y(n_641) );
OAI21xp33_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_611), .B(n_612), .Y(n_609) );
AND2x2_ASAP7_75t_L g674 ( .A(n_613), .B(n_632), .Y(n_674) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g652 ( .A(n_615), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g657 ( .A(n_617), .Y(n_657) );
NAND3xp33_ASAP7_75t_SL g620 ( .A(n_621), .B(n_641), .C(n_654), .Y(n_620) );
AOI211xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B(n_625), .C(n_633), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g691 ( .A(n_628), .Y(n_691) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g651 ( .A(n_630), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_630), .B(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B(n_636), .C(n_637), .Y(n_633) );
INVx2_ASAP7_75t_SL g645 ( .A(n_635), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_636), .A2(n_647), .B1(n_649), .B2(n_650), .Y(n_646) );
OAI21xp33_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B(n_658), .C(n_665), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVxp33_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g708 ( .A(n_662), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g667 ( .A(n_668), .B(n_683), .C(n_696), .D(n_701), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B(n_672), .C(n_679), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B(n_677), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g692 ( .A1(n_673), .A2(n_693), .B(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_680), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_700), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g717 ( .A(n_709), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_711), .Y(n_718) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx3_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
endmodule