module real_jpeg_2876_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_1),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_130),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_87),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_3),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_3),
.A2(n_63),
.B1(n_64),
.B2(n_87),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_27),
.C(n_29),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_4),
.A2(n_23),
.B1(n_42),
.B2(n_48),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_4),
.A2(n_29),
.B1(n_42),
.B2(n_52),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_4),
.A2(n_42),
.B1(n_63),
.B2(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_4),
.B(n_51),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_4),
.B(n_60),
.C(n_64),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_4),
.B(n_38),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_4),
.B(n_78),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_4),
.B(n_35),
.C(n_79),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_4),
.B(n_66),
.Y(n_174)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_7),
.A2(n_23),
.B1(n_40),
.B2(n_48),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_7),
.A2(n_29),
.B1(n_40),
.B2(n_52),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_7),
.A2(n_40),
.B1(n_63),
.B2(n_64),
.Y(n_83)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_212),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_191),
.B(n_211),
.Y(n_14)
);

OAI211xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_110),
.B(n_133),
.C(n_134),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_99),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_17),
.B(n_99),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_70),
.B2(n_71),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_18),
.B(n_73),
.C(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_43),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_20),
.B(n_45),
.C(n_55),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_21),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_26),
.Y(n_22)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_48),
.B(n_50),
.C(n_51),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_48),
.Y(n_50)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_27),
.A2(n_29),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_29),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_29),
.A2(n_52),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_29),
.B(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_31),
.A2(n_32),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_32),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_32),
.B(n_162),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_32),
.B(n_132),
.C(n_174),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_33),
.B(n_41),
.Y(n_89)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_34),
.A2(n_35),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_35),
.B(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_39),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_41),
.B(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_55),
.B2(n_69),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_44),
.A2(n_45),
.B1(n_92),
.B2(n_103),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_44),
.B(n_92),
.C(n_197),
.Y(n_234)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_51),
.B2(n_54),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_49),
.Y(n_226)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_54),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_107),
.C(n_108),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_55),
.A2(n_69),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_55),
.A2(n_230),
.B(n_233),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_55),
.B(n_230),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_66),
.B2(n_67),
.Y(n_55)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_66),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_68),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_58),
.A2(n_62),
.B(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

AOI22x1_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_64),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_64),
.B(n_167),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_90),
.B2(n_91),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_84),
.B2(n_85),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_85),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_74),
.A2(n_75),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_74),
.B(n_168),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_74),
.A2(n_75),
.B1(n_92),
.B2(n_103),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_74),
.B(n_92),
.C(n_182),
.Y(n_188)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_77),
.B(n_82),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_76),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_76),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_77),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_78),
.A2(n_209),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_82),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_88),
.B(n_89),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_88),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

OA21x2_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_89),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_88),
.B(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.C(n_95),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_94),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_96),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_95),
.B(n_118),
.C(n_123),
.Y(n_194)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_97),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.C(n_106),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_106),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_108),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_135),
.C(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_114),
.B(n_116),
.C(n_125),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_124),
.B2(n_125),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_127),
.B(n_131),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_129),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_132),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_131),
.A2(n_132),
.B1(n_146),
.B2(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_141),
.C(n_146),
.Y(n_140)
);

OAI21x1_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_153),
.B(n_190),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_140),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

NOR2xp67_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_165),
.Y(n_169)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_184),
.B(n_189),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_178),
.B(n_183),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_170),
.B(n_177),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_164),
.B(n_169),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_161),
.B(n_163),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_166),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_176),
.Y(n_177)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_180),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_188),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_193),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_196),
.C(n_201),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_210),
.Y(n_201)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_205),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_210),
.B1(n_224),
.B2(n_227),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_235),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_216),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_234),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_228),
.B2(n_229),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_224),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);


endmodule