module fake_jpeg_7085_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx5_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_2),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_23),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_7),
.A2(n_14),
.B1(n_13),
.B2(n_8),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

AOI322xp5_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_3),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_8),
.A2(n_4),
.B1(n_9),
.B2(n_12),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_11),
.A2(n_7),
.B1(n_10),
.B2(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_17),
.Y(n_38)
);

AND2x6_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_11),
.Y(n_34)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_12),
.C(n_11),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_21),
.B(n_18),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.C(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_39),
.Y(n_40)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_33),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_34),
.A3(n_37),
.B1(n_33),
.B2(n_40),
.C1(n_32),
.C2(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_42),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_43),
.B(n_16),
.C(n_26),
.Y(n_46)
);


endmodule