module fake_netlist_1_646_n_650 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_650);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_650;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_75), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_43), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_41), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_53), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_9), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_72), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_74), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_1), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_60), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_63), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_76), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_28), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_51), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_52), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_48), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_46), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_10), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_54), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_10), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_6), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_9), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_50), .Y(n_99) );
NOR2xp67_ASAP7_75t_L g100 ( .A(n_71), .B(n_11), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_5), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_73), .Y(n_102) );
INVxp33_ASAP7_75t_L g103 ( .A(n_42), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_18), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_38), .Y(n_105) );
INVxp33_ASAP7_75t_L g106 ( .A(n_33), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_44), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_23), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_22), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_57), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_35), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_13), .Y(n_112) );
INVxp33_ASAP7_75t_L g113 ( .A(n_58), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_18), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_59), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_13), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_27), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_6), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_29), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_16), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_30), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_32), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_34), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_65), .Y(n_124) );
INVxp33_ASAP7_75t_SL g125 ( .A(n_39), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_110), .B(n_94), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_116), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_98), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_99), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_123), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_114), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_121), .B(n_0), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_105), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_80), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_116), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_116), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_80), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_103), .B(n_0), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_78), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_78), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_125), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_95), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_88), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_87), .B(n_1), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_85), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_85), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_95), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_79), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
BUFx2_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_95), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_87), .B(n_2), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_89), .B(n_3), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_121), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_89), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_102), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_106), .B(n_4), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_90), .Y(n_161) );
BUFx2_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_83), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_90), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_88), .B(n_5), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_121), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_86), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_166), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_166), .B(n_112), .Y(n_171) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_166), .B(n_124), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_139), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_139), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_168), .B(n_113), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_145), .A2(n_82), .B1(n_120), .B2(n_101), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_126), .B(n_124), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_152), .B(n_101), .Y(n_180) );
AO22x2_ASAP7_75t_L g181 ( .A1(n_166), .A2(n_91), .B1(n_119), .B2(n_93), .Y(n_181) );
OAI21xp33_ASAP7_75t_L g182 ( .A1(n_141), .A2(n_91), .B(n_92), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_128), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_152), .B(n_112), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_144), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_162), .B(n_104), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_153), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_162), .B(n_104), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_159), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_159), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g194 ( .A1(n_147), .A2(n_97), .B1(n_118), .B2(n_119), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_159), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_133), .Y(n_196) );
AND2x4_ASAP7_75t_SL g197 ( .A(n_140), .B(n_97), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_157), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_141), .B(n_108), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_131), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_133), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_142), .B(n_108), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_132), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_142), .B(n_118), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_136), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_148), .B(n_92), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_150), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_157), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_158), .B(n_93), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_158), .B(n_109), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_157), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_136), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_135), .B(n_109), .Y(n_215) );
OR2x2_ASAP7_75t_SL g216 ( .A(n_146), .B(n_117), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_149), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_149), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_127), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_140), .B(n_111), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_127), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_151), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_137), .Y(n_223) );
BUFx4f_ASAP7_75t_L g224 ( .A(n_161), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_151), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_143), .B(n_111), .Y(n_226) );
XOR2xp5_ASAP7_75t_L g227 ( .A(n_129), .B(n_7), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_161), .B(n_165), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_209), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_185), .B(n_160), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_173), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_185), .B(n_160), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_209), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_220), .B(n_163), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_220), .B(n_165), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_173), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_184), .B(n_130), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_213), .Y(n_238) );
INVx1_ASAP7_75t_SL g239 ( .A(n_200), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_181), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_178), .Y(n_241) );
AOI22xp5_ASAP7_75t_SL g242 ( .A1(n_227), .A2(n_188), .B1(n_185), .B2(n_208), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_213), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_218), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_172), .A2(n_147), .B1(n_154), .B2(n_155), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_172), .Y(n_246) );
NAND2xp33_ASAP7_75t_L g247 ( .A(n_172), .B(n_121), .Y(n_247) );
BUFx10_ASAP7_75t_L g248 ( .A(n_185), .Y(n_248) );
BUFx12f_ASAP7_75t_L g249 ( .A(n_208), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_188), .B(n_100), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_213), .Y(n_251) );
INVx4_ASAP7_75t_L g252 ( .A(n_203), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_178), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_198), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_186), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_186), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_207), .B(n_138), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_189), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_188), .Y(n_260) );
AND2x6_ASAP7_75t_SL g261 ( .A(n_215), .B(n_115), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_198), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_188), .B(n_137), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_207), .B(n_138), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_224), .B(n_117), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_197), .B(n_115), .Y(n_266) );
NOR3xp33_ASAP7_75t_SL g267 ( .A(n_194), .B(n_134), .C(n_81), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_204), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_218), .Y(n_269) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_228), .A2(n_122), .B(n_102), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_181), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_182), .A2(n_122), .B(n_102), .C(n_107), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_224), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_205), .B(n_84), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_205), .B(n_122), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_189), .Y(n_276) );
O2A1O1Ixp5_ASAP7_75t_L g277 ( .A1(n_224), .A2(n_107), .B(n_164), .C(n_156), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_190), .Y(n_278) );
CKINVDCx8_ASAP7_75t_R g279 ( .A(n_171), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_190), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_197), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_195), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_197), .B(n_107), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_195), .Y(n_284) );
INVx1_ASAP7_75t_SL g285 ( .A(n_180), .Y(n_285) );
INVx4_ASAP7_75t_L g286 ( .A(n_203), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_171), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_203), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_180), .B(n_7), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_203), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_219), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_291), .A2(n_169), .B(n_171), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_230), .B(n_191), .Y(n_293) );
OR2x6_ASAP7_75t_L g294 ( .A(n_246), .B(n_181), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_248), .B(n_191), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_239), .B(n_177), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_230), .B(n_205), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_230), .B(n_205), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_240), .A2(n_181), .B1(n_171), .B2(n_169), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_237), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_291), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_246), .B(n_211), .Y(n_302) );
INVx4_ASAP7_75t_SL g303 ( .A(n_246), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_248), .B(n_211), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_231), .Y(n_305) );
INVx5_ASAP7_75t_L g306 ( .A(n_252), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_231), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_236), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_230), .B(n_232), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_260), .B(n_211), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_240), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_248), .B(n_211), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_252), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_236), .Y(n_314) );
OAI22xp5_ASAP7_75t_SL g315 ( .A1(n_249), .A2(n_227), .B1(n_194), .B2(n_177), .Y(n_315) );
AOI22x1_ASAP7_75t_L g316 ( .A1(n_241), .A2(n_174), .B1(n_170), .B2(n_187), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_252), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_271), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_232), .B(n_179), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_271), .A2(n_182), .B1(n_223), .B2(n_221), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_285), .B(n_176), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_252), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_241), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_232), .B(n_226), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_253), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_232), .B(n_199), .Y(n_326) );
INVx4_ASAP7_75t_L g327 ( .A(n_248), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_260), .A2(n_223), .B1(n_221), .B2(n_219), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_253), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_259), .Y(n_330) );
OR2x6_ASAP7_75t_L g331 ( .A(n_287), .B(n_202), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_259), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_286), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_255), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_290), .A2(n_210), .B(n_170), .Y(n_335) );
BUFx10_ASAP7_75t_L g336 ( .A(n_268), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_286), .Y(n_337) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_245), .A2(n_201), .B(n_206), .C(n_174), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_290), .A2(n_193), .B(n_183), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g340 ( .A(n_267), .B(n_201), .C(n_206), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_255), .Y(n_341) );
OR2x6_ASAP7_75t_L g342 ( .A(n_287), .B(n_214), .Y(n_342) );
OAI21xp33_ASAP7_75t_L g343 ( .A1(n_321), .A2(n_234), .B(n_237), .Y(n_343) );
BUFx2_ASAP7_75t_SL g344 ( .A(n_306), .Y(n_344) );
OA21x2_ASAP7_75t_L g345 ( .A1(n_316), .A2(n_272), .B(n_277), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_295), .B(n_289), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_294), .A2(n_279), .B1(n_281), .B2(n_235), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_301), .Y(n_348) );
NAND3xp33_ASAP7_75t_L g349 ( .A(n_338), .B(n_247), .C(n_242), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_305), .Y(n_350) );
AO31x2_ASAP7_75t_L g351 ( .A1(n_301), .A2(n_299), .A3(n_314), .B(n_334), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_306), .Y(n_352) );
AOI221x1_ASAP7_75t_L g353 ( .A1(n_305), .A2(n_250), .B1(n_275), .B2(n_151), .C(n_167), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_296), .A2(n_287), .B1(n_289), .B2(n_266), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_303), .B(n_286), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_292), .A2(n_256), .B(n_258), .Y(n_356) );
AOI22xp33_ASAP7_75t_SL g357 ( .A1(n_300), .A2(n_242), .B1(n_249), .B2(n_266), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_303), .B(n_286), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_296), .A2(n_250), .B1(n_283), .B2(n_263), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_315), .A2(n_250), .B1(n_283), .B2(n_263), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_315), .A2(n_250), .B1(n_264), .B2(n_274), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g362 ( .A1(n_335), .A2(n_278), .B(n_284), .Y(n_362) );
INVx4_ASAP7_75t_L g363 ( .A(n_294), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_314), .Y(n_364) );
AOI322xp5_ASAP7_75t_L g365 ( .A1(n_293), .A2(n_264), .A3(n_257), .B1(n_261), .B2(n_217), .C1(n_187), .C2(n_183), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_295), .B(n_256), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_294), .A2(n_258), .B1(n_284), .B2(n_282), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_336), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_336), .Y(n_369) );
AND2x6_ASAP7_75t_L g370 ( .A(n_302), .B(n_279), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_327), .B(n_273), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_319), .B(n_216), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_294), .A2(n_282), .B1(n_280), .B2(n_278), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_329), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_326), .B(n_261), .Y(n_375) );
NOR2x1_ASAP7_75t_L g376 ( .A(n_344), .B(n_331), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_343), .A2(n_331), .B1(n_324), .B2(n_311), .Y(n_377) );
AOI33xp33_ASAP7_75t_L g378 ( .A1(n_361), .A2(n_328), .A3(n_193), .B1(n_192), .B2(n_217), .B3(n_216), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_360), .A2(n_309), .B1(n_298), .B2(n_297), .C(n_329), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_363), .B(n_307), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_363), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_350), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_368), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_363), .A2(n_311), .B1(n_318), .B2(n_331), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_375), .A2(n_334), .B1(n_340), .B2(n_341), .C(n_307), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_357), .A2(n_331), .B1(n_318), .B2(n_302), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_367), .A2(n_320), .B1(n_341), .B2(n_323), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_365), .B(n_302), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_350), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_359), .A2(n_308), .B1(n_323), .B2(n_325), .C(n_276), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_370), .A2(n_312), .B1(n_304), .B2(n_336), .Y(n_391) );
OA21x2_ASAP7_75t_L g392 ( .A1(n_353), .A2(n_316), .B(n_325), .Y(n_392) );
OA21x2_ASAP7_75t_L g393 ( .A1(n_353), .A2(n_308), .B(n_320), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_370), .A2(n_304), .B1(n_312), .B2(n_310), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_373), .A2(n_310), .B1(n_276), .B2(n_280), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_362), .A2(n_339), .B(n_322), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_347), .A2(n_310), .B1(n_342), .B2(n_306), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_370), .A2(n_342), .B1(n_265), .B2(n_327), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_366), .B(n_303), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_370), .A2(n_342), .B1(n_327), .B2(n_306), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_364), .B(n_306), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_368), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_348), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_399), .B(n_364), .Y(n_404) );
AND2x2_ASAP7_75t_SL g405 ( .A(n_381), .B(n_355), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_403), .B(n_348), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_380), .Y(n_407) );
OAI31xp33_ASAP7_75t_SL g408 ( .A1(n_384), .A2(n_349), .A3(n_366), .B(n_374), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_382), .Y(n_409) );
OAI21xp33_ASAP7_75t_L g410 ( .A1(n_378), .A2(n_354), .B(n_346), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_403), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_379), .A2(n_370), .B1(n_372), .B2(n_344), .Y(n_412) );
OAI21xp5_ASAP7_75t_SL g413 ( .A1(n_386), .A2(n_369), .B(n_358), .Y(n_413) );
BUFx2_ASAP7_75t_L g414 ( .A(n_376), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_392), .A2(n_356), .B(n_345), .Y(n_415) );
OR2x6_ASAP7_75t_L g416 ( .A(n_397), .B(n_355), .Y(n_416) );
AND2x4_ASAP7_75t_SL g417 ( .A(n_399), .B(n_355), .Y(n_417) );
OAI322xp33_ASAP7_75t_L g418 ( .A1(n_388), .A2(n_372), .A3(n_374), .B1(n_214), .B2(n_196), .C1(n_192), .C2(n_167), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_397), .A2(n_370), .B1(n_352), .B2(n_358), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_376), .Y(n_420) );
AOI222xp33_ASAP7_75t_L g421 ( .A1(n_385), .A2(n_303), .B1(n_358), .B2(n_352), .C1(n_214), .C2(n_196), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_377), .A2(n_395), .B1(n_399), .B2(n_394), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_380), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_403), .B(n_351), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_382), .B(n_351), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_389), .B(n_351), .Y(n_426) );
NOR2xp67_ASAP7_75t_L g427 ( .A(n_401), .B(n_352), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_401), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_389), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_399), .B(n_330), .Y(n_430) );
NAND2xp33_ASAP7_75t_R g431 ( .A(n_381), .B(n_8), .Y(n_431) );
OAI33xp33_ASAP7_75t_L g432 ( .A1(n_395), .A2(n_371), .A3(n_11), .B1(n_12), .B2(n_14), .B3(n_15), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g433 ( .A1(n_387), .A2(n_270), .B(n_342), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_396), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_390), .B(n_351), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_391), .B(n_351), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_396), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_402), .B(n_270), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_412), .A2(n_387), .B1(n_383), .B2(n_400), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_425), .B(n_393), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_405), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_424), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_425), .B(n_393), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_424), .Y(n_444) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_428), .Y(n_445) );
AND2x6_ASAP7_75t_L g446 ( .A(n_435), .B(n_313), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_409), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_411), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_409), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_416), .Y(n_451) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_413), .A2(n_398), .B1(n_196), .B2(n_214), .C(n_393), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_405), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_434), .Y(n_454) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_405), .A2(n_393), .B1(n_392), .B2(n_333), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_429), .B(n_270), .Y(n_456) );
AOI33xp33_ASAP7_75t_L g457 ( .A1(n_422), .A2(n_8), .A3(n_12), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_416), .B(n_164), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_429), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_426), .B(n_392), .Y(n_461) );
AND2x4_ASAP7_75t_SL g462 ( .A(n_416), .B(n_337), .Y(n_462) );
AOI21xp5_ASAP7_75t_SL g463 ( .A1(n_416), .A2(n_392), .B(n_332), .Y(n_463) );
INVx3_ASAP7_75t_L g464 ( .A(n_416), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_423), .B(n_436), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_434), .Y(n_466) );
AND2x2_ASAP7_75t_SL g467 ( .A(n_408), .B(n_345), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_437), .Y(n_468) );
NAND4xp25_ASAP7_75t_L g469 ( .A(n_431), .B(n_408), .C(n_413), .D(n_410), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_406), .B(n_17), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_406), .B(n_17), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_414), .B(n_164), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_437), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_427), .Y(n_474) );
AOI33xp33_ASAP7_75t_L g475 ( .A1(n_419), .A2(n_222), .A3(n_225), .B1(n_262), .B2(n_254), .B3(n_333), .Y(n_475) );
AND2x2_ASAP7_75t_SL g476 ( .A(n_435), .B(n_345), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_414), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_438), .B(n_196), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_420), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_427), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_404), .B(n_345), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_404), .B(n_254), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_421), .B(n_151), .C(n_164), .Y(n_483) );
NAND2x1_ASAP7_75t_SL g484 ( .A(n_404), .B(n_337), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_404), .B(n_156), .Y(n_485) );
BUFx2_ASAP7_75t_L g486 ( .A(n_417), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_460), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_447), .B(n_410), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_470), .B(n_417), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_447), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_449), .Y(n_491) );
INVx2_ASAP7_75t_SL g492 ( .A(n_486), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_449), .B(n_415), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_459), .B(n_433), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_445), .Y(n_495) );
AND2x2_ASAP7_75t_SL g496 ( .A(n_486), .B(n_417), .Y(n_496) );
NOR2x1p5_ASAP7_75t_L g497 ( .A(n_469), .B(n_418), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_465), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_479), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_456), .B(n_430), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_483), .A2(n_418), .B(n_432), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_456), .B(n_156), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_469), .B(n_19), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_479), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_471), .B(n_20), .Y(n_505) );
AND2x2_ASAP7_75t_SL g506 ( .A(n_451), .B(n_337), .Y(n_506) );
NAND2xp33_ASAP7_75t_R g507 ( .A(n_451), .B(n_21), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_439), .A2(n_164), .B1(n_167), .B2(n_156), .C(n_262), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_471), .Y(n_509) );
AOI22xp33_ASAP7_75t_R g510 ( .A1(n_474), .A2(n_24), .B1(n_25), .B2(n_26), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_442), .B(n_167), .Y(n_511) );
AND3x1_ASAP7_75t_L g512 ( .A(n_457), .B(n_313), .C(n_317), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_442), .B(n_167), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_484), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_480), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_485), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_444), .B(n_167), .Y(n_517) );
NAND2xp33_ASAP7_75t_SL g518 ( .A(n_441), .B(n_313), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_444), .B(n_164), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_485), .Y(n_520) );
NAND2x1_ASAP7_75t_L g521 ( .A(n_441), .B(n_322), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_458), .Y(n_522) );
BUFx3_ASAP7_75t_L g523 ( .A(n_482), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_448), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_453), .B(n_31), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_453), .B(n_330), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_440), .B(n_332), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_440), .B(n_244), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_448), .B(n_244), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_443), .B(n_36), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_475), .B(n_175), .C(n_212), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_450), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_450), .B(n_244), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g534 ( .A(n_458), .B(n_322), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_450), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_498), .B(n_443), .Y(n_536) );
BUFx2_ASAP7_75t_SL g537 ( .A(n_509), .Y(n_537) );
OAI221xp5_ASAP7_75t_L g538 ( .A1(n_503), .A2(n_452), .B1(n_483), .B2(n_464), .C(n_484), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_495), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_487), .Y(n_540) );
NAND2x1_ASAP7_75t_SL g541 ( .A(n_522), .B(n_464), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_515), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_501), .A2(n_463), .B(n_455), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_497), .A2(n_464), .B1(n_462), .B2(n_458), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_512), .A2(n_446), .B1(n_464), .B2(n_458), .Y(n_545) );
OAI222xp33_ASAP7_75t_L g546 ( .A1(n_489), .A2(n_478), .B1(n_477), .B2(n_481), .C1(n_472), .C2(n_461), .Y(n_546) );
NAND4xp25_ASAP7_75t_L g547 ( .A(n_507), .B(n_463), .C(n_478), .D(n_481), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_490), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_496), .A2(n_462), .B1(n_477), .B2(n_467), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_491), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_501), .A2(n_467), .B(n_472), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_520), .B(n_477), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_506), .A2(n_467), .B1(n_455), .B2(n_476), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_499), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_516), .A2(n_446), .B1(n_476), .B2(n_472), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_505), .A2(n_446), .B1(n_476), .B2(n_461), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_492), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_504), .B(n_446), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_523), .A2(n_473), .B1(n_468), .B2(n_466), .Y(n_559) );
AOI21xp33_ASAP7_75t_L g560 ( .A1(n_502), .A2(n_473), .B(n_468), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_500), .B(n_446), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_502), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_488), .B(n_446), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_519), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_524), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_534), .A2(n_473), .B1(n_468), .B2(n_466), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_494), .B(n_446), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_527), .B(n_466), .Y(n_568) );
NAND3xp33_ASAP7_75t_L g569 ( .A(n_510), .B(n_454), .C(n_175), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_493), .B(n_454), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_494), .B(n_454), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_518), .A2(n_317), .B1(n_244), .B2(n_273), .Y(n_572) );
INVx2_ASAP7_75t_SL g573 ( .A(n_534), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_510), .B(n_175), .C(n_212), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_532), .Y(n_575) );
OAI321xp33_ASAP7_75t_L g576 ( .A1(n_525), .A2(n_212), .A3(n_175), .B1(n_225), .B2(n_222), .C(n_49), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_535), .B(n_37), .Y(n_577) );
INVxp33_ASAP7_75t_L g578 ( .A(n_530), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_565), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_539), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_568), .B(n_522), .Y(n_581) );
NOR3xp33_ASAP7_75t_SL g582 ( .A(n_569), .B(n_531), .C(n_508), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_536), .B(n_528), .Y(n_583) );
AOI211x1_ASAP7_75t_L g584 ( .A1(n_551), .A2(n_511), .B(n_513), .C(n_517), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_537), .Y(n_585) );
AOI21xp33_ASAP7_75t_L g586 ( .A1(n_578), .A2(n_514), .B(n_521), .Y(n_586) );
AOI21xp33_ASAP7_75t_SL g587 ( .A1(n_544), .A2(n_549), .B(n_553), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_543), .B(n_514), .Y(n_588) );
OAI22xp33_ASAP7_75t_SL g589 ( .A1(n_557), .A2(n_526), .B1(n_511), .B2(n_529), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_554), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_540), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_542), .B(n_533), .Y(n_592) );
NOR4xp25_ASAP7_75t_SL g593 ( .A(n_538), .B(n_508), .C(n_45), .D(n_47), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_548), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_550), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_562), .B(n_40), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_575), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_552), .B(n_55), .Y(n_598) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_574), .B(n_317), .Y(n_599) );
OAI21xp33_ASAP7_75t_SL g600 ( .A1(n_545), .A2(n_56), .B(n_61), .Y(n_600) );
NOR3xp33_ASAP7_75t_SL g601 ( .A(n_547), .B(n_62), .C(n_64), .Y(n_601) );
NOR4xp25_ASAP7_75t_SL g602 ( .A(n_576), .B(n_66), .C(n_67), .D(n_68), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_571), .Y(n_603) );
NOR2x1_ASAP7_75t_L g604 ( .A(n_546), .B(n_269), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_556), .B(n_212), .C(n_175), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_570), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_570), .B(n_69), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_567), .B(n_70), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_559), .Y(n_609) );
NAND3x2_ASAP7_75t_L g610 ( .A(n_583), .B(n_541), .C(n_555), .Y(n_610) );
BUFx2_ASAP7_75t_L g611 ( .A(n_585), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_609), .A2(n_561), .B1(n_563), .B2(n_564), .Y(n_612) );
OA22x2_ASAP7_75t_L g613 ( .A1(n_588), .A2(n_573), .B1(n_558), .B2(n_566), .Y(n_613) );
AOI221x1_ASAP7_75t_L g614 ( .A1(n_587), .A2(n_560), .B1(n_577), .B2(n_572), .C(n_212), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_588), .A2(n_577), .B(n_269), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_606), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_589), .B(n_233), .Y(n_617) );
OAI21xp5_ASAP7_75t_SL g618 ( .A1(n_604), .A2(n_288), .B(n_77), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_599), .Y(n_619) );
BUFx2_ASAP7_75t_L g620 ( .A(n_581), .Y(n_620) );
AOI31xp33_ASAP7_75t_SL g621 ( .A1(n_586), .A2(n_243), .A3(n_251), .B(n_238), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_603), .B(n_175), .Y(n_622) );
OAI21xp33_ASAP7_75t_SL g623 ( .A1(n_581), .A2(n_243), .B(n_251), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_600), .A2(n_259), .B(n_269), .Y(n_624) );
OAI21xp33_ASAP7_75t_SL g625 ( .A1(n_591), .A2(n_580), .B(n_594), .Y(n_625) );
OAI222xp33_ASAP7_75t_L g626 ( .A1(n_613), .A2(n_592), .B1(n_595), .B2(n_590), .C1(n_598), .C2(n_608), .Y(n_626) );
NOR2x1p5_ASAP7_75t_L g627 ( .A(n_613), .B(n_605), .Y(n_627) );
XNOR2x1_ASAP7_75t_L g628 ( .A(n_610), .B(n_608), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_616), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_625), .A2(n_601), .B(n_582), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_620), .Y(n_631) );
NAND2xp33_ASAP7_75t_SL g632 ( .A(n_617), .B(n_593), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_614), .A2(n_607), .B(n_596), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_612), .A2(n_584), .B1(n_597), .B2(n_579), .C(n_602), .Y(n_634) );
NAND5xp2_ASAP7_75t_L g635 ( .A(n_615), .B(n_229), .C(n_233), .D(n_288), .E(n_619), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_623), .A2(n_229), .B1(n_621), .B2(n_622), .C(n_624), .Y(n_636) );
OA22x2_ASAP7_75t_L g637 ( .A1(n_611), .A2(n_229), .B1(n_585), .B2(n_537), .Y(n_637) );
AOI211xp5_ASAP7_75t_L g638 ( .A1(n_618), .A2(n_229), .B(n_587), .C(n_625), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_631), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_629), .Y(n_640) );
AOI211xp5_ASAP7_75t_L g641 ( .A1(n_630), .A2(n_632), .B(n_626), .C(n_634), .Y(n_641) );
XNOR2xp5_ASAP7_75t_L g642 ( .A(n_628), .B(n_627), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_637), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_639), .Y(n_644) );
NOR3xp33_ASAP7_75t_SL g645 ( .A(n_642), .B(n_632), .C(n_635), .Y(n_645) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_644), .Y(n_646) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_644), .Y(n_647) );
OAI22xp5_ASAP7_75t_SL g648 ( .A1(n_646), .A2(n_641), .B1(n_643), .B2(n_645), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_648), .A2(n_647), .B1(n_638), .B2(n_640), .Y(n_649) );
AOI21xp33_ASAP7_75t_L g650 ( .A1(n_649), .A2(n_633), .B(n_636), .Y(n_650) );
endmodule