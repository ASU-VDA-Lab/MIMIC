module fake_jpeg_7704_n_90 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_2),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_59),
.Y(n_70)
);

AND2x4_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_0),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_64),
.B(n_66),
.C(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_56),
.B1(n_48),
.B2(n_53),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_47),
.B1(n_45),
.B2(n_44),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_76),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_0),
.B1(n_3),
.B2(n_6),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_78),
.B(n_79),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_77),
.B1(n_74),
.B2(n_75),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_75),
.B(n_72),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_82),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_12),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_13),
.C(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_17),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_18),
.A3(n_20),
.B1(n_22),
.B2(n_24),
.C1(n_25),
.C2(n_28),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_30),
.C(n_33),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_35),
.B(n_36),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_38),
.C(n_39),
.Y(n_90)
);


endmodule