module fake_jpeg_17733_n_216 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g16 ( 
.A(n_1),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_40),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_25),
.Y(n_51)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_25),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_58),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_22),
.B1(n_17),
.B2(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_41),
.B1(n_38),
.B2(n_39),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_22),
.B1(n_17),
.B2(n_24),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_53),
.A2(n_54),
.B1(n_41),
.B2(n_38),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_22),
.B1(n_30),
.B2(n_24),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_26),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_57),
.B1(n_39),
.B2(n_44),
.Y(n_102)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_64),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_79),
.Y(n_93)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_77),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_23),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_21),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_21),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_89),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_57),
.B1(n_39),
.B2(n_46),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_20),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_53),
.B(n_36),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_43),
.B(n_36),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_28),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_44),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_55),
.B1(n_57),
.B2(n_46),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_104),
.B1(n_90),
.B2(n_87),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_102),
.B1(n_114),
.B2(n_49),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_36),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_36),
.C(n_35),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_46),
.B1(n_44),
.B2(n_43),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_36),
.B(n_67),
.Y(n_135)
);

BUFx24_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_111),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_28),
.B1(n_27),
.B2(n_30),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_117),
.B1(n_126),
.B2(n_97),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_95),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_136),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_78),
.B(n_76),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_76),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_111),
.C(n_35),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_69),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_124),
.B(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_76),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_84),
.B1(n_91),
.B2(n_70),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_68),
.Y(n_127)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_94),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_68),
.Y(n_130)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_63),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_133),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_65),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_138),
.B(n_108),
.Y(n_150)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_108),
.Y(n_152)
);

NAND2x1_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_49),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_109),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_150),
.B(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_132),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_123),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_145),
.C(n_158),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_136),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_92),
.C(n_104),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_138),
.C(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_117),
.B1(n_121),
.B2(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

NAND4xp25_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_77),
.C(n_132),
.D(n_64),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

XOR2x1_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_163),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_151),
.A2(n_134),
.B(n_119),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_164),
.A2(n_165),
.B(n_170),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_151),
.A2(n_122),
.B1(n_113),
.B2(n_72),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_113),
.B1(n_74),
.B2(n_27),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_166),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_111),
.B(n_33),
.C(n_29),
.D(n_19),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_158),
.B(n_147),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_10),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_149),
.B(n_143),
.Y(n_177)
);

OA21x2_ASAP7_75t_SL g172 ( 
.A1(n_140),
.A2(n_12),
.B(n_11),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_154),
.Y(n_184)
);

OAI321xp33_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_19),
.A3(n_33),
.B1(n_29),
.B2(n_11),
.C(n_5),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_139),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_145),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_182),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_183),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_148),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_147),
.B(n_155),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_185),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_1),
.C(n_2),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_173),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_187),
.A2(n_193),
.B(n_194),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_163),
.B(n_165),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_160),
.B(n_171),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_167),
.C(n_148),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_203),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_169),
.C(n_190),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_182),
.C(n_176),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_202),
.C(n_159),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_144),
.C(n_180),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_188),
.B(n_192),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_206),
.C(n_208),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_196),
.C(n_190),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_180),
.Y(n_210)
);

NAND3xp33_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_211),
.C(n_212),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_205),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_162),
.B1(n_198),
.B2(n_6),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_SL g213 ( 
.A(n_209),
.B(n_162),
.C(n_4),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_213),
.A2(n_3),
.B1(n_7),
.B2(n_42),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_214),
.Y(n_216)
);


endmodule