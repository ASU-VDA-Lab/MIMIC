module fake_jpeg_16372_n_96 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_96);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVxp67_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_27),
.Y(n_33)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_30),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_13),
.B1(n_22),
.B2(n_20),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_40),
.B1(n_29),
.B2(n_14),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_13),
.B1(n_22),
.B2(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_13),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_1),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_19),
.B(n_16),
.C(n_15),
.Y(n_51)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_52),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_43),
.B(n_37),
.C(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_32),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_62),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_41),
.C(n_33),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_60),
.C(n_48),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_31),
.C(n_36),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_68),
.C(n_60),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_45),
.B(n_51),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_67),
.B(n_57),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_53),
.B1(n_39),
.B2(n_50),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_42),
.B(n_54),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_47),
.C(n_31),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_57),
.B(n_59),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_71),
.Y(n_79)
);

AOI322xp5_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_42),
.A3(n_12),
.B1(n_23),
.B2(n_19),
.C1(n_16),
.C2(n_15),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_73),
.Y(n_77)
);

OA21x2_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_39),
.B(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_75),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_31),
.C(n_17),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_80),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_52),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_80),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_68),
.C(n_74),
.Y(n_84)
);

AOI321xp33_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_78),
.A3(n_73),
.B1(n_72),
.B2(n_10),
.C(n_11),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_2),
.B(n_3),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_88),
.B(n_2),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_76),
.B1(n_52),
.B2(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_87),
.B(n_83),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_52),
.B1(n_44),
.B2(n_38),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_84),
.C(n_17),
.Y(n_91)
);

AOI322xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_91),
.A3(n_92),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_6),
.C(n_8),
.Y(n_94)
);

NOR4xp25_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_9),
.C(n_6),
.D(n_8),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_9),
.Y(n_96)
);


endmodule