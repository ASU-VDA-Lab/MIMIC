module real_aes_6904_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_769;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_785;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_314;
wire n_283;
wire n_741;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_371;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_SL g492 ( .A1(n_0), .A2(n_241), .B1(n_493), .B2(n_494), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_1), .A2(n_105), .B1(n_496), .B2(n_498), .Y(n_495) );
AOI22xp33_ASAP7_75t_SL g646 ( .A1(n_2), .A2(n_252), .B1(n_455), .B2(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_3), .A2(n_256), .B1(n_409), .B2(n_815), .Y(n_814) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_4), .A2(n_38), .B1(n_740), .B2(n_753), .C(n_754), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_5), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_6), .B(n_525), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_7), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_8), .B(n_440), .Y(n_668) );
AOI22xp5_ASAP7_75t_SL g456 ( .A1(n_9), .A2(n_59), .B1(n_457), .B2(n_459), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_10), .A2(n_22), .B1(n_417), .B2(n_418), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_11), .A2(n_168), .B1(n_309), .B2(n_653), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_12), .A2(n_74), .B1(n_314), .B2(n_320), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_13), .A2(n_267), .B1(n_525), .B2(n_526), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_14), .A2(n_126), .B1(n_403), .B2(n_526), .Y(n_747) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_15), .A2(n_119), .B1(n_309), .B2(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_SL g500 ( .A1(n_16), .A2(n_223), .B1(n_501), .B2(n_502), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_17), .A2(n_143), .B1(n_434), .B2(n_481), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_18), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g768 ( .A1(n_19), .A2(n_228), .B1(n_402), .B2(n_769), .C(n_770), .Y(n_768) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_20), .A2(n_23), .B1(n_753), .B2(n_858), .C(n_860), .Y(n_857) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_21), .A2(n_192), .B1(n_396), .B2(n_559), .Y(n_672) );
INVx1_ASAP7_75t_L g586 ( .A(n_24), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_25), .A2(n_287), .B1(n_383), .B2(n_384), .Y(n_286) );
INVx1_ASAP7_75t_L g384 ( .A(n_25), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_26), .A2(n_264), .B1(n_409), .B2(n_482), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_27), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_28), .A2(n_179), .B1(n_493), .B2(n_504), .Y(n_743) );
AOI22xp5_ASAP7_75t_SL g453 ( .A1(n_29), .A2(n_266), .B1(n_454), .B2(n_455), .Y(n_453) );
AO22x2_ASAP7_75t_L g296 ( .A1(n_30), .A2(n_85), .B1(n_297), .B2(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g793 ( .A(n_30), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_31), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_32), .A2(n_35), .B1(n_374), .B2(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_33), .A2(n_63), .B1(n_652), .B2(n_653), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_34), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_36), .A2(n_79), .B1(n_336), .B2(n_340), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_37), .A2(n_197), .B1(n_613), .B2(n_614), .Y(n_612) );
AOI22xp5_ASAP7_75t_SL g446 ( .A1(n_39), .A2(n_140), .B1(n_415), .B2(n_447), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_40), .A2(n_261), .B1(n_309), .B2(n_532), .Y(n_531) );
AO22x1_ASAP7_75t_L g589 ( .A1(n_41), .A2(n_590), .B1(n_619), .B2(n_620), .Y(n_589) );
INVx1_ASAP7_75t_L g619 ( .A(n_41), .Y(n_619) );
AOI222xp33_ASAP7_75t_L g420 ( .A1(n_42), .A2(n_128), .B1(n_198), .B2(n_421), .C1(n_422), .C2(n_424), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_43), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_44), .A2(n_227), .B1(n_391), .B2(n_617), .Y(n_616) );
AO22x2_ASAP7_75t_L g300 ( .A1(n_45), .A2(n_86), .B1(n_297), .B2(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g794 ( .A(n_45), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_46), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_47), .A2(n_200), .B1(n_457), .B2(n_507), .Y(n_733) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_48), .A2(n_208), .B1(n_410), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_49), .A2(n_99), .B1(n_340), .B2(n_613), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_50), .A2(n_67), .B1(n_409), .B2(n_522), .Y(n_748) );
AOI222xp33_ASAP7_75t_L g749 ( .A1(n_51), .A2(n_160), .B1(n_218), .B2(n_373), .C1(n_517), .C2(n_695), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_52), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g853 ( .A1(n_53), .A2(n_269), .B1(n_705), .B2(n_740), .C(n_854), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_54), .Y(n_472) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_55), .A2(n_81), .B1(n_642), .B2(n_643), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_56), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_57), .A2(n_242), .B1(n_413), .B2(n_415), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_58), .A2(n_257), .B1(n_610), .B2(n_611), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_60), .A2(n_630), .B1(n_631), .B2(n_655), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_60), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_61), .A2(n_137), .B1(n_407), .B2(n_409), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_62), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_64), .A2(n_204), .B1(n_493), .B2(n_707), .Y(n_809) );
INVx1_ASAP7_75t_L g861 ( .A(n_65), .Y(n_861) );
AOI22xp33_ASAP7_75t_SL g700 ( .A1(n_66), .A2(n_130), .B1(n_415), .B2(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_68), .A2(n_191), .B1(n_316), .B2(n_559), .Y(n_558) );
AOI222xp33_ASAP7_75t_L g774 ( .A1(n_69), .A2(n_90), .B1(n_155), .B2(n_434), .C1(n_518), .C2(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_70), .B(n_403), .Y(n_553) );
AOI22xp33_ASAP7_75t_SL g702 ( .A1(n_71), .A2(n_115), .B1(n_451), .B2(n_676), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_72), .A2(n_129), .B1(n_396), .B2(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_73), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_75), .A2(n_127), .B1(n_705), .B2(n_761), .C(n_762), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g442 ( .A1(n_76), .A2(n_254), .B1(n_443), .B2(n_444), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_77), .A2(n_158), .B1(n_546), .B2(n_547), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_78), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_80), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_82), .A2(n_217), .B1(n_314), .B2(n_507), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_83), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_84), .A2(n_151), .B1(n_498), .B2(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_87), .A2(n_183), .B1(n_314), .B2(n_530), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_88), .B(n_402), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_89), .Y(n_851) );
INVx1_ASAP7_75t_L g277 ( .A(n_91), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_92), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_93), .A2(n_144), .B1(n_374), .B2(n_423), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_94), .A2(n_189), .B1(n_546), .B2(n_547), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_95), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_96), .A2(n_112), .B1(n_391), .B2(n_392), .Y(n_390) );
INVx1_ASAP7_75t_L g274 ( .A(n_97), .Y(n_274) );
INVx1_ASAP7_75t_L g863 ( .A(n_98), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_100), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_101), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_102), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_103), .A2(n_123), .B1(n_392), .B2(n_504), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_104), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_106), .Y(n_856) );
OA22x2_ASAP7_75t_L g683 ( .A1(n_107), .A2(n_684), .B1(n_685), .B2(n_686), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_107), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_108), .A2(n_145), .B1(n_340), .B2(n_417), .Y(n_741) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_109), .A2(n_110), .B1(n_336), .B2(n_498), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_111), .A2(n_133), .B1(n_407), .B2(n_476), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_113), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_114), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_116), .A2(n_125), .B1(n_392), .B2(n_740), .Y(n_739) );
AOI22xp33_ASAP7_75t_SL g433 ( .A1(n_117), .A2(n_173), .B1(n_374), .B2(n_434), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_118), .A2(n_163), .B1(n_394), .B2(n_396), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_120), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_121), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_122), .A2(n_222), .B1(n_310), .B2(n_450), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_124), .Y(n_572) );
XOR2x2_ASAP7_75t_L g712 ( .A(n_131), .B(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_132), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_134), .A2(n_220), .B1(n_504), .B2(n_507), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_135), .Y(n_486) );
XNOR2x2_ASAP7_75t_L g736 ( .A(n_136), .B(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_138), .Y(n_432) );
INVx2_ASAP7_75t_L g278 ( .A(n_139), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_141), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_142), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_146), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_147), .Y(n_823) );
INVx1_ASAP7_75t_L g835 ( .A(n_148), .Y(n_835) );
AO22x1_ASAP7_75t_L g837 ( .A1(n_148), .A2(n_835), .B1(n_838), .B2(n_864), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_149), .A2(n_224), .B1(n_530), .B2(n_566), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_150), .Y(n_842) );
INVx1_ASAP7_75t_L g678 ( .A(n_152), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_153), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_154), .B(n_440), .Y(n_554) );
AND2x6_ASAP7_75t_L g273 ( .A(n_156), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_156), .Y(n_787) );
AO22x2_ASAP7_75t_L g304 ( .A1(n_157), .A2(n_233), .B1(n_297), .B2(n_301), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_159), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_161), .A2(n_797), .B1(n_824), .B2(n_825), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_161), .Y(n_824) );
AOI22xp5_ASAP7_75t_SL g448 ( .A1(n_162), .A2(n_231), .B1(n_449), .B2(n_451), .Y(n_448) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_164), .A2(n_271), .B(n_279), .C(n_795), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_165), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_166), .A2(n_243), .B1(n_454), .B2(n_705), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_167), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_169), .A2(n_253), .B1(n_444), .B2(n_522), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_170), .B(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_171), .A2(n_216), .B1(n_356), .B2(n_407), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_172), .B(n_402), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_174), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_175), .A2(n_250), .B1(n_419), .B2(n_496), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_176), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_177), .B(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_178), .A2(n_232), .B1(n_391), .B2(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_180), .A2(n_193), .B1(n_532), .B2(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_181), .B(n_373), .Y(n_849) );
AO22x2_ASAP7_75t_L g306 ( .A1(n_182), .A2(n_245), .B1(n_297), .B2(n_298), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_184), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_185), .Y(n_595) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_186), .A2(n_213), .B1(n_373), .B2(n_423), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_187), .B(n_639), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_188), .A2(n_229), .B1(n_316), .B2(n_501), .Y(n_673) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_190), .A2(n_210), .B1(n_517), .B2(n_518), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_194), .Y(n_398) );
INVx1_ASAP7_75t_L g460 ( .A(n_195), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_196), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_199), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_201), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_202), .A2(n_225), .B1(n_459), .B2(n_745), .Y(n_744) );
AO22x1_ASAP7_75t_L g750 ( .A1(n_203), .A2(n_751), .B1(n_776), .B2(n_777), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_203), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_205), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_206), .A2(n_262), .B1(n_417), .B2(n_498), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_207), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_209), .Y(n_846) );
AOI22xp33_ASAP7_75t_SL g654 ( .A1(n_211), .A2(n_212), .B1(n_459), .B2(n_532), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_214), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_215), .Y(n_813) );
OA22x2_ASAP7_75t_L g509 ( .A1(n_219), .A2(n_510), .B1(n_511), .B2(n_536), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_219), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_221), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_226), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_230), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_233), .B(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_234), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_235), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_236), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_237), .Y(n_802) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_238), .A2(n_268), .B1(n_292), .B2(n_506), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_239), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_240), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_244), .Y(n_550) );
INVx1_ASAP7_75t_L g790 ( .A(n_245), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g855 ( .A(n_246), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_247), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_248), .B(n_423), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_249), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_251), .B(n_402), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_255), .Y(n_471) );
INVx1_ASAP7_75t_L g297 ( .A(n_258), .Y(n_297) );
INVx1_ASAP7_75t_L g299 ( .A(n_258), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_259), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_260), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_263), .B(n_438), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_265), .Y(n_605) );
INVx2_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_274), .Y(n_786) );
OA21x2_ASAP7_75t_L g833 ( .A1(n_275), .A2(n_785), .B(n_834), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_623), .B1(n_780), .B2(n_781), .C(n_782), .Y(n_279) );
INVx1_ASAP7_75t_L g780 ( .A(n_280), .Y(n_780) );
AOI22xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_589), .B1(n_621), .B2(n_622), .Y(n_280) );
INVx1_ASAP7_75t_L g621 ( .A(n_281), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_539), .B2(n_588), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI22xp5_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_285), .B1(n_462), .B2(n_463), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_385), .B1(n_386), .B2(n_461), .Y(n_285) );
INVx2_ASAP7_75t_L g461 ( .A(n_286), .Y(n_461) );
INVx1_ASAP7_75t_L g383 ( .A(n_287), .Y(n_383) );
AND2x2_ASAP7_75t_SL g287 ( .A(n_288), .B(n_343), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_325), .Y(n_288) );
OAI221xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_307), .B1(n_308), .B2(n_312), .C(n_313), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g391 ( .A(n_291), .Y(n_391) );
INVx5_ASAP7_75t_SL g501 ( .A(n_291), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_291), .A2(n_414), .B1(n_569), .B2(n_570), .Y(n_568) );
INVx4_ASAP7_75t_L g745 ( .A(n_291), .Y(n_745) );
INVx11_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx11_ASAP7_75t_L g458 ( .A(n_292), .Y(n_458) );
AND2x6_ASAP7_75t_L g292 ( .A(n_293), .B(n_302), .Y(n_292) );
AND2x4_ASAP7_75t_L g405 ( .A(n_293), .B(n_328), .Y(n_405) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g348 ( .A(n_294), .B(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_300), .Y(n_294) );
AND2x2_ASAP7_75t_L g311 ( .A(n_295), .B(n_300), .Y(n_311) );
AND2x2_ASAP7_75t_L g318 ( .A(n_295), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g359 ( .A(n_296), .B(n_304), .Y(n_359) );
AND2x2_ASAP7_75t_L g363 ( .A(n_296), .B(n_300), .Y(n_363) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g301 ( .A(n_299), .Y(n_301) );
INVx2_ASAP7_75t_L g319 ( .A(n_300), .Y(n_319) );
INVx1_ASAP7_75t_L g342 ( .A(n_300), .Y(n_342) );
AND2x4_ASAP7_75t_L g310 ( .A(n_302), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g317 ( .A(n_302), .B(n_318), .Y(n_317) );
AND2x6_ASAP7_75t_L g362 ( .A(n_302), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
AND2x2_ASAP7_75t_L g328 ( .A(n_303), .B(n_306), .Y(n_328) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g323 ( .A(n_304), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_304), .B(n_306), .Y(n_333) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g324 ( .A(n_306), .Y(n_324) );
INVx1_ASAP7_75t_L g358 ( .A(n_306), .Y(n_358) );
INVx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx6_ASAP7_75t_L g414 ( .A(n_310), .Y(n_414) );
BUFx3_ASAP7_75t_L g494 ( .A(n_310), .Y(n_494) );
BUFx3_ASAP7_75t_L g707 ( .A(n_310), .Y(n_707) );
AND2x2_ASAP7_75t_L g339 ( .A(n_311), .B(n_323), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_311), .B(n_328), .Y(n_352) );
AND2x6_ASAP7_75t_L g440 ( .A(n_311), .B(n_328), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g765 ( .A(n_311), .B(n_323), .Y(n_765) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_315), .A2(n_572), .B1(n_573), .B2(n_574), .Y(n_571) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx3_ASAP7_75t_L g493 ( .A(n_316), .Y(n_493) );
BUFx3_ASAP7_75t_L g610 ( .A(n_316), .Y(n_610) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_316), .Y(n_652) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g395 ( .A(n_317), .Y(n_395) );
BUFx2_ASAP7_75t_SL g447 ( .A(n_317), .Y(n_447) );
BUFx2_ASAP7_75t_SL g753 ( .A(n_317), .Y(n_753) );
AND2x2_ASAP7_75t_L g322 ( .A(n_318), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g327 ( .A(n_318), .B(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g331 ( .A(n_318), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_318), .B(n_323), .Y(n_576) );
AND2x2_ASAP7_75t_L g357 ( .A(n_319), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g368 ( .A(n_319), .Y(n_368) );
BUFx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g396 ( .A(n_322), .Y(n_396) );
BUFx3_ASAP7_75t_L g454 ( .A(n_322), .Y(n_454) );
BUFx3_ASAP7_75t_L g506 ( .A(n_322), .Y(n_506) );
INVx1_ASAP7_75t_L g382 ( .A(n_324), .Y(n_382) );
OAI221xp5_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_329), .B1(n_330), .B2(n_334), .C(n_335), .Y(n_325) );
INVx1_ASAP7_75t_L g611 ( .A(n_326), .Y(n_611) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx3_ASAP7_75t_L g415 ( .A(n_327), .Y(n_415) );
BUFx3_ASAP7_75t_L g508 ( .A(n_327), .Y(n_508) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_327), .Y(n_546) );
BUFx3_ASAP7_75t_L g566 ( .A(n_327), .Y(n_566) );
INVx1_ASAP7_75t_L g349 ( .A(n_328), .Y(n_349) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx3_ASAP7_75t_L g392 ( .A(n_331), .Y(n_392) );
BUFx2_ASAP7_75t_L g455 ( .A(n_331), .Y(n_455) );
BUFx2_ASAP7_75t_SL g502 ( .A(n_331), .Y(n_502) );
BUFx2_ASAP7_75t_SL g530 ( .A(n_331), .Y(n_530) );
BUFx3_ASAP7_75t_L g559 ( .A(n_331), .Y(n_559) );
BUFx3_ASAP7_75t_L g705 ( .A(n_331), .Y(n_705) );
AND2x2_ASAP7_75t_L g547 ( .A(n_332), .B(n_368), .Y(n_547) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x6_ASAP7_75t_L g341 ( .A(n_333), .B(n_342), .Y(n_341) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx3_ASAP7_75t_L g417 ( .A(n_338), .Y(n_417) );
INVx4_ASAP7_75t_L g450 ( .A(n_338), .Y(n_450) );
INVx5_ASAP7_75t_L g676 ( .A(n_338), .Y(n_676) );
INVx2_ASAP7_75t_L g805 ( .A(n_338), .Y(n_805) );
INVx8_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx6_ASAP7_75t_SL g419 ( .A(n_341), .Y(n_419) );
INVx1_ASAP7_75t_SL g498 ( .A(n_341), .Y(n_498) );
INVx1_ASAP7_75t_L g408 ( .A(n_342), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_353), .C(n_370), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B1(n_350), .B2(n_351), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_346), .A2(n_841), .B1(n_842), .B2(n_843), .Y(n_840) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g594 ( .A(n_347), .Y(n_594) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_348), .Y(n_470) );
BUFx3_ASAP7_75t_L g690 ( .A(n_348), .Y(n_690) );
OAI22xp5_ASAP7_75t_SL g469 ( .A1(n_351), .A2(n_470), .B1(n_471), .B2(n_472), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_351), .A2(n_689), .B1(n_690), .B2(n_691), .Y(n_688) );
INVx2_ASAP7_75t_L g719 ( .A(n_351), .Y(n_719) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g400 ( .A(n_352), .Y(n_400) );
OAI222xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_360), .B1(n_361), .B2(n_364), .C1(n_365), .C2(n_369), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx4f_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_356), .Y(n_423) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_356), .Y(n_476) );
BUFx2_ASAP7_75t_L g517 ( .A(n_356), .Y(n_517) );
BUFx6f_ASAP7_75t_L g818 ( .A(n_356), .Y(n_818) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g376 ( .A(n_358), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_359), .B(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g375 ( .A(n_359), .B(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g407 ( .A(n_359), .B(n_408), .Y(n_407) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_361), .A2(n_662), .B(n_663), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g720 ( .A1(n_361), .A2(n_602), .B1(n_721), .B2(n_722), .C(n_723), .Y(n_720) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_362), .Y(n_421) );
INVx4_ASAP7_75t_L g431 ( .A(n_362), .Y(n_431) );
INVx2_ASAP7_75t_SL g478 ( .A(n_362), .Y(n_478) );
INVx2_ASAP7_75t_L g514 ( .A(n_362), .Y(n_514) );
BUFx3_ASAP7_75t_L g695 ( .A(n_362), .Y(n_695) );
INVx1_ASAP7_75t_L g380 ( .A(n_363), .Y(n_380) );
AND2x4_ASAP7_75t_L g410 ( .A(n_363), .B(n_382), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_365), .A2(n_487), .B1(n_851), .B2(n_852), .Y(n_850) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx4_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g485 ( .A(n_367), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_367), .A2(n_379), .B1(n_697), .B2(n_698), .Y(n_696) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_367), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_377), .B2(n_378), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx4f_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g425 ( .A(n_374), .Y(n_425) );
BUFx12f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_375), .Y(n_482) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_375), .Y(n_519) );
BUFx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_379), .Y(n_488) );
OR2x6_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
XNOR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_427), .Y(n_386) );
XOR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_426), .Y(n_387) );
NAND4xp75_ASAP7_75t_L g388 ( .A(n_389), .B(n_397), .C(n_411), .D(n_420), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_393), .Y(n_389) );
INVx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g701 ( .A(n_395), .Y(n_701) );
OA211x2_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B(n_401), .C(n_406), .Y(n_397) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g596 ( .A(n_400), .Y(n_596) );
INVx1_ASAP7_75t_SL g843 ( .A(n_400), .Y(n_843) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx5_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g525 ( .A(n_404), .Y(n_525) );
INVx2_ASAP7_75t_L g667 ( .A(n_404), .Y(n_667) );
INVx4_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g443 ( .A(n_407), .Y(n_443) );
INVx1_ASAP7_75t_L g523 ( .A(n_407), .Y(n_523) );
BUFx2_ASAP7_75t_L g815 ( .A(n_407), .Y(n_815) );
INVx1_ASAP7_75t_SL g644 ( .A(n_409), .Y(n_644) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx2_ASAP7_75t_SL g444 ( .A(n_410), .Y(n_444) );
BUFx3_ASAP7_75t_L g664 ( .A(n_410), .Y(n_664) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_416), .Y(n_411) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g459 ( .A(n_414), .Y(n_459) );
INVx2_ASAP7_75t_L g617 ( .A(n_414), .Y(n_617) );
INVx2_ASAP7_75t_L g757 ( .A(n_414), .Y(n_757) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g451 ( .A(n_419), .Y(n_451) );
BUFx4f_ASAP7_75t_SL g614 ( .A(n_419), .Y(n_614) );
INVx2_ASAP7_75t_SL g600 ( .A(n_421), .Y(n_600) );
INVx2_ASAP7_75t_L g634 ( .A(n_421), .Y(n_634) );
BUFx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx4_ASAP7_75t_L g435 ( .A(n_423), .Y(n_435) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
XOR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_460), .Y(n_427) );
NAND3x1_ASAP7_75t_L g428 ( .A(n_429), .B(n_445), .C(n_452), .Y(n_428) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_436), .Y(n_429) );
OAI21xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_432), .B(n_433), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_431), .A2(n_550), .B(n_551), .Y(n_549) );
OAI21xp5_ASAP7_75t_SL g578 ( .A1(n_431), .A2(n_579), .B(n_580), .Y(n_578) );
INVx4_ASAP7_75t_L g775 ( .A(n_431), .Y(n_775) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_441), .C(n_442), .Y(n_436) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g526 ( .A(n_439), .Y(n_526) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g583 ( .A(n_440), .Y(n_583) );
BUFx2_ASAP7_75t_L g639 ( .A(n_440), .Y(n_639) );
BUFx4f_ASAP7_75t_L g769 ( .A(n_440), .Y(n_769) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g497 ( .A(n_450), .Y(n_497) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_450), .Y(n_613) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g859 ( .A(n_454), .Y(n_859) );
INVx2_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx4_ASAP7_75t_L g532 ( .A(n_458), .Y(n_532) );
INVx3_ASAP7_75t_L g761 ( .A(n_458), .Y(n_761) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_509), .B1(n_537), .B2(n_538), .Y(n_464) );
INVx2_ASAP7_75t_L g537 ( .A(n_465), .Y(n_537) );
XNOR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_490), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .C(n_484), .Y(n_468) );
OAI221xp5_ASAP7_75t_SL g811 ( .A1(n_470), .A2(n_718), .B1(n_812), .B2(n_813), .C(n_814), .Y(n_811) );
OAI222xp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_477), .B1(n_478), .B2(n_479), .C1(n_480), .C2(n_483), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_SL g847 ( .A(n_475), .Y(n_847) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx4f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI22xp5_ASAP7_75t_SL g484 ( .A1(n_485), .A2(n_486), .B1(n_487), .B2(n_489), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_485), .A2(n_487), .B1(n_605), .B2(n_606), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_485), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_487), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_724) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g773 ( .A(n_488), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_499), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_495), .Y(n_491) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_503), .Y(n_499) );
INVx1_ASAP7_75t_L g801 ( .A(n_502), .Y(n_801) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx4f_ASAP7_75t_SL g653 ( .A(n_506), .Y(n_653) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g538 ( .A(n_509), .Y(n_538) );
INVx2_ASAP7_75t_L g536 ( .A(n_511), .Y(n_536) );
NAND2x1_ASAP7_75t_L g511 ( .A(n_512), .B(n_527), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_520), .Y(n_512) );
OAI21xp5_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_515), .B(n_516), .Y(n_513) );
INVx1_ASAP7_75t_L g598 ( .A(n_517), .Y(n_598) );
INVx2_ASAP7_75t_L g602 ( .A(n_518), .Y(n_602) );
BUFx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx2_ASAP7_75t_L g822 ( .A(n_519), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_524), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g642 ( .A(n_523), .Y(n_642) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx1_ASAP7_75t_L g862 ( .A(n_532), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g588 ( .A(n_539), .Y(n_588) );
OA22x2_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B1(n_561), .B2(n_587), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_540), .A2(n_541), .B1(n_682), .B2(n_683), .Y(n_681) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
XOR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_560), .Y(n_541) );
NAND3x1_ASAP7_75t_SL g542 ( .A(n_543), .B(n_548), .C(n_556), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
INVx4_ASAP7_75t_L g648 ( .A(n_546), .Y(n_648) );
NOR2x1_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .C(n_555), .Y(n_552) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g587 ( .A(n_561), .Y(n_587) );
XOR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_586), .Y(n_561) );
AND2x2_ASAP7_75t_SL g562 ( .A(n_563), .B(n_577), .Y(n_562) );
NOR3xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .C(n_571), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
BUFx2_ASAP7_75t_L g808 ( .A(n_566), .Y(n_808) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g759 ( .A(n_575), .Y(n_759) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .C(n_585), .Y(n_581) );
INVx1_ASAP7_75t_L g622 ( .A(n_589), .Y(n_622) );
INVx1_ASAP7_75t_SL g620 ( .A(n_590), .Y(n_620) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_607), .Y(n_590) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_597), .C(n_604), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_594), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_715) );
OAI222xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_600), .B2(n_601), .C1(n_602), .C2(n_603), .Y(n_597) );
OAI222xp33_ASAP7_75t_L g816 ( .A1(n_600), .A2(n_817), .B1(n_819), .B2(n_820), .C1(n_821), .C2(n_823), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_615), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_612), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_614), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g781 ( .A(n_623), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B1(n_680), .B2(n_779), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_627), .B1(n_656), .B2(n_679), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g655 ( .A(n_631), .Y(n_655) );
NAND3x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_645), .C(n_650), .Y(n_631) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_633), .B(n_637), .Y(n_632) );
OAI21xp5_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_635), .B(n_636), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .C(n_641), .Y(n_637) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_649), .Y(n_645) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx4_ASAP7_75t_L g740 ( .A(n_648), .Y(n_740) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g679 ( .A(n_656), .Y(n_679) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
XOR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_678), .Y(n_658) );
NAND2x1p5_ASAP7_75t_L g659 ( .A(n_660), .B(n_670), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_665), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .C(n_669), .Y(n_665) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_674), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx1_ASAP7_75t_L g779 ( .A(n_680), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_708), .B1(n_709), .B2(n_778), .Y(n_680) );
CKINVDCx14_ASAP7_75t_R g778 ( .A(n_681), .Y(n_778) );
INVx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND3x1_ASAP7_75t_L g686 ( .A(n_687), .B(n_699), .C(n_703), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_692), .C(n_696), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx3_ASAP7_75t_L g845 ( .A(n_695), .Y(n_845) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
XOR2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_750), .Y(n_709) );
OAI22xp5_ASAP7_75t_SL g710 ( .A1(n_711), .A2(n_712), .B1(n_735), .B2(n_736), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_728), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_720), .C(n_724), .Y(n_714) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_732), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND4xp75_ASAP7_75t_L g737 ( .A(n_738), .B(n_742), .C(n_746), .D(n_749), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .Y(n_738) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
AND2x2_ASAP7_75t_SL g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g777 ( .A(n_751), .Y(n_777) );
AND4x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_760), .C(n_768), .D(n_774), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B1(n_758), .B2(n_759), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_756), .A2(n_861), .B1(n_862), .B2(n_863), .Y(n_860) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OAI221xp5_ASAP7_75t_SL g799 ( .A1(n_759), .A2(n_800), .B1(n_801), .B2(n_802), .C(n_803), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B1(n_766), .B2(n_767), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_764), .A2(n_767), .B1(n_855), .B2(n_856), .Y(n_854) );
BUFx2_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
NOR2x1_ASAP7_75t_L g783 ( .A(n_784), .B(n_788), .Y(n_783) );
OR2x2_ASAP7_75t_SL g867 ( .A(n_784), .B(n_789), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_787), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_785), .Y(n_827) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_786), .B(n_830), .Y(n_834) );
CKINVDCx16_ASAP7_75t_R g830 ( .A(n_787), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
OAI322xp33_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_826), .A3(n_828), .B1(n_831), .B2(n_835), .C1(n_836), .C2(n_865), .Y(n_795) );
INVx1_ASAP7_75t_L g825 ( .A(n_797), .Y(n_825) );
AND2x2_ASAP7_75t_SL g797 ( .A(n_798), .B(n_810), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_806), .Y(n_798) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_809), .Y(n_806) );
NOR2xp33_ASAP7_75t_SL g810 ( .A(n_811), .B(n_816), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
INVxp67_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g864 ( .A(n_838), .Y(n_864) );
AND3x1_ASAP7_75t_L g838 ( .A(n_839), .B(n_853), .C(n_857), .Y(n_838) );
NOR3xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_844), .C(n_850), .Y(n_839) );
OAI221xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B1(n_847), .B2(n_848), .C(n_849), .Y(n_844) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_866), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_867), .Y(n_866) );
endmodule