module fake_jpeg_1635_n_310 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVxp33_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_7),
.B(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_15),
.B(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_9),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_52),
.B(n_54),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_11),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_11),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_62),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_7),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_59),
.B(n_66),
.Y(n_107)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_60),
.Y(n_136)
);

NAND2x1_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_0),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_85),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_30),
.B(n_12),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_26),
.B(n_4),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_68),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_20),
.A2(n_13),
.B(n_15),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_67),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_3),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_26),
.B(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_76),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_47),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_74),
.Y(n_152)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_13),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_81),
.Y(n_132)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_14),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_83),
.B(n_87),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_28),
.B(n_16),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_89),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_92),
.Y(n_117)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_101),
.B1(n_22),
.B2(n_43),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_23),
.B(n_0),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_94),
.Y(n_141)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_99),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_96),
.B(n_97),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_28),
.B(n_1),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_34),
.Y(n_105)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_23),
.B(n_1),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_29),
.Y(n_151)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_135),
.Y(n_172)
);

BUFx4f_ASAP7_75t_SL g163 ( 
.A(n_106),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_41),
.B1(n_40),
.B2(n_27),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_120),
.B1(n_121),
.B2(n_137),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_46),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_126),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_41),
.B1(n_40),
.B2(n_27),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_74),
.A2(n_46),
.B1(n_36),
.B2(n_33),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_61),
.B(n_33),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_62),
.A2(n_34),
.B1(n_38),
.B2(n_44),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_129),
.A2(n_130),
.B1(n_142),
.B2(n_143),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_92),
.B1(n_98),
.B2(n_96),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_75),
.B(n_38),
.C(n_44),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_57),
.A2(n_36),
.B1(n_38),
.B2(n_44),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_94),
.A2(n_78),
.B1(n_82),
.B2(n_70),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_51),
.A2(n_29),
.B1(n_21),
.B2(n_2),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_53),
.A2(n_29),
.B1(n_21),
.B2(n_1),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_71),
.B1(n_80),
.B2(n_91),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_60),
.A2(n_29),
.B(n_56),
.C(n_99),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_153),
.B(n_67),
.C(n_86),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_152),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_95),
.A2(n_29),
.B(n_58),
.C(n_64),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_84),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_84),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_156),
.B(n_169),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_160),
.Y(n_194)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_158),
.Y(n_214)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_117),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_181),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_164),
.Y(n_221)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_126),
.B(n_67),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_167),
.Y(n_196)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_132),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_150),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_171),
.B(n_177),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_123),
.A2(n_153),
.B(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_174),
.Y(n_197)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_104),
.A2(n_115),
.A3(n_123),
.B1(n_141),
.B2(n_105),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_112),
.B(n_149),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_102),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_186),
.Y(n_199)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_131),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g182 ( 
.A(n_122),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_110),
.A2(n_133),
.B1(n_122),
.B2(n_125),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_183),
.A2(n_188),
.B1(n_139),
.B2(n_138),
.Y(n_204)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_127),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_118),
.B(n_127),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_191),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_135),
.A2(n_146),
.B1(n_145),
.B2(n_116),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_129),
.A2(n_130),
.B1(n_146),
.B2(n_116),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_189),
.A2(n_172),
.B1(n_166),
.B2(n_173),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_L g190 ( 
.A1(n_131),
.A2(n_145),
.B1(n_124),
.B2(n_133),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_124),
.B1(n_119),
.B2(n_139),
.Y(n_200)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_136),
.B(n_128),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_167),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_154),
.A2(n_110),
.B1(n_128),
.B2(n_109),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_195),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_204),
.B1(n_210),
.B2(n_190),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_119),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_211),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_174),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_160),
.A2(n_166),
.B1(n_176),
.B2(n_172),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_183),
.B(n_189),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_220),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_176),
.B(n_186),
.Y(n_220)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_163),
.B(n_157),
.C(n_185),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_196),
.B(n_209),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

AOI22x1_ASAP7_75t_SL g224 ( 
.A1(n_197),
.A2(n_167),
.B1(n_163),
.B2(n_159),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_224),
.A2(n_225),
.B(n_238),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_211),
.B1(n_194),
.B2(n_199),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_230),
.B1(n_243),
.B2(n_193),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_180),
.C(n_170),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_228),
.C(n_207),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_161),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_205),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_234),
.Y(n_244)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_205),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_163),
.B1(n_157),
.B2(n_175),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_236),
.A2(n_201),
.B1(n_209),
.B2(n_200),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_194),
.A2(n_191),
.B(n_182),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_240),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_212),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_168),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_242),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_158),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_194),
.A2(n_157),
.B1(n_164),
.B2(n_165),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_248),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_196),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_253),
.C(n_258),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_255),
.B1(n_225),
.B2(n_231),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_203),
.A3(n_207),
.B1(n_193),
.B2(n_221),
.C1(n_198),
.C2(n_218),
.Y(n_251)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_203),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_236),
.B1(n_230),
.B2(n_224),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_271),
.B1(n_256),
.B2(n_250),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_264),
.A2(n_269),
.B1(n_245),
.B2(n_244),
.Y(n_274)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_272),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_227),
.C(n_234),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_270),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_243),
.B1(n_238),
.B2(n_237),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_229),
.C(n_241),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_248),
.A2(n_222),
.B1(n_233),
.B2(n_235),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_233),
.B(n_237),
.Y(n_272)
);

AOI321xp33_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_244),
.A3(n_253),
.B1(n_257),
.B2(n_252),
.C(n_267),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_275),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_265),
.B1(n_223),
.B2(n_218),
.Y(n_290)
);

AOI321xp33_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_253),
.A3(n_252),
.B1(n_256),
.B2(n_246),
.C(n_259),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_268),
.Y(n_278)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_246),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_269),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_260),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_247),
.B1(n_251),
.B2(n_239),
.Y(n_281)
);

AOI321xp33_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_260),
.A3(n_272),
.B1(n_265),
.B2(n_271),
.C(n_264),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_288),
.C(n_221),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_286),
.A2(n_282),
.B(n_277),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_260),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_287),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_262),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_280),
.B(n_281),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_290),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_294),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_202),
.B(n_223),
.C(n_214),
.Y(n_293)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_288),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_289),
.B(n_287),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_290),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_292),
.C(n_285),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_301),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_298),
.B(n_202),
.Y(n_307)
);

O2A1O1Ixp33_ASAP7_75t_SL g306 ( 
.A1(n_305),
.A2(n_300),
.B(n_297),
.C(n_296),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_307),
.B1(n_219),
.B2(n_213),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_219),
.B(n_213),
.C(n_164),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_213),
.Y(n_310)
);


endmodule