module fake_netlist_6_2346_n_4805 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4805);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4805;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_4730;
wire n_801;
wire n_4452;
wire n_3766;
wire n_1613;
wire n_4598;
wire n_1458;
wire n_2576;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_4649;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_4670;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_4620;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_4738;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_700;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_4504;
wire n_3844;
wire n_4395;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4388;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4517;
wire n_4168;
wire n_783;
wire n_2451;
wire n_1738;
wire n_4490;
wire n_2243;
wire n_1575;
wire n_798;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_4686;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_4699;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1930;
wire n_3706;
wire n_2405;
wire n_1743;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_2997;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1238;
wire n_4092;
wire n_4645;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_4755;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_4578;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_4777;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4591;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_4702;
wire n_2291;
wire n_4754;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_1371;
wire n_873;
wire n_2886;
wire n_2974;
wire n_1285;
wire n_3946;
wire n_4213;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_4474;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_4531;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2628;
wire n_3071;
wire n_2313;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1517;
wire n_1867;
wire n_1393;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_4666;
wire n_2470;
wire n_2321;
wire n_4446;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_4417;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_4501;
wire n_3678;
wire n_3440;
wire n_4617;
wire n_4733;
wire n_2129;
wire n_2340;
wire n_4764;
wire n_1261;
wire n_4724;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_4555;
wire n_4743;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_4696;
wire n_4692;
wire n_1572;
wire n_3979;
wire n_658;
wire n_616;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2739;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_3023;
wire n_2510;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_4602;
wire n_2212;
wire n_3929;
wire n_758;
wire n_3048;
wire n_1455;
wire n_3063;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_2418;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_943;
wire n_4060;
wire n_1550;
wire n_4767;
wire n_2703;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_4722;
wire n_4606;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_1094;
wire n_953;
wire n_3737;
wire n_3077;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_539;
wire n_4556;
wire n_3107;
wire n_4563;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_4687;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_4619;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4600;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_4646;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_4255;
wire n_4403;
wire n_3506;
wire n_4729;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_3413;
wire n_1230;
wire n_3850;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_4751;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_4605;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_4549;
wire n_4575;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_2113;
wire n_3871;
wire n_2190;
wire n_1918;
wire n_3603;
wire n_1641;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_4662;
wire n_1843;
wire n_619;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_1909;
wire n_2080;
wire n_813;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_1441;
wire n_606;
wire n_818;
wire n_3373;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_3910;
wire n_1699;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_4507;
wire n_630;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_541;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_4499;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_4677;
wire n_3272;
wire n_4765;
wire n_3193;
wire n_2522;
wire n_792;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_4732;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_2811;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_4372;
wire n_982;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_2832;
wire n_4581;
wire n_4226;
wire n_549;
wire n_1762;
wire n_4641;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2998;
wire n_2831;
wire n_4318;
wire n_4366;
wire n_3446;
wire n_4158;
wire n_4377;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_4259;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_4795;
wire n_3630;
wire n_4698;
wire n_3518;
wire n_4445;
wire n_3824;
wire n_4792;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3842;
wire n_4544;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_4772;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_4477;
wire n_966;
wire n_3888;
wire n_4511;
wire n_2908;
wire n_3168;
wire n_764;
wire n_4468;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_3092;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3492;
wire n_1233;
wire n_3966;
wire n_3895;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_4520;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_4502;
wire n_882;
wire n_4503;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_4375;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_4526;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_4319;
wire n_2434;
wire n_4613;
wire n_3369;
wire n_3419;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_4478;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_4717;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_612;
wire n_2641;
wire n_4585;
wire n_4731;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_4773;
wire n_3933;
wire n_702;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_4467;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_4427;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4386;
wire n_4485;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_4681;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_4523;
wire n_4752;
wire n_1801;
wire n_2347;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_928;
wire n_2092;
wire n_3917;
wire n_1654;
wire n_816;
wire n_4371;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_4552;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2519;
wire n_2319;
wire n_4043;
wire n_4673;
wire n_825;
wire n_4313;
wire n_728;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_4607;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_4510;
wire n_696;
wire n_1515;
wire n_4473;
wire n_961;
wire n_4356;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_4055;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_4362;
wire n_950;
wire n_4248;
wire n_2812;
wire n_4518;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_4589;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_4560;
wire n_590;
wire n_4737;
wire n_4685;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_4675;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_3073;
wire n_2431;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_595;
wire n_627;
wire n_1767;
wire n_3253;
wire n_1779;
wire n_1465;
wire n_3337;
wire n_3431;
wire n_3450;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_4603;
wire n_1391;
wire n_4663;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_1208;
wire n_2775;
wire n_1627;
wire n_1295;
wire n_1164;
wire n_4697;
wire n_2954;
wire n_3477;
wire n_4289;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4288;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_815;
wire n_3953;
wire n_1100;
wire n_4588;
wire n_585;
wire n_4653;
wire n_1487;
wire n_4435;
wire n_2691;
wire n_3614;
wire n_2913;
wire n_3421;
wire n_840;
wire n_874;
wire n_4471;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_4802;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_4728;
wire n_898;
wire n_4385;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_3423;
wire n_2573;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_1932;
wire n_925;
wire n_1101;
wire n_1026;
wire n_2535;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_4191;
wire n_4636;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_4701;
wire n_4651;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_4576;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_4615;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_2897;
wire n_851;
wire n_644;
wire n_682;
wire n_2537;
wire n_847;
wire n_3970;
wire n_4389;
wire n_4483;
wire n_4345;
wire n_2554;
wire n_996;
wire n_532;
wire n_4661;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_791;
wire n_1913;
wire n_4621;
wire n_4216;
wire n_3608;
wire n_837;
wire n_4540;
wire n_4315;
wire n_4664;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2643;
wire n_2590;
wire n_3353;
wire n_3018;
wire n_3150;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_4785;
wire n_3470;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4713;
wire n_4098;
wire n_4021;
wire n_4476;
wire n_765;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_4688;
wire n_3166;
wire n_4753;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_4775;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_4674;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_4481;
wire n_1246;
wire n_4528;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_4475;
wire n_899;
wire n_2012;
wire n_738;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_4669;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_4443;
wire n_3887;
wire n_4634;
wire n_1022;
wire n_614;
wire n_529;
wire n_2307;
wire n_2069;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_4123;
wire n_1431;
wire n_4096;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4587;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_947;
wire n_2936;
wire n_3224;
wire n_4718;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_4525;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_4440;
wire n_4402;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_3557;
wire n_927;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_4541;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4551;
wire n_4264;
wire n_4484;
wire n_2857;
wire n_3693;
wire n_4497;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_4459;
wire n_1299;
wire n_4545;
wire n_2896;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_4627;
wire n_3674;
wire n_2959;
wire n_2494;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_4464;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_4624;
wire n_2837;
wire n_4175;
wire n_4700;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_4659;
wire n_4771;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_4455;
wire n_4453;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_4514;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_4798;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4564;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_2424;
wire n_745;
wire n_1604;
wire n_2296;
wire n_3201;
wire n_1284;
wire n_3633;
wire n_3447;
wire n_4487;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_623;
wire n_1048;
wire n_1398;
wire n_716;
wire n_2354;
wire n_3032;
wire n_3103;
wire n_2682;
wire n_1201;
wire n_884;
wire n_3638;
wire n_4573;
wire n_4592;
wire n_2589;
wire n_4535;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_3393;
wire n_931;
wire n_811;
wire n_683;
wire n_2442;
wire n_1207;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_958;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_880;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_4695;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_4401;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_589;
wire n_4796;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_2966;
wire n_819;
wire n_2294;
wire n_1363;
wire n_3641;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_767;
wire n_2581;
wire n_1314;
wire n_600;
wire n_964;
wire n_2218;
wire n_2788;
wire n_831;
wire n_1837;
wire n_4533;
wire n_4756;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_1410;
wire n_4746;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_4658;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3944;
wire n_3909;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_3582;
wire n_4665;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_4431;
wire n_1602;
wire n_3270;
wire n_1136;
wire n_2421;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_4633;
wire n_4654;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_642;
wire n_1159;
wire n_995;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_4584;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_4430;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_1093;
wire n_4428;
wire n_4597;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3364;
wire n_3323;
wire n_4020;
wire n_4176;
wire n_4489;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_4404;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_4618;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_4679;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_4496;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_4063;
wire n_1679;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_4513;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_4706;
wire n_2648;
wire n_4747;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_4570;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_4410;
wire n_2462;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4056;
wire n_1617;
wire n_4034;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_4622;
wire n_4721;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_4693;
wire n_2928;
wire n_4206;
wire n_4448;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_2289;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_906;
wire n_3663;
wire n_4132;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_4609;
wire n_4438;
wire n_2135;
wire n_3956;
wire n_4707;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_858;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_4355;
wire n_956;
wire n_960;
wire n_3234;
wire n_2276;
wire n_4422;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_4647;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_3870;
wire n_4126;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_4632;
wire n_1429;
wire n_4655;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_4470;
wire n_587;
wire n_3466;
wire n_4801;
wire n_3554;
wire n_1593;
wire n_4546;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_4583;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_4704;
wire n_4714;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_828;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_4509;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_4374;
wire n_2201;
wire n_952;
wire n_725;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_4668;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4635;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3276;
wire n_3250;
wire n_1934;
wire n_3194;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_4582;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_2924;
wire n_807;
wire n_845;
wire n_4761;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_4420;
wire n_4710;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_4574;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_2598;
wire n_1916;
wire n_597;
wire n_1270;
wire n_2549;
wire n_4690;
wire n_1187;
wire n_4405;
wire n_610;
wire n_4234;
wire n_4304;
wire n_4413;
wire n_1403;
wire n_1669;
wire n_4558;
wire n_1852;
wire n_4488;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_4759;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_2302;
wire n_4211;
wire n_4667;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1397;
wire n_1037;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_750;
wire n_1499;
wire n_901;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_4230;
wire n_4656;
wire n_1841;
wire n_4660;
wire n_3839;
wire n_2823;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4637;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_4797;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_710;
wire n_3730;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_4611;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_4610;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_4472;
wire n_1943;
wire n_1216;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_4725;
wire n_4590;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_3132;
wire n_2486;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_3238;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3529;
wire n_2235;
wire n_4515;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_4614;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_2392;
wire n_3424;
wire n_2894;
wire n_1272;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_4565;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4195;
wire n_4159;
wire n_4567;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_782;
wire n_1539;
wire n_4554;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_4586;
wire n_4778;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_4595;
wire n_4626;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_4734;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_662;
wire n_3475;
wire n_4442;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_4434;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_4680;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_4689;
wire n_3845;
wire n_4616;
wire n_1682;
wire n_2017;
wire n_4516;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2046;
wire n_2272;
wire n_3029;
wire n_2200;
wire n_1695;
wire n_4547;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2760;
wire n_1940;
wire n_1979;
wire n_2560;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_4548;
wire n_4643;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_4601;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_3045;
wire n_936;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_4623;
wire n_885;
wire n_896;
wire n_3278;
wire n_2970;
wire n_2167;
wire n_2084;
wire n_2342;
wire n_3676;
wire n_4553;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_4739;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_3050;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_4135;
wire n_2871;
wire n_4209;
wire n_4279;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_4644;
wire n_4790;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_4561;
wire n_804;
wire n_4461;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_959;
wire n_879;
wire n_2310;
wire n_4608;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_4716;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_4757;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_4682;
wire n_3489;
wire n_4571;
wire n_4343;
wire n_2835;
wire n_4715;
wire n_4530;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_4694;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_4672;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2962;
wire n_2727;
wire n_3377;
wire n_4604;
wire n_2939;
wire n_560;
wire n_4782;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_1914;
wire n_1318;
wire n_737;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3932;
wire n_3469;
wire n_3958;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_4519;
wire n_2388;
wire n_3984;
wire n_4774;
wire n_2056;
wire n_790;
wire n_2901;
wire n_2611;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_4524;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_4469;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_4572;
wire n_3207;
wire n_2668;
wire n_672;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_1941;
wire n_3613;
wire n_3483;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_4726;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3855;
wire n_3743;
wire n_1872;
wire n_3091;
wire n_4736;
wire n_4317;
wire n_834;
wire n_4493;
wire n_4723;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_743;
wire n_766;
wire n_3124;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2923;
wire n_2761;
wire n_2885;
wire n_2888;
wire n_2715;
wire n_2671;
wire n_1804;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_4650;
wire n_4788;
wire n_660;
wire n_2062;
wire n_4539;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_4421;
wire n_4719;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_4793;
wire n_2874;
wire n_1200;
wire n_4498;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_4492;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_4799;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_897;
wire n_4789;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_841;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_3216;
wire n_1177;
wire n_3458;
wire n_4203;
wire n_3515;
wire n_1150;
wire n_4505;
wire n_3808;
wire n_1742;
wire n_3190;
wire n_4657;
wire n_4708;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_4512;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_4542;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_4462;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_4450;
wire n_4536;
wire n_4741;
wire n_4543;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4630;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_4550;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_4652;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_4534;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_4408;
wire n_4577;
wire n_1132;
wire n_4748;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_4439;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_4783;
wire n_955;
wire n_739;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_4639;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_3231;
wire n_1554;
wire n_789;
wire n_4083;
wire n_4494;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_2380;
wire n_769;
wire n_4786;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_4480;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_2746;
wire n_2946;
wire n_814;
wire n_4579;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_691;
wire n_535;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_3473;
wire n_1812;
wire n_957;
wire n_1994;
wire n_1652;
wire n_4557;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_4432;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_744;
wire n_971;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_946;
wire n_4593;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_4342;
wire n_4465;
wire n_3622;
wire n_4568;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_4495;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4436;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_4569;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_4559;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_4373;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_4711;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_4740;
wire n_2117;
wire n_2234;
wire n_4631;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_4720;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_2255;
wire n_2112;
wire n_3494;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_3584;
wire n_3486;
wire n_1414;
wire n_4678;
wire n_4086;
wire n_752;
wire n_908;
wire n_2721;
wire n_2649;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_4625;
wire n_4409;
wire n_2744;
wire n_4363;
wire n_4309;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_4521;
wire n_2437;
wire n_2444;
wire n_1215;
wire n_2743;
wire n_839;
wire n_3962;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_4766;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_1537;
wire n_779;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_854;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_870;
wire n_3362;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_904;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4744;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_3802;
wire n_1276;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_2118;
wire n_4266;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3697;
wire n_3643;
wire n_1584;
wire n_771;
wire n_2425;
wire n_924;
wire n_3461;
wire n_3408;
wire n_1582;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3690;
wire n_3468;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_4532;
wire n_1972;
wire n_719;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_4491;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_2666;
wire n_4105;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_4486;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1156;
wire n_1362;
wire n_911;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_4612;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_4787;
wire n_878;
wire n_620;
wire n_3285;
wire n_4208;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_4529;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_4537;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4351;
wire n_4346;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_4779;
wire n_4640;
wire n_3521;
wire n_3233;
wire n_4599;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_4437;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_4769;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_4628;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_4784;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4508;
wire n_4396;
wire n_1763;
wire n_4594;
wire n_1998;
wire n_3066;
wire n_4727;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_4451;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4108;
wire n_1133;
wire n_4460;
wire n_635;
wire n_3374;
wire n_1194;
wire n_4429;
wire n_4506;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_4538;
wire n_2640;
wire n_3695;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_3552;
wire n_941;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_553;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_849;
wire n_3709;
wire n_4684;
wire n_753;
wire n_4091;
wire n_3925;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_4580;
wire n_3330;
wire n_1479;
wire n_4768;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_1675;
wire n_4758;
wire n_4781;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4522;
wire n_4148;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_4057;
wire n_679;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_633;
wire n_1170;
wire n_1629;
wire n_665;
wire n_2221;
wire n_588;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_4447;
wire n_2891;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_4780;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_4763;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_4803;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_4463;
wire n_1417;
wire n_2185;
wire n_2086;
wire n_1242;
wire n_2927;
wire n_3673;
wire n_4750;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_4648;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_640;
wire n_1322;
wire n_4129;
wire n_4457;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_4804;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_4794;
wire n_722;
wire n_4500;
wire n_862;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_4039;
wire n_4745;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4566;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_4275;
wire n_4482;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_4426;
wire n_531;
wire n_827;
wire n_2912;
wire n_4703;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_4449;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_4762;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_4030;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g529 ( 
.A(n_32),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_268),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_343),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_485),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_265),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_498),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_224),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_401),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_133),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_136),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_474),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_156),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_489),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_29),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_290),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_167),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_407),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_29),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_256),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_108),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_225),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_343),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_517),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_95),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_450),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_203),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_231),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_86),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_525),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_298),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_24),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_23),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_16),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_470),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_194),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_229),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_275),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_437),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_195),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_286),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_211),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_442),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_514),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_245),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_308),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_136),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_416),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_403),
.Y(n_576)
);

CKINVDCx14_ASAP7_75t_R g577 ( 
.A(n_476),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_198),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_18),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_318),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_505),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_504),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_293),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_288),
.Y(n_584)
);

CKINVDCx14_ASAP7_75t_R g585 ( 
.A(n_518),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_101),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_477),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_49),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_252),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_363),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_28),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_102),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_365),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_22),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_521),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_175),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_18),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_208),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_5),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_184),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_244),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_138),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_506),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_324),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_173),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_54),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_397),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_47),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_111),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_510),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_344),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_107),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_512),
.Y(n_613)
);

BUFx8_ASAP7_75t_SL g614 ( 
.A(n_79),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_97),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_511),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_153),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_178),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_4),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_360),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_184),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_216),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_439),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_379),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_347),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_55),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_507),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_71),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_76),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_106),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_482),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_312),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_492),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_524),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_420),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_197),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_51),
.Y(n_637)
);

BUFx5_ASAP7_75t_L g638 ( 
.A(n_47),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_86),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_253),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_74),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_226),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_500),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_491),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_175),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_391),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_357),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_394),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_208),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_446),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_27),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_278),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_275),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_372),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_487),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_25),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_250),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_378),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_519),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_308),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_259),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_494),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_49),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_358),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_37),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_125),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_123),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_342),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_305),
.Y(n_669)
);

BUFx2_ASAP7_75t_R g670 ( 
.A(n_270),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_88),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_19),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_80),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_255),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_303),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_364),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_42),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_367),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_120),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_53),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_444),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_438),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_118),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_279),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_192),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_32),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_111),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_471),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_391),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_131),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_390),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_227),
.Y(n_692)
);

CKINVDCx16_ASAP7_75t_R g693 ( 
.A(n_210),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_318),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_453),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_488),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_483),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_144),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_139),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_481),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_89),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_245),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_351),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_189),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_145),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_1),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_99),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_134),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_69),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_347),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_456),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_122),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_290),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_424),
.Y(n_714)
);

BUFx5_ASAP7_75t_L g715 ( 
.A(n_316),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_193),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_316),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_148),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_164),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_195),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_145),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_371),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_178),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_345),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_50),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_406),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_499),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_231),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_325),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_21),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_198),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_144),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_335),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_56),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_70),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_98),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_37),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_221),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_272),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_314),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_508),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_352),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_138),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_200),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_171),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_262),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_143),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_25),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_397),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_303),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_281),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_192),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_122),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_79),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_4),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_263),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_390),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_486),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_354),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_99),
.Y(n_760)
);

BUFx5_ASAP7_75t_L g761 ( 
.A(n_526),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_377),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_520),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_244),
.Y(n_764)
);

BUFx10_ASAP7_75t_L g765 ( 
.A(n_409),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_172),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_243),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_152),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_165),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_9),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_256),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_473),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_186),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_190),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_105),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_430),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_313),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_309),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_9),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_232),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_356),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_353),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_207),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_132),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_55),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_22),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_404),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_211),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_92),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_327),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_445),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_87),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_385),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_296),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_479),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_417),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_6),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_151),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_513),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_385),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_12),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_480),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_228),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_288),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_181),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_104),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_395),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_254),
.Y(n_808)
);

BUFx5_ASAP7_75t_L g809 ( 
.A(n_312),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_24),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_6),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_88),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_96),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_286),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_281),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_361),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_85),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_139),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_91),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_493),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_168),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_207),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_392),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_412),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_394),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_467),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_527),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_10),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_509),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_135),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_300),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_432),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_159),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_17),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_176),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_388),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_324),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_58),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_23),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_147),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_177),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_190),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_515),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_249),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_282),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_100),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_314),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_75),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_153),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_45),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_325),
.Y(n_851)
);

CKINVDCx16_ASAP7_75t_R g852 ( 
.A(n_326),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_50),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_496),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_38),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_516),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_60),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_185),
.Y(n_858)
);

BUFx10_ASAP7_75t_L g859 ( 
.A(n_215),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_415),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_224),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_151),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_272),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_371),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_183),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_152),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_451),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_395),
.Y(n_868)
);

BUFx8_ASAP7_75t_SL g869 ( 
.A(n_21),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_354),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_337),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_221),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_377),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_7),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_484),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_240),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_114),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_117),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_52),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_309),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_76),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_118),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_276),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_269),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_393),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_497),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_396),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_388),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_91),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_234),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_141),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_130),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_523),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_502),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_361),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_522),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_133),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_202),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_113),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_248),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_154),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_478),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_163),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_61),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_93),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_154),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_181),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_271),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_356),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_204),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_253),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_501),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_26),
.Y(n_913)
);

BUFx5_ASAP7_75t_L g914 ( 
.A(n_287),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_276),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_402),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_115),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_243),
.Y(n_918)
);

CKINVDCx16_ASAP7_75t_R g919 ( 
.A(n_367),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_328),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_503),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_366),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_121),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_234),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_358),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_495),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_301),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_172),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_296),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_218),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_289),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_39),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_74),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_201),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_398),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_213),
.Y(n_936)
);

INVxp33_ASAP7_75t_R g937 ( 
.A(n_251),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_372),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_166),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_121),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_43),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_36),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_387),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_490),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_257),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_163),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_472),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_528),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_475),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_93),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_68),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_594),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_638),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_638),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_638),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_638),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_638),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_638),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_553),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_638),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_638),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_594),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_610),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_695),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_638),
.Y(n_965)
);

INVxp33_ASAP7_75t_SL g966 ( 
.A(n_649),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_680),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_614),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_715),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_680),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_715),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_715),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_613),
.Y(n_973)
);

BUFx10_ASAP7_75t_L g974 ( 
.A(n_807),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_715),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_715),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_715),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_696),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_715),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_715),
.Y(n_980)
);

INVxp33_ASAP7_75t_L g981 ( 
.A(n_877),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_697),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_715),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_758),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_809),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_809),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_809),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_809),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_809),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_869),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_809),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_809),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_809),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_809),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_689),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_947),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_914),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_914),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_914),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_914),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_914),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_914),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_693),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_914),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_914),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_689),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_914),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_773),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_947),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_537),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_537),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_537),
.Y(n_1012)
);

CKINVDCx14_ASAP7_75t_R g1013 ( 
.A(n_577),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_537),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_537),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_622),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_622),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_622),
.Y(n_1018)
);

INVxp67_ASAP7_75t_SL g1019 ( 
.A(n_902),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_622),
.Y(n_1020)
);

INVxp67_ASAP7_75t_SL g1021 ( 
.A(n_902),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_852),
.Y(n_1022)
);

INVxp67_ASAP7_75t_SL g1023 ( 
.A(n_800),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_773),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_777),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_800),
.Y(n_1026)
);

INVxp67_ASAP7_75t_SL g1027 ( 
.A(n_800),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_882),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_622),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_919),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_787),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_765),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_539),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_777),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_531),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_626),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_529),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_626),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_626),
.Y(n_1039)
);

INVxp33_ASAP7_75t_SL g1040 ( 
.A(n_535),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_538),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_626),
.Y(n_1042)
);

CKINVDCx14_ASAP7_75t_R g1043 ( 
.A(n_585),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_626),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_868),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_540),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_868),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_543),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_765),
.Y(n_1049)
);

CKINVDCx14_ASAP7_75t_R g1050 ( 
.A(n_542),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_532),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_642),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_642),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_642),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_642),
.Y(n_1055)
);

CKINVDCx14_ASAP7_75t_R g1056 ( 
.A(n_542),
.Y(n_1056)
);

INVxp33_ASAP7_75t_SL g1057 ( 
.A(n_544),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_868),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_546),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_642),
.Y(n_1060)
);

CKINVDCx16_ASAP7_75t_R g1061 ( 
.A(n_542),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_548),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_654),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_534),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_654),
.Y(n_1065)
);

CKINVDCx16_ASAP7_75t_R g1066 ( 
.A(n_542),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_549),
.Y(n_1067)
);

NOR2xp67_ASAP7_75t_L g1068 ( 
.A(n_595),
.B(n_0),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_654),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_654),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_654),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_660),
.Y(n_1072)
);

INVxp67_ASAP7_75t_SL g1073 ( 
.A(n_595),
.Y(n_1073)
);

INVxp33_ASAP7_75t_SL g1074 ( 
.A(n_550),
.Y(n_1074)
);

INVxp33_ASAP7_75t_SL g1075 ( 
.A(n_554),
.Y(n_1075)
);

INVxp67_ASAP7_75t_SL g1076 ( 
.A(n_595),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_660),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_556),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_660),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_660),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_545),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_558),
.Y(n_1082)
);

CKINVDCx16_ASAP7_75t_R g1083 ( 
.A(n_646),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_545),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_551),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_551),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_765),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_557),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_557),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_581),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_613),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_660),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_581),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_582),
.Y(n_1094)
);

INVxp67_ASAP7_75t_SL g1095 ( 
.A(n_801),
.Y(n_1095)
);

INVx4_ASAP7_75t_R g1096 ( 
.A(n_832),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_582),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_552),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_627),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_627),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_662),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_662),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_688),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_688),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_561),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_563),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_801),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_801),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_567),
.Y(n_1109)
);

INVxp67_ASAP7_75t_SL g1110 ( 
.A(n_801),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_700),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_569),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_700),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_772),
.Y(n_1114)
);

INVxp67_ASAP7_75t_SL g1115 ( 
.A(n_801),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_772),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_573),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_536),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_574),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_799),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_799),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_827),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_827),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_765),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_829),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_829),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_867),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_867),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_578),
.Y(n_1129)
);

CKINVDCx16_ASAP7_75t_R g1130 ( 
.A(n_646),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_875),
.Y(n_1131)
);

CKINVDCx16_ASAP7_75t_R g1132 ( 
.A(n_646),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_875),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_886),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_886),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_893),
.Y(n_1136)
);

INVxp33_ASAP7_75t_SL g1137 ( 
.A(n_584),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_559),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_893),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_916),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_916),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_588),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_589),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_926),
.Y(n_1144)
);

INVxp67_ASAP7_75t_L g1145 ( 
.A(n_529),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_926),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_591),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_838),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_838),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_559),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_579),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_579),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_625),
.Y(n_1153)
);

INVxp67_ASAP7_75t_SL g1154 ( 
.A(n_838),
.Y(n_1154)
);

INVxp67_ASAP7_75t_SL g1155 ( 
.A(n_838),
.Y(n_1155)
);

CKINVDCx16_ASAP7_75t_R g1156 ( 
.A(n_646),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_625),
.Y(n_1157)
);

INVxp33_ASAP7_75t_SL g1158 ( 
.A(n_593),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_596),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_838),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_597),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_816),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_541),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_816),
.Y(n_1164)
);

INVxp33_ASAP7_75t_SL g1165 ( 
.A(n_599),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_934),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_934),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_580),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_844),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_844),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_851),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_844),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_600),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_844),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_601),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_844),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_653),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_761),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_533),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_604),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_533),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_547),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_547),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_555),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_605),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_609),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_555),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_560),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_560),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_564),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_564),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_565),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_611),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_565),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_617),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_655),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_651),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_572),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_562),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_572),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_586),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_586),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_761),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_590),
.Y(n_1204)
);

CKINVDCx14_ASAP7_75t_R g1205 ( 
.A(n_851),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_590),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_761),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_592),
.B(n_0),
.Y(n_1208)
);

INVxp67_ASAP7_75t_SL g1209 ( 
.A(n_896),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_615),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_761),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_592),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_602),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_602),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_612),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_612),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_761),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_619),
.Y(n_1218)
);

CKINVDCx16_ASAP7_75t_R g1219 ( 
.A(n_851),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_620),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_761),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_620),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_628),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_624),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_896),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_761),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_624),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_629),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_630),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_632),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_632),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_636),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_761),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_639),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_761),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_637),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_583),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_583),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_598),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_598),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_607),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_607),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_608),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_608),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_730),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_678),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_730),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_640),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_786),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_786),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_566),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_805),
.Y(n_1252)
);

INVxp67_ASAP7_75t_SL g1253 ( 
.A(n_568),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_639),
.B(n_1),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_570),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_805),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_810),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_810),
.Y(n_1258)
);

BUFx5_ASAP7_75t_L g1259 ( 
.A(n_641),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_571),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_641),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_645),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_815),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_815),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_872),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_575),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_576),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_872),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_645),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_883),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_692),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_648),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_648),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_883),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_647),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_656),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_656),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_658),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_657),
.Y(n_1279)
);

CKINVDCx16_ASAP7_75t_R g1280 ( 
.A(n_851),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_661),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_657),
.Y(n_1282)
);

INVxp67_ASAP7_75t_SL g1283 ( 
.A(n_811),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_663),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_663),
.Y(n_1285)
);

INVxp67_ASAP7_75t_SL g1286 ( 
.A(n_862),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_667),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_667),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_672),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_672),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_664),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_690),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_690),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_699),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_666),
.Y(n_1295)
);

NOR2xp67_ASAP7_75t_L g1296 ( 
.A(n_618),
.B(n_2),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_699),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_669),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_671),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_702),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_673),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_674),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_702),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_675),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_705),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_705),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_613),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_706),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_587),
.Y(n_1309)
);

INVxp67_ASAP7_75t_SL g1310 ( 
.A(n_832),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_613),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_706),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_709),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_676),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_709),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_712),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_712),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_677),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_723),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_679),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_683),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1067),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1095),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1310),
.B(n_603),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1110),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_959),
.Y(n_1326)
);

CKINVDCx16_ASAP7_75t_R g1327 ( 
.A(n_1050),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1115),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1154),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1073),
.B(n_1076),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1155),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_996),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1051),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1064),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1169),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1118),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1163),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1170),
.Y(n_1338)
);

CKINVDCx16_ASAP7_75t_R g1339 ( 
.A(n_1056),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1172),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_996),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1003),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_1009),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1199),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1003),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_963),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1251),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1255),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1174),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_964),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1176),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1010),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1019),
.B(n_616),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1021),
.B(n_623),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1010),
.Y(n_1355)
);

INVxp67_ASAP7_75t_SL g1356 ( 
.A(n_1009),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1011),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_1035),
.B(n_631),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1011),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1260),
.Y(n_1360)
);

INVxp33_ASAP7_75t_L g1361 ( 
.A(n_1228),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1196),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_978),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1012),
.Y(n_1364)
);

INVxp67_ASAP7_75t_SL g1365 ( 
.A(n_1023),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_982),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1266),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1267),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1012),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1014),
.Y(n_1370)
);

INVxp67_ASAP7_75t_SL g1371 ( 
.A(n_1027),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1014),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1309),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1040),
.B(n_633),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1033),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_984),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1015),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1031),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1080),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1013),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1043),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1015),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1016),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_SL g1384 ( 
.A(n_1032),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1016),
.Y(n_1385)
);

CKINVDCx16_ASAP7_75t_R g1386 ( 
.A(n_1205),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_968),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1017),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1017),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1018),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1061),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1018),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1066),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1020),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1040),
.B(n_634),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_968),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1020),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1029),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1080),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1029),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1036),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_990),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_990),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1036),
.Y(n_1404)
);

CKINVDCx16_ASAP7_75t_R g1405 ( 
.A(n_1083),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1130),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1038),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1132),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1038),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1039),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1039),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1156),
.Y(n_1412)
);

INVxp67_ASAP7_75t_SL g1413 ( 
.A(n_1209),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1035),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1057),
.B(n_635),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1042),
.Y(n_1416)
);

INVxp67_ASAP7_75t_SL g1417 ( 
.A(n_1307),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1042),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1044),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1022),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1041),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1044),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1041),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1098),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1052),
.Y(n_1425)
);

CKINVDCx16_ASAP7_75t_R g1426 ( 
.A(n_1219),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1052),
.Y(n_1427)
);

CKINVDCx20_ASAP7_75t_R g1428 ( 
.A(n_1280),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1046),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1053),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1053),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1054),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1054),
.Y(n_1433)
);

INVxp67_ASAP7_75t_SL g1434 ( 
.A(n_1307),
.Y(n_1434)
);

INVxp33_ASAP7_75t_SL g1435 ( 
.A(n_1022),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1232),
.B(n_859),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1055),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1057),
.B(n_643),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1046),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1048),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1307),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1055),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1048),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1060),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1028),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1059),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1028),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1059),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1060),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1062),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1063),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1063),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1030),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1030),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1065),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1168),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1195),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1062),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1078),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1065),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1069),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1069),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1078),
.Y(n_1463)
);

CKINVDCx20_ASAP7_75t_R g1464 ( 
.A(n_1197),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1082),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1196),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_1246),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1070),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1082),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1070),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1271),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1105),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_973),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1071),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1105),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1106),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_R g1477 ( 
.A(n_1106),
.B(n_644),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1092),
.Y(n_1478)
);

NAND2xp33_ASAP7_75t_R g1479 ( 
.A(n_1109),
.B(n_684),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1109),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_1112),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1071),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1112),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1072),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1117),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1117),
.Y(n_1486)
);

CKINVDCx20_ASAP7_75t_R g1487 ( 
.A(n_1119),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1119),
.Y(n_1488)
);

INVxp33_ASAP7_75t_L g1489 ( 
.A(n_1320),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1129),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1072),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1129),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1142),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_1142),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1092),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_1143),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1077),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1143),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1077),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1147),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1079),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1074),
.B(n_650),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1079),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1026),
.Y(n_1504)
);

NOR2xp67_ASAP7_75t_L g1505 ( 
.A(n_1147),
.B(n_659),
.Y(n_1505)
);

INVxp67_ASAP7_75t_SL g1506 ( 
.A(n_1321),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1159),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1159),
.Y(n_1508)
);

NOR2xp67_ASAP7_75t_L g1509 ( 
.A(n_1161),
.B(n_681),
.Y(n_1509)
);

INVxp33_ASAP7_75t_SL g1510 ( 
.A(n_1161),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1026),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1045),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1175),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1045),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1047),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1047),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1074),
.B(n_682),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1058),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_1175),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1058),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1107),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1180),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1180),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1107),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1075),
.B(n_711),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1108),
.Y(n_1526)
);

INVxp33_ASAP7_75t_L g1527 ( 
.A(n_967),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1108),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_973),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1150),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1032),
.B(n_859),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1186),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1148),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1186),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_SL g1535 ( 
.A(n_1049),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1148),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1149),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1149),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1193),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1160),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1160),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1081),
.Y(n_1542)
);

INVxp33_ASAP7_75t_L g1543 ( 
.A(n_970),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1259),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1259),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1084),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1259),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1193),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1210),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1085),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1210),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1218),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1218),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1223),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1086),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1088),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1223),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1229),
.Y(n_1558)
);

CKINVDCx20_ASAP7_75t_R g1559 ( 
.A(n_1229),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1049),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1089),
.Y(n_1561)
);

CKINVDCx20_ASAP7_75t_R g1562 ( 
.A(n_1236),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1236),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1248),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1090),
.Y(n_1565)
);

CKINVDCx16_ASAP7_75t_R g1566 ( 
.A(n_1087),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1093),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1094),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1097),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1099),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1100),
.Y(n_1571)
);

INVxp67_ASAP7_75t_SL g1572 ( 
.A(n_1087),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1173),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1151),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_1124),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1101),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_1248),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1275),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1275),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1278),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1102),
.Y(n_1581)
);

NOR2xp67_ASAP7_75t_L g1582 ( 
.A(n_1278),
.B(n_714),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1152),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_1281),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1281),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1103),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1291),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1291),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1295),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1104),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1111),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1295),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1124),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1113),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1259),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1298),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1075),
.B(n_726),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_973),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1114),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1298),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1299),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1116),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1299),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1120),
.Y(n_1604)
);

INVxp33_ASAP7_75t_SL g1605 ( 
.A(n_1302),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1302),
.Y(n_1606)
);

BUFx2_ASAP7_75t_SL g1607 ( 
.A(n_1171),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_1304),
.Y(n_1608)
);

INVxp33_ASAP7_75t_SL g1609 ( 
.A(n_1304),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1121),
.Y(n_1610)
);

NOR2xp67_ASAP7_75t_L g1611 ( 
.A(n_1314),
.B(n_727),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1137),
.B(n_741),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1253),
.B(n_948),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1122),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1123),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1125),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1126),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1259),
.Y(n_1618)
);

INVxp67_ASAP7_75t_SL g1619 ( 
.A(n_973),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1314),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1318),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1127),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1318),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1137),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1128),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1131),
.Y(n_1626)
);

CKINVDCx20_ASAP7_75t_R g1627 ( 
.A(n_1173),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1133),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1134),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_1185),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1135),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1136),
.Y(n_1632)
);

INVxp67_ASAP7_75t_SL g1633 ( 
.A(n_973),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1185),
.B(n_859),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1158),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1473),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1332),
.B(n_1244),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1379),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1379),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1542),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1473),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1332),
.B(n_1244),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1417),
.B(n_1225),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1546),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1434),
.B(n_1225),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1550),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_1456),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1555),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1330),
.A2(n_956),
.B(n_955),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1362),
.B(n_1250),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1424),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1473),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1441),
.B(n_957),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1556),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1413),
.B(n_960),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1362),
.B(n_1250),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1561),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1565),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1473),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1456),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1466),
.Y(n_1661)
);

AND2x2_ASAP7_75t_SL g1662 ( 
.A(n_1459),
.B(n_1208),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1560),
.B(n_1158),
.Y(n_1663)
);

INVx4_ASAP7_75t_L g1664 ( 
.A(n_1529),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1567),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1568),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1333),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1569),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1457),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1365),
.B(n_961),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_1457),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1399),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1570),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1466),
.B(n_1256),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1529),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1529),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1464),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1571),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1529),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1371),
.B(n_1256),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1566),
.B(n_1068),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1598),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1464),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1399),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1341),
.B(n_1343),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1467),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1467),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1576),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1581),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1586),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1598),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1478),
.Y(n_1692)
);

NAND2xp33_ASAP7_75t_L g1693 ( 
.A(n_1613),
.B(n_613),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1590),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1598),
.Y(n_1695)
);

BUFx6f_ASAP7_75t_L g1696 ( 
.A(n_1530),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1591),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1594),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_1471),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1599),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1323),
.B(n_965),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1530),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1575),
.B(n_1165),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1602),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1478),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1604),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1495),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1495),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1334),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1479),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1521),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1356),
.B(n_1265),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1471),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1524),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1325),
.B(n_969),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1574),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1610),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1614),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1607),
.B(n_1265),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1328),
.B(n_1329),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1506),
.A2(n_1573),
.B1(n_1322),
.B2(n_1354),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1504),
.B(n_1274),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1615),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1331),
.B(n_971),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1616),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1526),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1324),
.B(n_972),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1353),
.B(n_1165),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1617),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1544),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1622),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1574),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1528),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1336),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1533),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1625),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1536),
.Y(n_1737)
);

CKINVDCx16_ASAP7_75t_R g1738 ( 
.A(n_1327),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1626),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1583),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1339),
.B(n_1386),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1634),
.A2(n_1593),
.B1(n_1572),
.B2(n_966),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1619),
.B(n_975),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1583),
.B(n_1274),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1628),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1511),
.B(n_1139),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1512),
.B(n_1140),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1629),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1337),
.Y(n_1749)
);

AND2x2_ASAP7_75t_SL g1750 ( 
.A(n_1558),
.B(n_1208),
.Y(n_1750)
);

BUFx2_ASAP7_75t_L g1751 ( 
.A(n_1627),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1537),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1631),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1632),
.B(n_1312),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1352),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1355),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1357),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1359),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1538),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1540),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1544),
.Y(n_1761)
);

NOR2x1_ASAP7_75t_L g1762 ( 
.A(n_1358),
.B(n_1296),
.Y(n_1762)
);

INVx6_ASAP7_75t_L g1763 ( 
.A(n_1531),
.Y(n_1763)
);

AOI22x1_ASAP7_75t_SL g1764 ( 
.A1(n_1373),
.A2(n_721),
.B1(n_722),
.B2(n_707),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1514),
.B(n_1515),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1541),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1364),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1369),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_1370),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1505),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1372),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1516),
.B(n_1317),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1377),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1436),
.A2(n_966),
.B1(n_1286),
.B2(n_1283),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1382),
.Y(n_1775)
);

OAI21x1_ASAP7_75t_L g1776 ( 
.A1(n_1545),
.A2(n_979),
.B(n_977),
.Y(n_1776)
);

CKINVDCx20_ASAP7_75t_R g1777 ( 
.A(n_1326),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1383),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1374),
.B(n_1301),
.Y(n_1779)
);

CKINVDCx20_ASAP7_75t_R g1780 ( 
.A(n_1326),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1385),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1388),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1389),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1518),
.B(n_1141),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1390),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1395),
.A2(n_1301),
.B1(n_1006),
.B2(n_1025),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_1342),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1545),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1392),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1520),
.B(n_1308),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1335),
.B(n_1144),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1394),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1397),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1398),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1400),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1401),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_R g1797 ( 
.A(n_1396),
.B(n_763),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1633),
.B(n_980),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1404),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1509),
.B(n_983),
.Y(n_1800)
);

CKINVDCx20_ASAP7_75t_R g1801 ( 
.A(n_1346),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1547),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1407),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1409),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1410),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1415),
.A2(n_952),
.B1(n_1008),
.B2(n_962),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1582),
.B(n_985),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1411),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1345),
.Y(n_1809)
);

OA21x2_ASAP7_75t_L g1810 ( 
.A1(n_1416),
.A2(n_988),
.B(n_987),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1338),
.B(n_1146),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1418),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1419),
.Y(n_1813)
);

CKINVDCx8_ASAP7_75t_R g1814 ( 
.A(n_1405),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1422),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1425),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1427),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1430),
.Y(n_1818)
);

BUFx3_ASAP7_75t_L g1819 ( 
.A(n_1431),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_L g1820 ( 
.A(n_1438),
.B(n_1171),
.C(n_1024),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1432),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1611),
.B(n_953),
.Y(n_1822)
);

AOI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1502),
.A2(n_1525),
.B1(n_1597),
.B2(n_1517),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1612),
.B(n_953),
.Y(n_1824)
);

CKINVDCx20_ASAP7_75t_R g1825 ( 
.A(n_1346),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1433),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1620),
.A2(n_1034),
.B1(n_1254),
.B2(n_1024),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1510),
.A2(n_995),
.B1(n_606),
.B2(n_621),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1437),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1442),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1340),
.B(n_1308),
.Y(n_1831)
);

CKINVDCx16_ASAP7_75t_R g1832 ( 
.A(n_1426),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1547),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1444),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1595),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1449),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1451),
.Y(n_1837)
);

CKINVDCx20_ASAP7_75t_R g1838 ( 
.A(n_1350),
.Y(n_1838)
);

INVx3_ASAP7_75t_L g1839 ( 
.A(n_1595),
.Y(n_1839)
);

BUFx6f_ASAP7_75t_L g1840 ( 
.A(n_1452),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_1627),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1455),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1460),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1461),
.Y(n_1844)
);

BUFx2_ASAP7_75t_L g1845 ( 
.A(n_1630),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1462),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1349),
.B(n_1153),
.Y(n_1847)
);

BUFx2_ASAP7_75t_L g1848 ( 
.A(n_1630),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_R g1849 ( 
.A(n_1402),
.B(n_776),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1468),
.B(n_991),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1351),
.B(n_1313),
.Y(n_1851)
);

INVx1_ASAP7_75t_SL g1852 ( 
.A(n_1472),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1344),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1470),
.B(n_1157),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1474),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1482),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1484),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1491),
.B(n_1162),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1497),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1499),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1501),
.Y(n_1861)
);

OA21x2_ASAP7_75t_L g1862 ( 
.A1(n_1503),
.A2(n_992),
.B(n_991),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1361),
.B(n_981),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1618),
.B(n_992),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1347),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1489),
.B(n_995),
.Y(n_1866)
);

BUFx8_ASAP7_75t_L g1867 ( 
.A(n_1384),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1510),
.A2(n_665),
.B1(n_668),
.B2(n_530),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1618),
.B(n_1312),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1523),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1477),
.B(n_993),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1384),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1553),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1563),
.B(n_1313),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1605),
.B(n_993),
.Y(n_1875)
);

BUFx6f_ASAP7_75t_L g1876 ( 
.A(n_1420),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1384),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_R g1878 ( 
.A(n_1403),
.B(n_791),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1605),
.B(n_994),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1527),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1414),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1609),
.A2(n_1254),
.B1(n_686),
.B2(n_687),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1421),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1535),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1543),
.B(n_1164),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1535),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1535),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1348),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1423),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1472),
.A2(n_736),
.B1(n_770),
.B2(n_724),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1429),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1439),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1440),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1609),
.B(n_1259),
.Y(n_1894)
);

AND2x4_ASAP7_75t_L g1895 ( 
.A(n_1380),
.B(n_1317),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1450),
.B(n_974),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1463),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1465),
.B(n_974),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1469),
.Y(n_1899)
);

INVx4_ASAP7_75t_L g1900 ( 
.A(n_1380),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1475),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1476),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1483),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1360),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1485),
.Y(n_1905)
);

BUFx2_ASAP7_75t_L g1906 ( 
.A(n_1445),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_1367),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1486),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1488),
.B(n_974),
.Y(n_1909)
);

AND2x2_ASAP7_75t_SL g1910 ( 
.A(n_1435),
.B(n_723),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1381),
.B(n_1166),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1490),
.Y(n_1912)
);

INVx3_ASAP7_75t_L g1913 ( 
.A(n_1492),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1493),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1508),
.Y(n_1915)
);

CKINVDCx6p67_ASAP7_75t_R g1916 ( 
.A(n_1391),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1513),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1534),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1539),
.B(n_994),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1551),
.Y(n_1920)
);

AND2x4_ASAP7_75t_L g1921 ( 
.A(n_1381),
.B(n_1289),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1554),
.Y(n_1922)
);

CKINVDCx20_ASAP7_75t_R g1923 ( 
.A(n_1350),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1375),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1600),
.B(n_997),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1601),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1603),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1606),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1443),
.B(n_1289),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1435),
.B(n_1138),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1624),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1443),
.B(n_1167),
.Y(n_1932)
);

CKINVDCx20_ASAP7_75t_R g1933 ( 
.A(n_1363),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1446),
.Y(n_1934)
);

BUFx6f_ASAP7_75t_L g1935 ( 
.A(n_1446),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1448),
.B(n_1290),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1448),
.B(n_997),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1458),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1458),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1368),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1557),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1557),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1564),
.B(n_998),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1635),
.A2(n_817),
.B1(n_796),
.B2(n_802),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1564),
.B(n_998),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1578),
.Y(n_1946)
);

BUFx3_ASAP7_75t_L g1947 ( 
.A(n_1635),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1578),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1579),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1579),
.Y(n_1950)
);

INVx3_ASAP7_75t_L g1951 ( 
.A(n_1580),
.Y(n_1951)
);

BUFx2_ASAP7_75t_L g1952 ( 
.A(n_1445),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1580),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1585),
.Y(n_1954)
);

OA21x2_ASAP7_75t_L g1955 ( 
.A1(n_1623),
.A2(n_1000),
.B(n_999),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1585),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1588),
.Y(n_1957)
);

INVx3_ASAP7_75t_L g1958 ( 
.A(n_1588),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1621),
.B(n_1290),
.Y(n_1959)
);

BUFx6f_ASAP7_75t_L g1960 ( 
.A(n_1621),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1623),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1480),
.Y(n_1962)
);

INVx3_ASAP7_75t_L g1963 ( 
.A(n_1387),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1480),
.B(n_1292),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1387),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1373),
.B(n_999),
.Y(n_1966)
);

NAND2x1p5_ASAP7_75t_L g1967 ( 
.A(n_1481),
.B(n_1000),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1481),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1487),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1487),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1375),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_SL g1972 ( 
.A1(n_1494),
.A2(n_798),
.B1(n_823),
.B2(n_780),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1494),
.Y(n_1973)
);

INVxp67_ASAP7_75t_L g1974 ( 
.A(n_1651),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1824),
.B(n_1259),
.Y(n_1975)
);

INVxp67_ASAP7_75t_L g1976 ( 
.A(n_1863),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1650),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1776),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1776),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1650),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1823),
.B(n_1259),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1869),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1727),
.B(n_1002),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1696),
.Y(n_1984)
);

BUFx6f_ASAP7_75t_L g1985 ( 
.A(n_1696),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1650),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1869),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1728),
.A2(n_1498),
.B1(n_1500),
.B2(n_1496),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1862),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_L g1990 ( 
.A(n_1875),
.B(n_685),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1862),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1869),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1656),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1862),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1656),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1638),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1656),
.Y(n_1997)
);

BUFx8_ASAP7_75t_L g1998 ( 
.A(n_1677),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1680),
.B(n_1138),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1674),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1638),
.Y(n_2001)
);

INVx3_ASAP7_75t_L g2002 ( 
.A(n_1810),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1639),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1639),
.Y(n_2004)
);

OAI22xp5_ASAP7_75t_SL g2005 ( 
.A1(n_1890),
.A2(n_1366),
.B1(n_1363),
.B2(n_924),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1672),
.Y(n_2006)
);

BUFx3_ASAP7_75t_L g2007 ( 
.A(n_1661),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1674),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1674),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1879),
.B(n_795),
.Y(n_2010)
);

INVx1_ASAP7_75t_SL g2011 ( 
.A(n_1686),
.Y(n_2011)
);

XNOR2xp5_ASAP7_75t_L g2012 ( 
.A(n_1972),
.B(n_1366),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1672),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1684),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1637),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1637),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1684),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1692),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1637),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1642),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1692),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1642),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1642),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1744),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1696),
.Y(n_2025)
);

OAI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_1806),
.A2(n_652),
.B1(n_864),
.B2(n_618),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1744),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1719),
.B(n_1002),
.Y(n_2028)
);

OAI22xp5_ASAP7_75t_SL g2029 ( 
.A1(n_1647),
.A2(n_1671),
.B1(n_1687),
.B2(n_1660),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1929),
.B(n_820),
.Y(n_2030)
);

INVx6_ASAP7_75t_L g2031 ( 
.A(n_1867),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1719),
.B(n_1007),
.Y(n_2032)
);

AOI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1779),
.A2(n_1498),
.B1(n_1500),
.B2(n_1496),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1744),
.Y(n_2034)
);

BUFx6f_ASAP7_75t_L g2035 ( 
.A(n_1696),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_1702),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1655),
.B(n_1007),
.Y(n_2037)
);

AOI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_1710),
.A2(n_1685),
.B1(n_1943),
.B2(n_1937),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1945),
.B(n_691),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1705),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1765),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1680),
.B(n_1037),
.Y(n_2042)
);

AOI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1685),
.A2(n_1519),
.B1(n_1522),
.B2(n_1507),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1765),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1640),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1874),
.B(n_1145),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1644),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1646),
.Y(n_2048)
);

INVx1_ASAP7_75t_SL g2049 ( 
.A(n_1880),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1929),
.B(n_824),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1648),
.Y(n_2051)
);

BUFx2_ASAP7_75t_L g2052 ( 
.A(n_1677),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_1964),
.Y(n_2053)
);

AOI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_1685),
.A2(n_1519),
.B1(n_1522),
.B2(n_1507),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1705),
.Y(n_2055)
);

INVxp67_ASAP7_75t_L g2056 ( 
.A(n_1866),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1654),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1707),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1707),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1657),
.Y(n_2060)
);

OAI21x1_ASAP7_75t_L g2061 ( 
.A1(n_1649),
.A2(n_1203),
.B(n_1178),
.Y(n_2061)
);

NAND2xp33_ASAP7_75t_SL g2062 ( 
.A(n_1919),
.B(n_830),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1658),
.Y(n_2063)
);

CKINVDCx11_ASAP7_75t_R g2064 ( 
.A(n_1814),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1665),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1708),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1670),
.B(n_826),
.Y(n_2067)
);

BUFx6f_ASAP7_75t_L g2068 ( 
.A(n_1702),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1666),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1874),
.B(n_1261),
.Y(n_2070)
);

AND2x6_ASAP7_75t_L g2071 ( 
.A(n_1872),
.B(n_728),
.Y(n_2071)
);

INVx1_ASAP7_75t_SL g2072 ( 
.A(n_1647),
.Y(n_2072)
);

BUFx8_ASAP7_75t_L g2073 ( 
.A(n_1683),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1668),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1673),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1678),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1688),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1874),
.B(n_1269),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1689),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_1925),
.B(n_694),
.Y(n_2080)
);

BUFx6f_ASAP7_75t_L g2081 ( 
.A(n_1702),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1690),
.Y(n_2082)
);

OAI22xp5_ASAP7_75t_SL g2083 ( 
.A1(n_1660),
.A2(n_932),
.B1(n_945),
.B2(n_929),
.Y(n_2083)
);

BUFx4f_ASAP7_75t_L g2084 ( 
.A(n_1955),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1694),
.Y(n_2085)
);

INVx4_ASAP7_75t_L g2086 ( 
.A(n_1691),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1810),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1708),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1810),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1711),
.Y(n_2090)
);

INVxp67_ASAP7_75t_L g2091 ( 
.A(n_1930),
.Y(n_2091)
);

INVx3_ASAP7_75t_L g2092 ( 
.A(n_1682),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1929),
.B(n_1292),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1711),
.Y(n_2094)
);

INVxp67_ASAP7_75t_L g2095 ( 
.A(n_1663),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1697),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_1966),
.B(n_698),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1936),
.B(n_843),
.Y(n_2098)
);

HB1xp67_ASAP7_75t_L g2099 ( 
.A(n_1964),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_1894),
.A2(n_1548),
.B1(n_1549),
.B2(n_1532),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1871),
.B(n_854),
.Y(n_2101)
);

AND2x6_ASAP7_75t_L g2102 ( 
.A(n_1872),
.B(n_728),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1714),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_1661),
.B(n_1179),
.Y(n_2104)
);

NAND2x1_ASAP7_75t_L g2105 ( 
.A(n_1682),
.B(n_1096),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1714),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1698),
.Y(n_2107)
);

INVxp67_ASAP7_75t_L g2108 ( 
.A(n_1885),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1700),
.Y(n_2109)
);

AND3x1_ASAP7_75t_L g2110 ( 
.A(n_1828),
.B(n_937),
.C(n_732),
.Y(n_2110)
);

INVx1_ASAP7_75t_SL g2111 ( 
.A(n_1671),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_1712),
.B(n_1704),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1726),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_1936),
.B(n_1959),
.Y(n_2114)
);

BUFx6f_ASAP7_75t_SL g2115 ( 
.A(n_1900),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1726),
.Y(n_2116)
);

OAI22xp33_ASAP7_75t_SL g2117 ( 
.A1(n_1763),
.A2(n_731),
.B1(n_734),
.B2(n_732),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1936),
.B(n_856),
.Y(n_2118)
);

BUFx2_ASAP7_75t_L g2119 ( 
.A(n_1683),
.Y(n_2119)
);

AOI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_1894),
.A2(n_1548),
.B1(n_1549),
.B2(n_1532),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1706),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1822),
.B(n_860),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_1712),
.B(n_1181),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1717),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1733),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1643),
.B(n_894),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1645),
.B(n_912),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1718),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1723),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1733),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1959),
.B(n_921),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1712),
.B(n_944),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1735),
.Y(n_2133)
);

AND2x4_ASAP7_75t_L g2134 ( 
.A(n_1725),
.B(n_1182),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1729),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1800),
.B(n_949),
.Y(n_2136)
);

AOI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_1742),
.A2(n_1559),
.B1(n_1562),
.B2(n_1552),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1731),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1736),
.Y(n_2139)
);

NAND2xp33_ASAP7_75t_R g2140 ( 
.A(n_1955),
.B(n_1376),
.Y(n_2140)
);

OAI22xp5_ASAP7_75t_SL g2141 ( 
.A1(n_1687),
.A2(n_1699),
.B1(n_1559),
.B2(n_1562),
.Y(n_2141)
);

NAND2xp33_ASAP7_75t_SL g2142 ( 
.A(n_1959),
.B(n_652),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1739),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1745),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_1662),
.B(n_954),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1735),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_SL g2147 ( 
.A1(n_1699),
.A2(n_1577),
.B1(n_1584),
.B2(n_1552),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1748),
.Y(n_2148)
);

INVx3_ASAP7_75t_L g2149 ( 
.A(n_1682),
.Y(n_2149)
);

AOI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_1763),
.A2(n_1584),
.B1(n_1587),
.B2(n_1577),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1753),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1807),
.B(n_954),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1746),
.Y(n_2153)
);

OAI22xp5_ASAP7_75t_SL g2154 ( 
.A1(n_1910),
.A2(n_1589),
.B1(n_1592),
.B2(n_1587),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1737),
.Y(n_2155)
);

INVxp67_ASAP7_75t_L g2156 ( 
.A(n_1885),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1746),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1747),
.Y(n_2158)
);

NAND2xp33_ASAP7_75t_L g2159 ( 
.A(n_1864),
.B(n_1091),
.Y(n_2159)
);

BUFx6f_ASAP7_75t_L g2160 ( 
.A(n_1702),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1737),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1747),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1784),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1784),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_1662),
.B(n_958),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1750),
.B(n_958),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1754),
.Y(n_2167)
);

BUFx6f_ASAP7_75t_L g2168 ( 
.A(n_1716),
.Y(n_2168)
);

HB1xp67_ASAP7_75t_L g2169 ( 
.A(n_1964),
.Y(n_2169)
);

HB1xp67_ASAP7_75t_L g2170 ( 
.A(n_1713),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1752),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_1750),
.B(n_976),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1754),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_1716),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1754),
.Y(n_2175)
);

HB1xp67_ASAP7_75t_L g2176 ( 
.A(n_1713),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1847),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1847),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1752),
.Y(n_2179)
);

INVx3_ASAP7_75t_L g2180 ( 
.A(n_1730),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_1669),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1701),
.B(n_976),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1921),
.B(n_986),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1854),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1854),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1858),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_1858),
.B(n_1293),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1715),
.B(n_986),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1722),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_1955),
.B(n_1293),
.Y(n_2190)
);

AND2x4_ASAP7_75t_L g2191 ( 
.A(n_1716),
.B(n_1732),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1921),
.B(n_989),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1722),
.Y(n_2193)
);

BUFx6f_ASAP7_75t_L g2194 ( 
.A(n_1716),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_1732),
.B(n_1183),
.Y(n_2195)
);

AOI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_1763),
.A2(n_1592),
.B1(n_1596),
.B2(n_1589),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1791),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1791),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_1730),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1811),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_1763),
.B(n_1294),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_1667),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_1811),
.B(n_1294),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1831),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1831),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1831),
.Y(n_2206)
);

BUFx3_ASAP7_75t_L g2207 ( 
.A(n_1732),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1759),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1759),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_1820),
.B(n_701),
.Y(n_2210)
);

INVx3_ASAP7_75t_L g2211 ( 
.A(n_1730),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1760),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1851),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1851),
.Y(n_2214)
);

BUFx2_ASAP7_75t_L g2215 ( 
.A(n_1876),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_SL g2216 ( 
.A(n_1921),
.B(n_989),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1851),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1799),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1760),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1799),
.Y(n_2220)
);

INVxp67_ASAP7_75t_L g2221 ( 
.A(n_1932),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_1895),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1766),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1818),
.Y(n_2224)
);

OAI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_1774),
.A2(n_703),
.B1(n_708),
.B2(n_704),
.Y(n_2225)
);

BUFx2_ASAP7_75t_L g2226 ( 
.A(n_1876),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1910),
.B(n_1932),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1766),
.Y(n_2228)
);

INVx3_ASAP7_75t_L g2229 ( 
.A(n_1761),
.Y(n_2229)
);

NAND2x1_ASAP7_75t_L g2230 ( 
.A(n_1664),
.B(n_1091),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_1895),
.B(n_1297),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1818),
.Y(n_2232)
);

INVx3_ASAP7_75t_L g2233 ( 
.A(n_1761),
.Y(n_2233)
);

BUFx6f_ASAP7_75t_L g2234 ( 
.A(n_1732),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1724),
.B(n_1001),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1819),
.Y(n_2236)
);

BUFx6f_ASAP7_75t_L g2237 ( 
.A(n_1740),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_1895),
.Y(n_2238)
);

NOR2x1_ASAP7_75t_L g2239 ( 
.A(n_1931),
.B(n_1596),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1772),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1772),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_1967),
.B(n_1297),
.Y(n_2242)
);

NOR2xp33_ASAP7_75t_L g2243 ( 
.A(n_1721),
.B(n_710),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_1761),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_1740),
.B(n_1184),
.Y(n_2245)
);

HB1xp67_ASAP7_75t_L g2246 ( 
.A(n_1876),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1819),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1772),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1755),
.Y(n_2249)
);

INVxp67_ASAP7_75t_L g2250 ( 
.A(n_1896),
.Y(n_2250)
);

OAI22xp5_ASAP7_75t_SL g2251 ( 
.A1(n_1777),
.A2(n_1608),
.B1(n_1453),
.B2(n_1454),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1756),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1757),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1758),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1767),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1790),
.Y(n_2256)
);

NOR2x1_ASAP7_75t_L g2257 ( 
.A(n_1900),
.B(n_1608),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1771),
.Y(n_2258)
);

INVx3_ASAP7_75t_L g2259 ( 
.A(n_1788),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1790),
.Y(n_2260)
);

OAI22xp5_ASAP7_75t_SL g2261 ( 
.A1(n_1777),
.A2(n_1453),
.B1(n_1454),
.B2(n_1447),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1778),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1790),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1781),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1782),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1792),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1794),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_1788),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1796),
.Y(n_2269)
);

NAND2xp33_ASAP7_75t_SL g2270 ( 
.A(n_1770),
.B(n_864),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_1967),
.B(n_1300),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1803),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_1740),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_1653),
.B(n_1001),
.Y(n_2274)
);

BUFx6f_ASAP7_75t_L g2275 ( 
.A(n_1740),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1788),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1802),
.B(n_1004),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1804),
.Y(n_2278)
);

BUFx6f_ASAP7_75t_L g2279 ( 
.A(n_1636),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_SL g2280 ( 
.A(n_1769),
.B(n_1004),
.Y(n_2280)
);

INVx3_ASAP7_75t_L g2281 ( 
.A(n_1802),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_1802),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1833),
.B(n_1005),
.Y(n_2283)
);

OAI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_1786),
.A2(n_713),
.B1(n_717),
.B2(n_716),
.Y(n_2284)
);

INVx3_ASAP7_75t_L g2285 ( 
.A(n_1833),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_1833),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1805),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1812),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1815),
.Y(n_2289)
);

AOI22xp5_ASAP7_75t_L g2290 ( 
.A1(n_1681),
.A2(n_1447),
.B1(n_1393),
.B2(n_1406),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_1835),
.Y(n_2291)
);

OAI22xp5_ASAP7_75t_SL g2292 ( 
.A1(n_1780),
.A2(n_1378),
.B1(n_1376),
.B2(n_1391),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1817),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1835),
.B(n_1005),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1826),
.Y(n_2295)
);

INVx3_ASAP7_75t_L g2296 ( 
.A(n_1835),
.Y(n_2296)
);

CKINVDCx20_ASAP7_75t_R g2297 ( 
.A(n_1780),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1834),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_1967),
.B(n_1300),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_1769),
.B(n_1178),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1836),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_1787),
.B(n_1303),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1843),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1844),
.Y(n_2304)
);

NOR2x1_ASAP7_75t_L g2305 ( 
.A(n_1900),
.B(n_731),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_1787),
.B(n_1303),
.Y(n_2306)
);

AND2x4_ASAP7_75t_L g2307 ( 
.A(n_1855),
.B(n_1856),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1839),
.Y(n_2308)
);

CKINVDCx8_ASAP7_75t_R g2309 ( 
.A(n_1738),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1839),
.B(n_1091),
.Y(n_2310)
);

INVxp33_ASAP7_75t_L g2311 ( 
.A(n_1827),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1859),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_1839),
.B(n_1091),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_1636),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1860),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1768),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1768),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1773),
.Y(n_2318)
);

INVx4_ASAP7_75t_SL g2319 ( 
.A(n_2071),
.Y(n_2319)
);

AOI22xp5_ASAP7_75t_L g2320 ( 
.A1(n_2038),
.A2(n_1939),
.B1(n_1941),
.B2(n_1934),
.Y(n_2320)
);

INVx5_ASAP7_75t_L g2321 ( 
.A(n_1989),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2240),
.Y(n_2322)
);

CKINVDCx8_ASAP7_75t_R g2323 ( 
.A(n_2202),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2039),
.B(n_1762),
.Y(n_2324)
);

INVx3_ASAP7_75t_L g2325 ( 
.A(n_2092),
.Y(n_2325)
);

NOR2xp33_ASAP7_75t_L g2326 ( 
.A(n_2095),
.B(n_2091),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2039),
.B(n_1720),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_1978),
.Y(n_2328)
);

INVx4_ASAP7_75t_L g2329 ( 
.A(n_1984),
.Y(n_2329)
);

NAND2x1p5_ASAP7_75t_L g2330 ( 
.A(n_2226),
.B(n_1938),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2240),
.Y(n_2331)
);

CKINVDCx5p33_ASAP7_75t_R g2332 ( 
.A(n_2202),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2241),
.Y(n_2333)
);

INVx5_ASAP7_75t_L g2334 ( 
.A(n_1989),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_1978),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2084),
.B(n_2114),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_2279),
.Y(n_2337)
);

BUFx6f_ASAP7_75t_L g2338 ( 
.A(n_2279),
.Y(n_2338)
);

AND2x4_ASAP7_75t_L g2339 ( 
.A(n_2007),
.B(n_1877),
.Y(n_2339)
);

BUFx4f_ASAP7_75t_L g2340 ( 
.A(n_2031),
.Y(n_2340)
);

BUFx2_ASAP7_75t_L g2341 ( 
.A(n_2052),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_2279),
.Y(n_2342)
);

INVx1_ASAP7_75t_SL g2343 ( 
.A(n_2049),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_1979),
.Y(n_2344)
);

BUFx3_ASAP7_75t_L g2345 ( 
.A(n_2226),
.Y(n_2345)
);

AND2x4_ASAP7_75t_SL g2346 ( 
.A(n_2114),
.B(n_1876),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2241),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_2064),
.Y(n_2348)
);

BUFx4f_ASAP7_75t_L g2349 ( 
.A(n_2031),
.Y(n_2349)
);

BUFx6f_ASAP7_75t_L g2350 ( 
.A(n_2279),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_1979),
.Y(n_2351)
);

CKINVDCx5p33_ASAP7_75t_R g2352 ( 
.A(n_2064),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1996),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_L g2354 ( 
.A(n_1976),
.B(n_1934),
.Y(n_2354)
);

INVx4_ASAP7_75t_L g2355 ( 
.A(n_1984),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_1999),
.B(n_1951),
.Y(n_2356)
);

NAND2x1p5_ASAP7_75t_L g2357 ( 
.A(n_2191),
.B(n_1938),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_1996),
.Y(n_2358)
);

INVx5_ASAP7_75t_L g2359 ( 
.A(n_1989),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_L g2360 ( 
.A(n_2056),
.B(n_1939),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_1999),
.B(n_1951),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_2297),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2001),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2248),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2001),
.Y(n_2365)
);

NAND2x1p5_ASAP7_75t_L g2366 ( 
.A(n_2191),
.B(n_1938),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2003),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2042),
.B(n_1951),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2003),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2084),
.B(n_1938),
.Y(n_2370)
);

OAI22xp5_ASAP7_75t_L g2371 ( 
.A1(n_2084),
.A2(n_1949),
.B1(n_1954),
.B2(n_1941),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2248),
.Y(n_2372)
);

INVxp33_ASAP7_75t_L g2373 ( 
.A(n_2046),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2256),
.Y(n_2374)
);

NAND3xp33_ASAP7_75t_L g2375 ( 
.A(n_1990),
.B(n_1909),
.C(n_1898),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2080),
.B(n_1773),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2256),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2011),
.B(n_1852),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2260),
.Y(n_2379)
);

INVx3_ASAP7_75t_L g2380 ( 
.A(n_2092),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2004),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2042),
.B(n_1956),
.Y(n_2382)
);

OR2x6_ASAP7_75t_L g2383 ( 
.A(n_2031),
.B(n_1881),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_2221),
.B(n_1962),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2260),
.Y(n_2385)
);

BUFx3_ASAP7_75t_L g2386 ( 
.A(n_2215),
.Y(n_2386)
);

INVx3_ASAP7_75t_L g2387 ( 
.A(n_2092),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_2149),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2004),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2263),
.Y(n_2390)
);

HB1xp67_ASAP7_75t_L g2391 ( 
.A(n_2222),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2080),
.B(n_1775),
.Y(n_2392)
);

CKINVDCx20_ASAP7_75t_R g2393 ( 
.A(n_2297),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2263),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_2311),
.B(n_2250),
.Y(n_2395)
);

AOI22xp33_ASAP7_75t_L g2396 ( 
.A1(n_1981),
.A2(n_735),
.B1(n_743),
.B2(n_734),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2024),
.Y(n_2397)
);

BUFx10_ASAP7_75t_L g2398 ( 
.A(n_2115),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2027),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2034),
.Y(n_2400)
);

AND2x6_ASAP7_75t_L g2401 ( 
.A(n_2089),
.B(n_1877),
.Y(n_2401)
);

BUFx3_ASAP7_75t_L g2402 ( 
.A(n_2007),
.Y(n_2402)
);

INVx1_ASAP7_75t_SL g2403 ( 
.A(n_2119),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2006),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_1977),
.Y(n_2405)
);

AO22x1_ASAP7_75t_L g2406 ( 
.A1(n_2311),
.A2(n_2243),
.B1(n_2210),
.B2(n_2227),
.Y(n_2406)
);

INVx4_ASAP7_75t_L g2407 ( 
.A(n_1984),
.Y(n_2407)
);

CKINVDCx20_ASAP7_75t_R g2408 ( 
.A(n_2261),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_1980),
.Y(n_2409)
);

AOI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_2145),
.A2(n_1954),
.B1(n_1949),
.B2(n_1889),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_1990),
.B(n_1775),
.Y(n_2411)
);

INVx2_ASAP7_75t_SL g2412 ( 
.A(n_2302),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_1986),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2006),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_2314),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1993),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_L g2417 ( 
.A(n_2108),
.B(n_1956),
.Y(n_2417)
);

INVx3_ASAP7_75t_L g2418 ( 
.A(n_2149),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2302),
.B(n_1956),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2097),
.B(n_1785),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_2149),
.Y(n_2421)
);

AND2x6_ASAP7_75t_L g2422 ( 
.A(n_2089),
.B(n_1884),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_1995),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_1997),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2306),
.B(n_1958),
.Y(n_2425)
);

OAI22xp33_ASAP7_75t_L g2426 ( 
.A1(n_2197),
.A2(n_1938),
.B1(n_1868),
.B2(n_1961),
.Y(n_2426)
);

BUFx3_ASAP7_75t_L g2427 ( 
.A(n_2246),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2013),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_2156),
.B(n_1958),
.Y(n_2429)
);

AND2x6_ASAP7_75t_L g2430 ( 
.A(n_1991),
.B(n_1884),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2000),
.Y(n_2431)
);

NAND2x1p5_ASAP7_75t_L g2432 ( 
.A(n_2191),
.B(n_1935),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2306),
.B(n_1958),
.Y(n_2433)
);

INVx5_ASAP7_75t_L g2434 ( 
.A(n_1991),
.Y(n_2434)
);

AND3x1_ASAP7_75t_L g2435 ( 
.A(n_2243),
.B(n_1962),
.C(n_1944),
.Y(n_2435)
);

AOI22xp33_ASAP7_75t_L g2436 ( 
.A1(n_1981),
.A2(n_743),
.B1(n_744),
.B2(n_735),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2046),
.B(n_2070),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2008),
.Y(n_2438)
);

AND2x2_ASAP7_75t_SL g2439 ( 
.A(n_2227),
.B(n_1693),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2013),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2070),
.B(n_1913),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2097),
.B(n_2201),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_SL g2443 ( 
.A(n_2028),
.B(n_1935),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2201),
.B(n_1785),
.Y(n_2444)
);

BUFx10_ASAP7_75t_L g2445 ( 
.A(n_2210),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_L g2446 ( 
.A(n_2238),
.B(n_1942),
.Y(n_2446)
);

NOR2xp33_ASAP7_75t_L g2447 ( 
.A(n_2053),
.B(n_1946),
.Y(n_2447)
);

HB1xp67_ASAP7_75t_L g2448 ( 
.A(n_2099),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_SL g2449 ( 
.A(n_2032),
.B(n_1950),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_L g2450 ( 
.A(n_2314),
.Y(n_2450)
);

OR2x6_ASAP7_75t_L g2451 ( 
.A(n_2029),
.B(n_1881),
.Y(n_2451)
);

INVx4_ASAP7_75t_L g2452 ( 
.A(n_1984),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2014),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2014),
.Y(n_2454)
);

AND2x4_ASAP7_75t_L g2455 ( 
.A(n_2112),
.B(n_2307),
.Y(n_2455)
);

OR2x2_ASAP7_75t_L g2456 ( 
.A(n_2072),
.B(n_1924),
.Y(n_2456)
);

NOR2xp33_ASAP7_75t_L g2457 ( 
.A(n_2169),
.B(n_1948),
.Y(n_2457)
);

AND2x4_ASAP7_75t_L g2458 ( 
.A(n_2112),
.B(n_1886),
.Y(n_2458)
);

BUFx6f_ASAP7_75t_L g2459 ( 
.A(n_2314),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_1983),
.B(n_1789),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2017),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2170),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2009),
.Y(n_2463)
);

INVx3_ASAP7_75t_L g2464 ( 
.A(n_1985),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_2112),
.B(n_1886),
.Y(n_2465)
);

INVx3_ASAP7_75t_L g2466 ( 
.A(n_1985),
.Y(n_2466)
);

BUFx3_ASAP7_75t_L g2467 ( 
.A(n_2207),
.Y(n_2467)
);

INVx4_ASAP7_75t_L g2468 ( 
.A(n_1985),
.Y(n_2468)
);

INVx3_ASAP7_75t_L g2469 ( 
.A(n_1985),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2078),
.B(n_1913),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2242),
.B(n_1789),
.Y(n_2471)
);

NOR2xp33_ASAP7_75t_L g2472 ( 
.A(n_2242),
.B(n_1953),
.Y(n_2472)
);

BUFx3_ASAP7_75t_L g2473 ( 
.A(n_2207),
.Y(n_2473)
);

BUFx10_ASAP7_75t_L g2474 ( 
.A(n_2115),
.Y(n_2474)
);

CKINVDCx5p33_ASAP7_75t_R g2475 ( 
.A(n_2309),
.Y(n_2475)
);

INVx4_ASAP7_75t_L g2476 ( 
.A(n_2025),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2015),
.Y(n_2477)
);

INVx3_ASAP7_75t_L g2478 ( 
.A(n_2025),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_2314),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2017),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2018),
.Y(n_2481)
);

CKINVDCx8_ASAP7_75t_R g2482 ( 
.A(n_2071),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_2309),
.Y(n_2483)
);

INVx6_ASAP7_75t_L g2484 ( 
.A(n_1998),
.Y(n_2484)
);

AND2x4_ASAP7_75t_L g2485 ( 
.A(n_2307),
.B(n_1887),
.Y(n_2485)
);

INVx3_ASAP7_75t_L g2486 ( 
.A(n_2025),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2271),
.B(n_1793),
.Y(n_2487)
);

OAI22xp5_ASAP7_75t_L g2488 ( 
.A1(n_1982),
.A2(n_1957),
.B1(n_1914),
.B2(n_1915),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2078),
.B(n_1913),
.Y(n_2489)
);

INVx1_ASAP7_75t_SL g2490 ( 
.A(n_2111),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2018),
.Y(n_2491)
);

BUFx3_ASAP7_75t_L g2492 ( 
.A(n_2025),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2271),
.B(n_1793),
.Y(n_2493)
);

INVxp67_ASAP7_75t_SL g2494 ( 
.A(n_2035),
.Y(n_2494)
);

NOR2xp33_ASAP7_75t_L g2495 ( 
.A(n_2299),
.B(n_1889),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2231),
.B(n_1935),
.Y(n_2496)
);

AND2x6_ASAP7_75t_L g2497 ( 
.A(n_1991),
.B(n_1887),
.Y(n_2497)
);

AND2x2_ASAP7_75t_SL g2498 ( 
.A(n_2190),
.B(n_1693),
.Y(n_2498)
);

AND2x4_ASAP7_75t_L g2499 ( 
.A(n_2307),
.B(n_1914),
.Y(n_2499)
);

BUFx3_ASAP7_75t_L g2500 ( 
.A(n_2035),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2231),
.B(n_1935),
.Y(n_2501)
);

AO21x2_ASAP7_75t_L g2502 ( 
.A1(n_2145),
.A2(n_1649),
.B(n_1681),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_L g2503 ( 
.A(n_2299),
.B(n_1915),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2021),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2021),
.Y(n_2505)
);

INVx1_ASAP7_75t_SL g2506 ( 
.A(n_2176),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2016),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2093),
.B(n_1950),
.Y(n_2508)
);

INVx4_ASAP7_75t_L g2509 ( 
.A(n_2035),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2040),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2019),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2203),
.B(n_1795),
.Y(n_2512)
);

BUFx8_ASAP7_75t_SL g2513 ( 
.A(n_2115),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_1982),
.B(n_1950),
.Y(n_2514)
);

INVx4_ASAP7_75t_L g2515 ( 
.A(n_2035),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2020),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_1974),
.B(n_1920),
.Y(n_2517)
);

AO21x2_ASAP7_75t_L g2518 ( 
.A1(n_2165),
.A2(n_1850),
.B(n_1798),
.Y(n_2518)
);

BUFx6f_ASAP7_75t_L g2519 ( 
.A(n_2036),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_2218),
.B(n_1920),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2040),
.Y(n_2521)
);

AND2x6_ASAP7_75t_L g2522 ( 
.A(n_1994),
.B(n_1950),
.Y(n_2522)
);

INVx4_ASAP7_75t_L g2523 ( 
.A(n_2036),
.Y(n_2523)
);

NAND2xp33_ASAP7_75t_L g2524 ( 
.A(n_2036),
.B(n_1960),
.Y(n_2524)
);

AOI22xp33_ASAP7_75t_L g2525 ( 
.A1(n_2190),
.A2(n_746),
.B1(n_749),
.B2(n_744),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_1987),
.B(n_1960),
.Y(n_2526)
);

INVx4_ASAP7_75t_L g2527 ( 
.A(n_2036),
.Y(n_2527)
);

BUFx2_ASAP7_75t_L g2528 ( 
.A(n_2181),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2022),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2055),
.Y(n_2530)
);

BUFx3_ASAP7_75t_L g2531 ( 
.A(n_2068),
.Y(n_2531)
);

AND2x6_ASAP7_75t_L g2532 ( 
.A(n_1994),
.B(n_1960),
.Y(n_2532)
);

BUFx4f_ASAP7_75t_L g2533 ( 
.A(n_2071),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2093),
.B(n_2203),
.Y(n_2534)
);

OR2x6_ASAP7_75t_L g2535 ( 
.A(n_2141),
.B(n_1881),
.Y(n_2535)
);

OR2x2_ASAP7_75t_L g2536 ( 
.A(n_2033),
.B(n_1832),
.Y(n_2536)
);

BUFx3_ASAP7_75t_L g2537 ( 
.A(n_2068),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2023),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_1987),
.B(n_1960),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_1992),
.Y(n_2540)
);

AND2x6_ASAP7_75t_L g2541 ( 
.A(n_1994),
.B(n_1961),
.Y(n_2541)
);

OR2x2_ASAP7_75t_L g2542 ( 
.A(n_2198),
.B(n_1809),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_1992),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2055),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2058),
.Y(n_2545)
);

INVx4_ASAP7_75t_SL g2546 ( 
.A(n_2071),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2183),
.B(n_2192),
.Y(n_2547)
);

INVx4_ASAP7_75t_L g2548 ( 
.A(n_2068),
.Y(n_2548)
);

CKINVDCx20_ASAP7_75t_R g2549 ( 
.A(n_2251),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2167),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_SL g2551 ( 
.A(n_2068),
.B(n_1961),
.Y(n_2551)
);

AND2x4_ASAP7_75t_L g2552 ( 
.A(n_2220),
.B(n_1927),
.Y(n_2552)
);

HB1xp67_ASAP7_75t_L g2553 ( 
.A(n_2104),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2173),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_2165),
.B(n_1927),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2175),
.Y(n_2556)
);

AND2x4_ASAP7_75t_L g2557 ( 
.A(n_2224),
.B(n_1881),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2204),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_2166),
.B(n_1891),
.Y(n_2559)
);

BUFx3_ASAP7_75t_L g2560 ( 
.A(n_2081),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2058),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_SL g2562 ( 
.A(n_2081),
.B(n_1961),
.Y(n_2562)
);

INVx4_ASAP7_75t_L g2563 ( 
.A(n_2081),
.Y(n_2563)
);

AND2x6_ASAP7_75t_L g2564 ( 
.A(n_2002),
.B(n_1965),
.Y(n_2564)
);

BUFx6f_ASAP7_75t_L g2565 ( 
.A(n_2081),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2205),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2183),
.B(n_1795),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2059),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_L g2569 ( 
.A(n_2166),
.B(n_1892),
.Y(n_2569)
);

INVx3_ASAP7_75t_L g2570 ( 
.A(n_2160),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2206),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2187),
.B(n_1809),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2059),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2192),
.B(n_1808),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2213),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2214),
.Y(n_2576)
);

BUFx6f_ASAP7_75t_L g2577 ( 
.A(n_2160),
.Y(n_2577)
);

AOI22xp33_ASAP7_75t_L g2578 ( 
.A1(n_2187),
.A2(n_749),
.B1(n_750),
.B2(n_746),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2066),
.Y(n_2579)
);

INVx4_ASAP7_75t_L g2580 ( 
.A(n_2160),
.Y(n_2580)
);

AND2x6_ASAP7_75t_L g2581 ( 
.A(n_2002),
.B(n_1965),
.Y(n_2581)
);

INVx3_ASAP7_75t_L g2582 ( 
.A(n_2160),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2216),
.B(n_1808),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2217),
.Y(n_2584)
);

INVx3_ASAP7_75t_L g2585 ( 
.A(n_2168),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2090),
.Y(n_2586)
);

AND2x4_ASAP7_75t_L g2587 ( 
.A(n_2232),
.B(n_1883),
.Y(n_2587)
);

XOR2xp5_ASAP7_75t_L g2588 ( 
.A(n_2292),
.B(n_1378),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2216),
.B(n_1813),
.Y(n_2589)
);

BUFx6f_ASAP7_75t_L g2590 ( 
.A(n_2168),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2090),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2123),
.B(n_1813),
.Y(n_2592)
);

BUFx6f_ASAP7_75t_L g2593 ( 
.A(n_2168),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2200),
.B(n_1963),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_2168),
.B(n_1883),
.Y(n_2595)
);

INVx4_ASAP7_75t_L g2596 ( 
.A(n_2174),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2094),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2177),
.B(n_1751),
.Y(n_2598)
);

AND2x6_ASAP7_75t_L g2599 ( 
.A(n_2002),
.B(n_1965),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2123),
.B(n_1816),
.Y(n_2600)
);

HB1xp67_ASAP7_75t_L g2601 ( 
.A(n_2104),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2066),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2094),
.Y(n_2603)
);

BUFx2_ASAP7_75t_L g2604 ( 
.A(n_1998),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2103),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2088),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2123),
.B(n_1816),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2103),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2106),
.Y(n_2609)
);

INVx2_ASAP7_75t_SL g2610 ( 
.A(n_2104),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2088),
.Y(n_2611)
);

INVx3_ASAP7_75t_L g2612 ( 
.A(n_2174),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2317),
.Y(n_2613)
);

INVx3_ASAP7_75t_L g2614 ( 
.A(n_2174),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2041),
.B(n_1963),
.Y(n_2615)
);

AND2x4_ASAP7_75t_L g2616 ( 
.A(n_2236),
.B(n_1883),
.Y(n_2616)
);

AND2x4_ASAP7_75t_L g2617 ( 
.A(n_2247),
.B(n_1883),
.Y(n_2617)
);

INVx2_ASAP7_75t_SL g2618 ( 
.A(n_2134),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2106),
.Y(n_2619)
);

INVxp67_ASAP7_75t_L g2620 ( 
.A(n_2270),
.Y(n_2620)
);

INVx4_ASAP7_75t_L g2621 ( 
.A(n_2174),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2172),
.B(n_1897),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_SL g2623 ( 
.A(n_2194),
.B(n_1893),
.Y(n_2623)
);

NOR2xp33_ASAP7_75t_L g2624 ( 
.A(n_2172),
.B(n_1899),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2317),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2113),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2044),
.B(n_1963),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_SL g2628 ( 
.A(n_2194),
.B(n_1893),
.Y(n_2628)
);

AND3x2_ASAP7_75t_L g2629 ( 
.A(n_2178),
.B(n_1952),
.C(n_1906),
.Y(n_2629)
);

INVx3_ASAP7_75t_L g2630 ( 
.A(n_2194),
.Y(n_2630)
);

NOR2xp33_ASAP7_75t_L g2631 ( 
.A(n_2010),
.B(n_1901),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_2194),
.Y(n_2632)
);

NOR2xp33_ASAP7_75t_L g2633 ( 
.A(n_2010),
.B(n_1902),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2189),
.B(n_1846),
.Y(n_2634)
);

OR2x6_ASAP7_75t_L g2635 ( 
.A(n_2147),
.B(n_1893),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2113),
.Y(n_2636)
);

INVx3_ASAP7_75t_L g2637 ( 
.A(n_2234),
.Y(n_2637)
);

AND2x4_ASAP7_75t_L g2638 ( 
.A(n_2193),
.B(n_1893),
.Y(n_2638)
);

BUFx6f_ASAP7_75t_L g2639 ( 
.A(n_2234),
.Y(n_2639)
);

AND2x6_ASAP7_75t_L g2640 ( 
.A(n_2087),
.B(n_1965),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2116),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2116),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2125),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2125),
.Y(n_2644)
);

INVx1_ASAP7_75t_SL g2645 ( 
.A(n_2270),
.Y(n_2645)
);

AND2x6_ASAP7_75t_L g2646 ( 
.A(n_2087),
.B(n_1965),
.Y(n_2646)
);

AND2x4_ASAP7_75t_L g2647 ( 
.A(n_2045),
.B(n_1928),
.Y(n_2647)
);

HB1xp67_ASAP7_75t_L g2648 ( 
.A(n_2184),
.Y(n_2648)
);

INVx4_ASAP7_75t_SL g2649 ( 
.A(n_2071),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2130),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2185),
.B(n_1903),
.Y(n_2651)
);

BUFx6f_ASAP7_75t_L g2652 ( 
.A(n_2234),
.Y(n_2652)
);

BUFx6f_ASAP7_75t_L g2653 ( 
.A(n_2234),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2067),
.B(n_1846),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2130),
.Y(n_2655)
);

AOI22xp33_ASAP7_75t_L g2656 ( 
.A1(n_2087),
.A2(n_751),
.B1(n_754),
.B2(n_750),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2133),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_L g2658 ( 
.A(n_2186),
.B(n_1905),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2133),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2037),
.B(n_1857),
.Y(n_2660)
);

AND2x2_ASAP7_75t_SL g2661 ( 
.A(n_2110),
.B(n_1928),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2146),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2146),
.Y(n_2663)
);

AOI22xp5_ASAP7_75t_L g2664 ( 
.A1(n_2140),
.A2(n_1873),
.B1(n_1870),
.B2(n_1917),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2155),
.Y(n_2665)
);

AND2x4_ASAP7_75t_L g2666 ( 
.A(n_2047),
.B(n_1928),
.Y(n_2666)
);

O2A1O1Ixp33_ASAP7_75t_L g2667 ( 
.A1(n_2442),
.A2(n_2117),
.B(n_2157),
.C(n_2153),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_L g2668 ( 
.A1(n_2656),
.A2(n_2062),
.B1(n_2162),
.B2(n_2158),
.Y(n_2668)
);

BUFx6f_ASAP7_75t_L g2669 ( 
.A(n_2337),
.Y(n_2669)
);

NOR2xp67_ASAP7_75t_SL g2670 ( 
.A(n_2323),
.B(n_1928),
.Y(n_2670)
);

AOI22xp33_ASAP7_75t_L g2671 ( 
.A1(n_2656),
.A2(n_2062),
.B1(n_2164),
.B2(n_2163),
.Y(n_2671)
);

NOR2xp33_ASAP7_75t_L g2672 ( 
.A(n_2395),
.B(n_1667),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2353),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2327),
.B(n_2419),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2425),
.B(n_2255),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2433),
.B(n_2278),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_SL g2677 ( 
.A(n_2368),
.B(n_1908),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2534),
.B(n_2258),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2495),
.B(n_2272),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2572),
.B(n_1947),
.Y(n_2680)
);

BUFx12f_ASAP7_75t_SL g2681 ( 
.A(n_2383),
.Y(n_2681)
);

NAND2xp33_ASAP7_75t_L g2682 ( 
.A(n_2522),
.B(n_2532),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2322),
.Y(n_2683)
);

AOI21x1_ASAP7_75t_L g2684 ( 
.A1(n_2443),
.A2(n_2061),
.B(n_1975),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2495),
.B(n_2262),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_SL g2686 ( 
.A(n_2382),
.B(n_1912),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_L g2687 ( 
.A(n_2395),
.B(n_1709),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2503),
.B(n_2265),
.Y(n_2688)
);

NOR2xp33_ASAP7_75t_L g2689 ( 
.A(n_2326),
.B(n_1947),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_2499),
.B(n_1918),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2503),
.B(n_2252),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2331),
.Y(n_2692)
);

AOI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2406),
.A2(n_2140),
.B1(n_2142),
.B2(n_2050),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2333),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2356),
.B(n_2254),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_SL g2696 ( 
.A(n_2499),
.B(n_1922),
.Y(n_2696)
);

BUFx12f_ASAP7_75t_SL g2697 ( 
.A(n_2383),
.Y(n_2697)
);

INVx8_ASAP7_75t_L g2698 ( 
.A(n_2383),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2361),
.B(n_2249),
.Y(n_2699)
);

CKINVDCx5p33_ASAP7_75t_R g2700 ( 
.A(n_2332),
.Y(n_2700)
);

OAI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_2412),
.A2(n_2120),
.B1(n_2100),
.B2(n_2048),
.Y(n_2701)
);

BUFx3_ASAP7_75t_L g2702 ( 
.A(n_2341),
.Y(n_2702)
);

AOI21xp5_ASAP7_75t_L g2703 ( 
.A1(n_2321),
.A2(n_2274),
.B(n_2086),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2347),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2364),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2472),
.B(n_2360),
.Y(n_2706)
);

INVx5_ASAP7_75t_L g2707 ( 
.A(n_2522),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2499),
.B(n_2496),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2472),
.B(n_2301),
.Y(n_2709)
);

NOR2xp33_ASAP7_75t_L g2710 ( 
.A(n_2326),
.B(n_1926),
.Y(n_2710)
);

AOI22xp5_ASAP7_75t_L g2711 ( 
.A1(n_2437),
.A2(n_2142),
.B1(n_2050),
.B2(n_2098),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2360),
.B(n_2253),
.Y(n_2712)
);

OAI22xp5_ASAP7_75t_L g2713 ( 
.A1(n_2439),
.A2(n_2132),
.B1(n_2101),
.B2(n_2180),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2354),
.B(n_2266),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2354),
.B(n_2267),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2417),
.B(n_2303),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2417),
.B(n_2429),
.Y(n_2717)
);

INVx2_ASAP7_75t_SL g2718 ( 
.A(n_2343),
.Y(n_2718)
);

AOI22xp5_ASAP7_75t_L g2719 ( 
.A1(n_2631),
.A2(n_2098),
.B1(n_2118),
.B2(n_2030),
.Y(n_2719)
);

OR2x2_ASAP7_75t_L g2720 ( 
.A(n_2378),
.B(n_1751),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_SL g2721 ( 
.A(n_2501),
.B(n_1709),
.Y(n_2721)
);

INVx2_ASAP7_75t_SL g2722 ( 
.A(n_2462),
.Y(n_2722)
);

AOI22xp33_ASAP7_75t_L g2723 ( 
.A1(n_2525),
.A2(n_2026),
.B1(n_2161),
.B2(n_2155),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2429),
.B(n_2287),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_SL g2725 ( 
.A(n_2508),
.B(n_1734),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2372),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_SL g2727 ( 
.A(n_2455),
.B(n_1734),
.Y(n_2727)
);

NOR2xp67_ASAP7_75t_L g2728 ( 
.A(n_2375),
.B(n_1749),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2559),
.B(n_2289),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2353),
.Y(n_2730)
);

OAI22xp33_ASAP7_75t_L g2731 ( 
.A1(n_2320),
.A2(n_2057),
.B1(n_2060),
.B2(n_2051),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2358),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2559),
.B(n_2269),
.Y(n_2733)
);

AOI21xp5_ASAP7_75t_L g2734 ( 
.A1(n_2321),
.A2(n_2086),
.B(n_2182),
.Y(n_2734)
);

AOI22xp5_ASAP7_75t_L g2735 ( 
.A1(n_2631),
.A2(n_2118),
.B1(n_2131),
.B2(n_2030),
.Y(n_2735)
);

INVx2_ASAP7_75t_SL g2736 ( 
.A(n_2462),
.Y(n_2736)
);

OAI22xp33_ASAP7_75t_L g2737 ( 
.A1(n_2512),
.A2(n_2065),
.B1(n_2069),
.B2(n_2063),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2569),
.B(n_2264),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2569),
.B(n_2288),
.Y(n_2739)
);

NOR2xp33_ASAP7_75t_L g2740 ( 
.A(n_2373),
.B(n_1749),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_SL g2741 ( 
.A(n_2455),
.B(n_1853),
.Y(n_2741)
);

NOR2xp33_ASAP7_75t_L g2742 ( 
.A(n_2373),
.B(n_2043),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2374),
.Y(n_2743)
);

NOR2xp33_ASAP7_75t_L g2744 ( 
.A(n_2324),
.B(n_2054),
.Y(n_2744)
);

AOI22xp33_ASAP7_75t_L g2745 ( 
.A1(n_2525),
.A2(n_2171),
.B1(n_2179),
.B2(n_2161),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2622),
.B(n_2304),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2622),
.B(n_2293),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2441),
.B(n_1911),
.Y(n_2748)
);

NAND3xp33_ASAP7_75t_L g2749 ( 
.A(n_2517),
.B(n_1988),
.C(n_1971),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2358),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2624),
.B(n_2295),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2363),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2624),
.B(n_2312),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2470),
.B(n_2298),
.Y(n_2754)
);

AND2x2_ASAP7_75t_SL g2755 ( 
.A(n_2439),
.B(n_2237),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2377),
.Y(n_2756)
);

O2A1O1Ixp33_ASAP7_75t_L g2757 ( 
.A1(n_2411),
.A2(n_2315),
.B(n_2318),
.C(n_2316),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2363),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2489),
.B(n_2074),
.Y(n_2759)
);

A2O1A1Ixp33_ASAP7_75t_L g2760 ( 
.A1(n_2555),
.A2(n_2076),
.B(n_2077),
.C(n_2075),
.Y(n_2760)
);

INVx8_ASAP7_75t_L g2761 ( 
.A(n_2401),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2376),
.B(n_2079),
.Y(n_2762)
);

OAI22xp33_ASAP7_75t_L g2763 ( 
.A1(n_2410),
.A2(n_2085),
.B1(n_2096),
.B2(n_2082),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2392),
.B(n_2107),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2379),
.Y(n_2765)
);

NAND2x1_ASAP7_75t_L g2766 ( 
.A(n_2329),
.B(n_2180),
.Y(n_2766)
);

AOI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2633),
.A2(n_2131),
.B1(n_2305),
.B2(n_2239),
.Y(n_2767)
);

INVxp67_ASAP7_75t_L g2768 ( 
.A(n_2528),
.Y(n_2768)
);

INVx2_ASAP7_75t_SL g2769 ( 
.A(n_2403),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2420),
.B(n_2109),
.Y(n_2770)
);

BUFx3_ASAP7_75t_L g2771 ( 
.A(n_2386),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2365),
.Y(n_2772)
);

NOR2xp67_ASAP7_75t_L g2773 ( 
.A(n_2332),
.B(n_1853),
.Y(n_2773)
);

INVxp67_ASAP7_75t_L g2774 ( 
.A(n_2391),
.Y(n_2774)
);

OAI22xp5_ASAP7_75t_L g2775 ( 
.A1(n_2498),
.A2(n_2199),
.B1(n_2211),
.B2(n_2180),
.Y(n_2775)
);

O2A1O1Ixp33_ASAP7_75t_L g2776 ( 
.A1(n_2371),
.A2(n_2121),
.B(n_2128),
.C(n_2124),
.Y(n_2776)
);

NOR2xp33_ASAP7_75t_L g2777 ( 
.A(n_2517),
.B(n_1865),
.Y(n_2777)
);

AOI22xp5_ASAP7_75t_L g2778 ( 
.A1(n_2633),
.A2(n_2135),
.B1(n_2138),
.B2(n_2129),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2365),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_SL g2780 ( 
.A(n_2455),
.B(n_1865),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_SL g2781 ( 
.A(n_2426),
.B(n_1888),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2385),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2390),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2471),
.B(n_2139),
.Y(n_2784)
);

INVx1_ASAP7_75t_SL g2785 ( 
.A(n_2506),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2394),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_L g2787 ( 
.A(n_2490),
.B(n_1888),
.Y(n_2787)
);

AND2x4_ASAP7_75t_L g2788 ( 
.A(n_2346),
.B(n_2143),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2456),
.B(n_1904),
.Y(n_2789)
);

O2A1O1Ixp33_ASAP7_75t_L g2790 ( 
.A1(n_2460),
.A2(n_2148),
.B(n_2151),
.C(n_2144),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_L g2791 ( 
.A(n_2446),
.B(n_1904),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2487),
.B(n_2195),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2493),
.B(n_2195),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2555),
.B(n_2195),
.Y(n_2794)
);

NOR2xp33_ASAP7_75t_L g2795 ( 
.A(n_2446),
.B(n_1907),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2540),
.Y(n_2796)
);

CKINVDCx5p33_ASAP7_75t_R g2797 ( 
.A(n_2393),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2543),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2594),
.B(n_2615),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2648),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_L g2801 ( 
.A(n_2445),
.B(n_1907),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2648),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2627),
.B(n_2245),
.Y(n_2803)
);

OAI21xp5_ASAP7_75t_L g2804 ( 
.A1(n_2498),
.A2(n_2152),
.B(n_2188),
.Y(n_2804)
);

OAI22xp5_ASAP7_75t_SL g2805 ( 
.A1(n_2408),
.A2(n_2154),
.B1(n_2083),
.B2(n_2005),
.Y(n_2805)
);

AOI22xp5_ASAP7_75t_L g2806 ( 
.A1(n_2435),
.A2(n_2245),
.B1(n_1940),
.B2(n_2127),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2586),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_SL g2808 ( 
.A(n_2426),
.B(n_1940),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2591),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2651),
.B(n_2245),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2651),
.B(n_2126),
.Y(n_2811)
);

INVx2_ASAP7_75t_SL g2812 ( 
.A(n_2598),
.Y(n_2812)
);

AND2x6_ASAP7_75t_SL g2813 ( 
.A(n_2635),
.B(n_1968),
.Y(n_2813)
);

AOI22xp33_ASAP7_75t_SL g2814 ( 
.A1(n_2661),
.A2(n_1764),
.B1(n_1867),
.B2(n_2284),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_SL g2815 ( 
.A(n_2638),
.B(n_2257),
.Y(n_2815)
);

NOR2xp67_ASAP7_75t_L g2816 ( 
.A(n_2620),
.B(n_1971),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2658),
.B(n_2134),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2658),
.B(n_2134),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2445),
.B(n_1969),
.Y(n_2819)
);

HB1xp67_ASAP7_75t_L g2820 ( 
.A(n_2391),
.Y(n_2820)
);

AOI22xp33_ASAP7_75t_SL g2821 ( 
.A1(n_2661),
.A2(n_1867),
.B1(n_2073),
.B2(n_1998),
.Y(n_2821)
);

OAI221xp5_ASAP7_75t_L g2822 ( 
.A1(n_2664),
.A2(n_2225),
.B1(n_2457),
.B2(n_2447),
.C(n_2578),
.Y(n_2822)
);

NAND2xp33_ASAP7_75t_L g2823 ( 
.A(n_2522),
.B(n_2237),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2444),
.B(n_2071),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2367),
.Y(n_2825)
);

NAND2xp33_ASAP7_75t_L g2826 ( 
.A(n_2522),
.B(n_2237),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_SL g2827 ( 
.A(n_2638),
.B(n_2150),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2660),
.B(n_2102),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_SL g2829 ( 
.A(n_2638),
.B(n_2196),
.Y(n_2829)
);

AND2x4_ASAP7_75t_L g2830 ( 
.A(n_2346),
.B(n_2102),
.Y(n_2830)
);

AOI21xp5_ASAP7_75t_L g2831 ( 
.A1(n_2321),
.A2(n_2086),
.B(n_2235),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2634),
.B(n_2102),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2597),
.Y(n_2833)
);

INVx2_ASAP7_75t_SL g2834 ( 
.A(n_2384),
.Y(n_2834)
);

O2A1O1Ixp5_ASAP7_75t_L g2835 ( 
.A1(n_2443),
.A2(n_2449),
.B(n_2370),
.C(n_2514),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2367),
.Y(n_2836)
);

O2A1O1Ixp33_ASAP7_75t_L g2837 ( 
.A1(n_2449),
.A2(n_2171),
.B(n_2208),
.C(n_2179),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2603),
.Y(n_2838)
);

AOI22xp5_ASAP7_75t_L g2839 ( 
.A1(n_2618),
.A2(n_2102),
.B1(n_2136),
.B2(n_1911),
.Y(n_2839)
);

INVx2_ASAP7_75t_SL g2840 ( 
.A(n_2427),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2369),
.Y(n_2841)
);

CKINVDCx5p33_ASAP7_75t_R g2842 ( 
.A(n_2393),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_SL g2843 ( 
.A(n_2647),
.B(n_2237),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2605),
.Y(n_2844)
);

AOI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_2666),
.A2(n_2102),
.B1(n_2122),
.B2(n_1703),
.Y(n_2845)
);

NOR2xp33_ASAP7_75t_L g2846 ( 
.A(n_2447),
.B(n_1970),
.Y(n_2846)
);

AND2x4_ASAP7_75t_L g2847 ( 
.A(n_2402),
.B(n_2102),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2608),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2609),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2619),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2542),
.B(n_1703),
.Y(n_2851)
);

NOR2xp33_ASAP7_75t_L g2852 ( 
.A(n_2457),
.B(n_1973),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2654),
.B(n_2208),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2550),
.B(n_2209),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2554),
.B(n_2209),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2556),
.B(n_2212),
.Y(n_2856)
);

NAND2xp33_ASAP7_75t_SL g2857 ( 
.A(n_2475),
.B(n_2105),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2558),
.B(n_2212),
.Y(n_2858)
);

NOR2xp67_ASAP7_75t_L g2859 ( 
.A(n_2475),
.B(n_2483),
.Y(n_2859)
);

INVx2_ASAP7_75t_SL g2860 ( 
.A(n_2427),
.Y(n_2860)
);

INVxp67_ASAP7_75t_L g2861 ( 
.A(n_2448),
.Y(n_2861)
);

AOI22xp33_ASAP7_75t_SL g2862 ( 
.A1(n_2635),
.A2(n_2073),
.B1(n_1882),
.B2(n_1845),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2626),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2566),
.B(n_2223),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_SL g2865 ( 
.A(n_2348),
.B(n_1814),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_SL g2866 ( 
.A(n_2647),
.B(n_2273),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_L g2867 ( 
.A(n_2448),
.B(n_2137),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2571),
.B(n_2219),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2575),
.B(n_2219),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2576),
.B(n_2223),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2584),
.B(n_2228),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2397),
.B(n_2228),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2399),
.B(n_2273),
.Y(n_2873)
);

AND2x4_ASAP7_75t_SL g2874 ( 
.A(n_2398),
.B(n_1801),
.Y(n_2874)
);

NAND2xp33_ASAP7_75t_L g2875 ( 
.A(n_2522),
.B(n_2273),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2400),
.B(n_2273),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_L g2877 ( 
.A(n_2645),
.B(n_2290),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2405),
.B(n_2275),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2369),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2409),
.B(n_2275),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2413),
.B(n_2275),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2416),
.B(n_2275),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2636),
.Y(n_2883)
);

NAND2xp33_ASAP7_75t_L g2884 ( 
.A(n_2532),
.B(n_1797),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2641),
.Y(n_2885)
);

NOR2xp67_ASAP7_75t_L g2886 ( 
.A(n_2483),
.B(n_1741),
.Y(n_2886)
);

AOI22xp33_ASAP7_75t_L g2887 ( 
.A1(n_2396),
.A2(n_754),
.B1(n_755),
.B2(n_751),
.Y(n_2887)
);

AND2x4_ASAP7_75t_L g2888 ( 
.A(n_2402),
.B(n_1741),
.Y(n_2888)
);

AND2x6_ASAP7_75t_SL g2889 ( 
.A(n_2635),
.B(n_1916),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_L g2890 ( 
.A(n_2536),
.B(n_2012),
.Y(n_2890)
);

NOR3xp33_ASAP7_75t_L g2891 ( 
.A(n_2488),
.B(n_1952),
.C(n_1906),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2423),
.B(n_2424),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2381),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2431),
.B(n_2229),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2642),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2438),
.B(n_2229),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2381),
.Y(n_2897)
);

AOI22xp33_ASAP7_75t_L g2898 ( 
.A1(n_2396),
.A2(n_2436),
.B1(n_2578),
.B2(n_2336),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_SL g2899 ( 
.A(n_2647),
.B(n_2012),
.Y(n_2899)
);

OAI21xp33_ASAP7_75t_L g2900 ( 
.A1(n_2436),
.A2(n_1849),
.B(n_1797),
.Y(n_2900)
);

OR2x2_ASAP7_75t_L g2901 ( 
.A(n_2345),
.B(n_1841),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2389),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2463),
.B(n_2233),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2477),
.B(n_2233),
.Y(n_2904)
);

BUFx3_ASAP7_75t_L g2905 ( 
.A(n_2386),
.Y(n_2905)
);

BUFx6f_ASAP7_75t_L g2906 ( 
.A(n_2337),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2507),
.B(n_2233),
.Y(n_2907)
);

INVxp67_ASAP7_75t_L g2908 ( 
.A(n_2553),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2511),
.B(n_2244),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_2345),
.B(n_1841),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_SL g2911 ( 
.A(n_2666),
.B(n_1849),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2516),
.B(n_2199),
.Y(n_2912)
);

NOR2xp67_ASAP7_75t_L g2913 ( 
.A(n_2348),
.B(n_1857),
.Y(n_2913)
);

CKINVDCx5p33_ASAP7_75t_R g2914 ( 
.A(n_2362),
.Y(n_2914)
);

BUFx6f_ASAP7_75t_L g2915 ( 
.A(n_2337),
.Y(n_2915)
);

AOI22xp33_ASAP7_75t_L g2916 ( 
.A1(n_2336),
.A2(n_759),
.B1(n_766),
.B2(n_755),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_SL g2917 ( 
.A(n_2666),
.B(n_1878),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2389),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2643),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2650),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2655),
.Y(n_2921)
);

AOI22xp33_ASAP7_75t_L g2922 ( 
.A1(n_2547),
.A2(n_766),
.B1(n_768),
.B2(n_759),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2657),
.Y(n_2923)
);

AO221x1_ASAP7_75t_L g2924 ( 
.A1(n_2464),
.A2(n_1848),
.B1(n_1845),
.B2(n_771),
.C(n_778),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2553),
.B(n_1848),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_SL g2926 ( 
.A(n_2520),
.B(n_1878),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2529),
.B(n_2259),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_SL g2928 ( 
.A(n_2520),
.B(n_2073),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2538),
.B(n_2199),
.Y(n_2929)
);

OAI22x1_ASAP7_75t_SL g2930 ( 
.A1(n_2408),
.A2(n_1825),
.B1(n_1838),
.B2(n_1801),
.Y(n_2930)
);

INVx2_ASAP7_75t_SL g2931 ( 
.A(n_2362),
.Y(n_2931)
);

BUFx6f_ASAP7_75t_L g2932 ( 
.A(n_2337),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2404),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2663),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2613),
.Y(n_2935)
);

NOR2xp67_ASAP7_75t_SL g2936 ( 
.A(n_2482),
.B(n_2296),
.Y(n_2936)
);

NAND3xp33_ASAP7_75t_L g2937 ( 
.A(n_2601),
.B(n_1406),
.C(n_1393),
.Y(n_2937)
);

OR2x6_ASAP7_75t_L g2938 ( 
.A(n_2484),
.B(n_2330),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2592),
.B(n_2229),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2600),
.B(n_2211),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2404),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_SL g2942 ( 
.A(n_2352),
.B(n_1825),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2607),
.B(n_2244),
.Y(n_2943)
);

NAND2x1p5_ASAP7_75t_L g2944 ( 
.A(n_2338),
.B(n_2211),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2520),
.B(n_2259),
.Y(n_2945)
);

NOR2xp33_ASAP7_75t_L g2946 ( 
.A(n_2601),
.B(n_1838),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2613),
.Y(n_2947)
);

A2O1A1Ixp33_ASAP7_75t_L g2948 ( 
.A1(n_2552),
.A2(n_2259),
.B(n_2281),
.C(n_2244),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2552),
.B(n_2281),
.Y(n_2949)
);

NOR2xp33_ASAP7_75t_L g2950 ( 
.A(n_2552),
.B(n_1916),
.Y(n_2950)
);

AOI22xp33_ASAP7_75t_L g2951 ( 
.A1(n_2625),
.A2(n_771),
.B1(n_775),
.B2(n_768),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2625),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_SL g2953 ( 
.A(n_2352),
.B(n_1923),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2644),
.Y(n_2954)
);

BUFx6f_ASAP7_75t_SL g2955 ( 
.A(n_2535),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2458),
.B(n_2281),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2458),
.B(n_2285),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2414),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2610),
.B(n_1923),
.Y(n_2959)
);

INVxp67_ASAP7_75t_L g2960 ( 
.A(n_2557),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2414),
.Y(n_2961)
);

BUFx6f_ASAP7_75t_L g2962 ( 
.A(n_2338),
.Y(n_2962)
);

AOI22xp5_ASAP7_75t_L g2963 ( 
.A1(n_2458),
.A2(n_1933),
.B1(n_1408),
.B2(n_1428),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2428),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2428),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_SL g2966 ( 
.A(n_2557),
.B(n_2587),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2465),
.B(n_2285),
.Y(n_2967)
);

BUFx3_ASAP7_75t_L g2968 ( 
.A(n_2484),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2440),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2892),
.Y(n_2970)
);

INVx4_ASAP7_75t_L g2971 ( 
.A(n_2698),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2807),
.Y(n_2972)
);

CKINVDCx20_ASAP7_75t_R g2973 ( 
.A(n_2797),
.Y(n_2973)
);

INVx3_ASAP7_75t_L g2974 ( 
.A(n_2761),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2809),
.Y(n_2975)
);

AND2x6_ASAP7_75t_SL g2976 ( 
.A(n_2801),
.B(n_2535),
.Y(n_2976)
);

INVx5_ASAP7_75t_L g2977 ( 
.A(n_2698),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2674),
.B(n_2532),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_R g2979 ( 
.A(n_2700),
.B(n_1933),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2833),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2838),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2673),
.Y(n_2982)
);

INVx3_ASAP7_75t_L g2983 ( 
.A(n_2761),
.Y(n_2983)
);

NAND2x1p5_ASAP7_75t_L g2984 ( 
.A(n_2707),
.B(n_2492),
.Y(n_2984)
);

AND3x2_ASAP7_75t_SL g2985 ( 
.A(n_2930),
.B(n_2588),
.C(n_2629),
.Y(n_2985)
);

HB1xp67_ASAP7_75t_L g2986 ( 
.A(n_2718),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_SL g2987 ( 
.A(n_2777),
.B(n_2557),
.Y(n_2987)
);

OAI22xp5_ASAP7_75t_L g2988 ( 
.A1(n_2706),
.A2(n_2535),
.B1(n_2451),
.B2(n_2366),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_SL g2989 ( 
.A(n_2777),
.B(n_2587),
.Y(n_2989)
);

INVxp67_ASAP7_75t_L g2990 ( 
.A(n_2720),
.Y(n_2990)
);

AND2x4_ASAP7_75t_L g2991 ( 
.A(n_2938),
.B(n_2485),
.Y(n_2991)
);

AND2x6_ASAP7_75t_SL g2992 ( 
.A(n_2672),
.B(n_2687),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_SL g2993 ( 
.A(n_2791),
.B(n_2587),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2844),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_SL g2995 ( 
.A(n_2795),
.B(n_2616),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2848),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2811),
.B(n_2532),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2717),
.B(n_2532),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2730),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2849),
.Y(n_3000)
);

CKINVDCx5p33_ASAP7_75t_R g3001 ( 
.A(n_2842),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2732),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_SL g3003 ( 
.A(n_2689),
.B(n_2710),
.Y(n_3003)
);

NOR2x2_ASAP7_75t_L g3004 ( 
.A(n_2938),
.B(n_2451),
.Y(n_3004)
);

AOI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2744),
.A2(n_2822),
.B1(n_2742),
.B2(n_2877),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2712),
.B(n_2616),
.Y(n_3006)
);

INVx8_ASAP7_75t_L g3007 ( 
.A(n_2698),
.Y(n_3007)
);

AOI21xp5_ASAP7_75t_L g3008 ( 
.A1(n_2823),
.A2(n_2524),
.B(n_2334),
.Y(n_3008)
);

BUFx4f_ASAP7_75t_L g3009 ( 
.A(n_2938),
.Y(n_3009)
);

INVx1_ASAP7_75t_SL g3010 ( 
.A(n_2785),
.Y(n_3010)
);

AND2x6_ASAP7_75t_SL g3011 ( 
.A(n_2890),
.B(n_2451),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2850),
.Y(n_3012)
);

BUFx4f_ASAP7_75t_L g3013 ( 
.A(n_2874),
.Y(n_3013)
);

AOI22xp33_ASAP7_75t_L g3014 ( 
.A1(n_2744),
.A2(n_2485),
.B1(n_2465),
.B2(n_2616),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2863),
.Y(n_3015)
);

NAND2xp33_ASAP7_75t_L g3016 ( 
.A(n_2900),
.B(n_2432),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2714),
.B(n_2715),
.Y(n_3017)
);

AND2x2_ASAP7_75t_L g3018 ( 
.A(n_2748),
.B(n_2617),
.Y(n_3018)
);

CKINVDCx20_ASAP7_75t_R g3019 ( 
.A(n_2914),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2709),
.B(n_2617),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2710),
.B(n_2617),
.Y(n_3021)
);

INVx6_ASAP7_75t_L g3022 ( 
.A(n_2702),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2750),
.Y(n_3023)
);

AOI22xp33_ASAP7_75t_L g3024 ( 
.A1(n_2742),
.A2(n_2485),
.B1(n_2465),
.B2(n_2339),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2883),
.Y(n_3025)
);

HB1xp67_ASAP7_75t_L g3026 ( 
.A(n_2769),
.Y(n_3026)
);

INVx3_ASAP7_75t_L g3027 ( 
.A(n_2761),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_SL g3028 ( 
.A(n_2689),
.B(n_2340),
.Y(n_3028)
);

AOI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2826),
.A2(n_2524),
.B(n_2334),
.Y(n_3029)
);

INVx2_ASAP7_75t_SL g3030 ( 
.A(n_2771),
.Y(n_3030)
);

INVxp67_ASAP7_75t_L g3031 ( 
.A(n_2812),
.Y(n_3031)
);

AND2x4_ASAP7_75t_L g3032 ( 
.A(n_2788),
.B(n_2339),
.Y(n_3032)
);

BUFx2_ASAP7_75t_SL g3033 ( 
.A(n_2905),
.Y(n_3033)
);

AOI22xp33_ASAP7_75t_L g3034 ( 
.A1(n_2877),
.A2(n_2339),
.B1(n_2526),
.B2(n_2514),
.Y(n_3034)
);

BUFx3_ASAP7_75t_L g3035 ( 
.A(n_2968),
.Y(n_3035)
);

AND2x2_ASAP7_75t_L g3036 ( 
.A(n_2680),
.B(n_2330),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2752),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2885),
.Y(n_3038)
);

OAI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2898),
.A2(n_2366),
.B1(n_2357),
.B2(n_2432),
.Y(n_3039)
);

AOI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_2851),
.A2(n_2701),
.B1(n_2735),
.B2(n_2719),
.Y(n_3040)
);

BUFx6f_ASAP7_75t_L g3041 ( 
.A(n_2669),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2895),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2758),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2772),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2762),
.B(n_2541),
.Y(n_3045)
);

INVx3_ASAP7_75t_L g3046 ( 
.A(n_2669),
.Y(n_3046)
);

AOI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2875),
.A2(n_2334),
.B(n_2321),
.Y(n_3047)
);

AOI21xp5_ASAP7_75t_L g3048 ( 
.A1(n_2804),
.A2(n_2359),
.B(n_2334),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2779),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2846),
.B(n_1408),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2919),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2920),
.Y(n_3052)
);

INVx6_ASAP7_75t_L g3053 ( 
.A(n_2901),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2925),
.B(n_2467),
.Y(n_3054)
);

NOR3xp33_ASAP7_75t_SL g3055 ( 
.A(n_2749),
.B(n_719),
.C(n_718),
.Y(n_3055)
);

NOR2x2_ASAP7_75t_L g3056 ( 
.A(n_2805),
.B(n_670),
.Y(n_3056)
);

NAND3xp33_ASAP7_75t_SL g3057 ( 
.A(n_2767),
.B(n_1428),
.C(n_1412),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2921),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2867),
.B(n_2467),
.Y(n_3059)
);

BUFx6f_ASAP7_75t_L g3060 ( 
.A(n_2669),
.Y(n_3060)
);

HB1xp67_ASAP7_75t_L g3061 ( 
.A(n_2820),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2825),
.Y(n_3062)
);

AO21x1_ASAP7_75t_L g3063 ( 
.A1(n_2713),
.A2(n_2370),
.B(n_2526),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2923),
.Y(n_3064)
);

INVx4_ASAP7_75t_L g3065 ( 
.A(n_2669),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2934),
.Y(n_3066)
);

BUFx8_ASAP7_75t_L g3067 ( 
.A(n_2955),
.Y(n_3067)
);

AO22x1_ASAP7_75t_L g3068 ( 
.A1(n_2789),
.A2(n_2787),
.B1(n_2852),
.B2(n_2890),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2836),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2764),
.B(n_2541),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2841),
.Y(n_3071)
);

INVx1_ASAP7_75t_SL g3072 ( 
.A(n_2820),
.Y(n_3072)
);

AOI22xp5_ASAP7_75t_L g3073 ( 
.A1(n_2701),
.A2(n_2539),
.B1(n_2623),
.B2(n_2595),
.Y(n_3073)
);

AOI22xp5_ASAP7_75t_L g3074 ( 
.A1(n_2867),
.A2(n_2539),
.B1(n_2623),
.B2(n_2595),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2879),
.Y(n_3075)
);

BUFx6f_ASAP7_75t_L g3076 ( 
.A(n_2906),
.Y(n_3076)
);

INVx2_ASAP7_75t_SL g3077 ( 
.A(n_2722),
.Y(n_3077)
);

BUFx2_ASAP7_75t_L g3078 ( 
.A(n_2768),
.Y(n_3078)
);

NOR2xp33_ASAP7_75t_L g3079 ( 
.A(n_2852),
.B(n_1412),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2893),
.Y(n_3080)
);

BUFx2_ASAP7_75t_L g3081 ( 
.A(n_2768),
.Y(n_3081)
);

NOR2x2_ASAP7_75t_L g3082 ( 
.A(n_2969),
.B(n_2549),
.Y(n_3082)
);

NAND2x1p5_ASAP7_75t_L g3083 ( 
.A(n_2707),
.B(n_2492),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2897),
.Y(n_3084)
);

BUFx6f_ASAP7_75t_L g3085 ( 
.A(n_2906),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2770),
.B(n_2541),
.Y(n_3086)
);

BUFx6f_ASAP7_75t_L g3087 ( 
.A(n_2906),
.Y(n_3087)
);

AND2x4_ASAP7_75t_L g3088 ( 
.A(n_2788),
.B(n_2473),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2817),
.B(n_2473),
.Y(n_3089)
);

AND2x4_ASAP7_75t_L g3090 ( 
.A(n_2966),
.B(n_2500),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2818),
.B(n_2357),
.Y(n_3091)
);

BUFx4f_ASAP7_75t_L g3092 ( 
.A(n_2888),
.Y(n_3092)
);

INVx2_ASAP7_75t_SL g3093 ( 
.A(n_2736),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2902),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2918),
.Y(n_3095)
);

INVx3_ASAP7_75t_L g3096 ( 
.A(n_2906),
.Y(n_3096)
);

BUFx6f_ASAP7_75t_L g3097 ( 
.A(n_2915),
.Y(n_3097)
);

AND2x6_ASAP7_75t_L g3098 ( 
.A(n_2830),
.B(n_2325),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2679),
.B(n_2628),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_SL g3100 ( 
.A(n_2740),
.B(n_2340),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2685),
.B(n_2628),
.Y(n_3101)
);

NAND3xp33_ASAP7_75t_L g3102 ( 
.A(n_2891),
.B(n_2629),
.C(n_2562),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2933),
.Y(n_3103)
);

CKINVDCx20_ASAP7_75t_R g3104 ( 
.A(n_2963),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2941),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_2959),
.B(n_2349),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2688),
.B(n_2567),
.Y(n_3107)
);

AOI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_2810),
.A2(n_2562),
.B1(n_2551),
.B2(n_2502),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_SL g3109 ( 
.A(n_2773),
.B(n_2349),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2958),
.Y(n_3110)
);

AND2x4_ASAP7_75t_L g3111 ( 
.A(n_2840),
.B(n_2860),
.Y(n_3111)
);

CKINVDCx11_ASAP7_75t_R g3112 ( 
.A(n_2889),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_2915),
.Y(n_3113)
);

NAND2x1p5_ASAP7_75t_L g3114 ( 
.A(n_2707),
.B(n_2500),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2691),
.B(n_2574),
.Y(n_3115)
);

NOR3xp33_ASAP7_75t_L g3116 ( 
.A(n_2781),
.B(n_2604),
.C(n_2551),
.Y(n_3116)
);

AND2x4_ASAP7_75t_L g3117 ( 
.A(n_2960),
.B(n_2531),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2729),
.B(n_2583),
.Y(n_3118)
);

CKINVDCx5p33_ASAP7_75t_R g3119 ( 
.A(n_2813),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2961),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2733),
.B(n_2589),
.Y(n_3121)
);

INVx5_ASAP7_75t_L g3122 ( 
.A(n_2915),
.Y(n_3122)
);

NAND3xp33_ASAP7_75t_SL g3123 ( 
.A(n_2806),
.B(n_2549),
.C(n_725),
.Y(n_3123)
);

INVx3_ASAP7_75t_L g3124 ( 
.A(n_2915),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2964),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2965),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2935),
.Y(n_3127)
);

INVx5_ASAP7_75t_L g3128 ( 
.A(n_2932),
.Y(n_3128)
);

CKINVDCx5p33_ASAP7_75t_R g3129 ( 
.A(n_2931),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2738),
.B(n_2541),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_2834),
.B(n_2398),
.Y(n_3131)
);

BUFx2_ASAP7_75t_L g3132 ( 
.A(n_2681),
.Y(n_3132)
);

INVx2_ASAP7_75t_SL g3133 ( 
.A(n_2888),
.Y(n_3133)
);

NOR2xp33_ASAP7_75t_L g3134 ( 
.A(n_2827),
.B(n_2513),
.Y(n_3134)
);

AND2x4_ASAP7_75t_L g3135 ( 
.A(n_2960),
.B(n_2531),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_2808),
.A2(n_2502),
.B1(n_2422),
.B2(n_2401),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2947),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2739),
.B(n_2541),
.Y(n_3138)
);

BUFx2_ASAP7_75t_L g3139 ( 
.A(n_2697),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2952),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2954),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2746),
.B(n_2644),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2747),
.B(n_2659),
.Y(n_3143)
);

BUFx6f_ASAP7_75t_L g3144 ( 
.A(n_2932),
.Y(n_3144)
);

OR2x6_ASAP7_75t_L g3145 ( 
.A(n_2928),
.B(n_2484),
.Y(n_3145)
);

INVx5_ASAP7_75t_L g3146 ( 
.A(n_2932),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2683),
.Y(n_3147)
);

NOR2xp33_ASAP7_75t_L g3148 ( 
.A(n_2829),
.B(n_2513),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_L g3149 ( 
.A(n_2910),
.B(n_2398),
.Y(n_3149)
);

BUFx6f_ASAP7_75t_L g3150 ( 
.A(n_2932),
.Y(n_3150)
);

AOI22xp5_ASAP7_75t_L g3151 ( 
.A1(n_2891),
.A2(n_2422),
.B1(n_2401),
.B2(n_2430),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2751),
.B(n_2659),
.Y(n_3152)
);

CKINVDCx5p33_ASAP7_75t_R g3153 ( 
.A(n_2910),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_SL g3154 ( 
.A(n_2728),
.B(n_2859),
.Y(n_3154)
);

AOI22xp33_ASAP7_75t_L g3155 ( 
.A1(n_2899),
.A2(n_2422),
.B1(n_2401),
.B2(n_2564),
.Y(n_3155)
);

AOI22xp5_ASAP7_75t_L g3156 ( 
.A1(n_2693),
.A2(n_2422),
.B1(n_2401),
.B2(n_2430),
.Y(n_3156)
);

AND2x4_ASAP7_75t_L g3157 ( 
.A(n_2847),
.B(n_2908),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2692),
.Y(n_3158)
);

INVx2_ASAP7_75t_SL g3159 ( 
.A(n_2800),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2753),
.B(n_2662),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2694),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2704),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_SL g3163 ( 
.A(n_2670),
.B(n_2474),
.Y(n_3163)
);

OAI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_2835),
.A2(n_2061),
.B(n_2662),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2705),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2726),
.Y(n_3166)
);

CKINVDCx5p33_ASAP7_75t_R g3167 ( 
.A(n_2946),
.Y(n_3167)
);

BUFx12f_ASAP7_75t_L g3168 ( 
.A(n_2847),
.Y(n_3168)
);

INVx4_ASAP7_75t_L g3169 ( 
.A(n_2962),
.Y(n_3169)
);

INVx3_ASAP7_75t_L g3170 ( 
.A(n_2962),
.Y(n_3170)
);

A2O1A1Ixp33_ASAP7_75t_L g3171 ( 
.A1(n_2711),
.A2(n_2533),
.B(n_2380),
.C(n_2387),
.Y(n_3171)
);

BUFx2_ASAP7_75t_L g3172 ( 
.A(n_2774),
.Y(n_3172)
);

AND2x4_ASAP7_75t_SL g3173 ( 
.A(n_2830),
.B(n_2474),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2743),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2756),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2765),
.Y(n_3176)
);

INVx1_ASAP7_75t_SL g3177 ( 
.A(n_2802),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_SL g3178 ( 
.A(n_2816),
.B(n_2474),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2784),
.B(n_2665),
.Y(n_3179)
);

INVxp67_ASAP7_75t_L g3180 ( 
.A(n_2942),
.Y(n_3180)
);

CKINVDCx5p33_ASAP7_75t_R g3181 ( 
.A(n_2819),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2782),
.Y(n_3182)
);

AND2x4_ASAP7_75t_L g3183 ( 
.A(n_2908),
.B(n_2537),
.Y(n_3183)
);

BUFx2_ASAP7_75t_L g3184 ( 
.A(n_2774),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_SL g3185 ( 
.A(n_2678),
.B(n_2338),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_SL g3186 ( 
.A(n_2953),
.B(n_2338),
.Y(n_3186)
);

INVx3_ASAP7_75t_L g3187 ( 
.A(n_2962),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2783),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2786),
.Y(n_3189)
);

AO21x1_ASAP7_75t_L g3190 ( 
.A1(n_2737),
.A2(n_2159),
.B(n_2280),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2796),
.Y(n_3191)
);

AND2x2_ASAP7_75t_SL g3192 ( 
.A(n_2755),
.B(n_2533),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2798),
.Y(n_3193)
);

INVx3_ASAP7_75t_L g3194 ( 
.A(n_2962),
.Y(n_3194)
);

NOR2xp33_ASAP7_75t_L g3195 ( 
.A(n_2861),
.B(n_2325),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_SL g3196 ( 
.A(n_3005),
.B(n_3003),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_3040),
.B(n_2737),
.Y(n_3197)
);

AND2x2_ASAP7_75t_L g3198 ( 
.A(n_3059),
.B(n_2950),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_SL g3199 ( 
.A(n_3040),
.B(n_2755),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_3017),
.B(n_2695),
.Y(n_3200)
);

NAND2xp33_ASAP7_75t_SL g3201 ( 
.A(n_2979),
.B(n_2955),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_SL g3202 ( 
.A(n_3021),
.B(n_2794),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3068),
.B(n_2699),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2970),
.B(n_2754),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_SL g3205 ( 
.A(n_3181),
.B(n_2821),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_SL g3206 ( 
.A(n_3153),
.B(n_2821),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_SL g3207 ( 
.A(n_3079),
.B(n_2778),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_SL g3208 ( 
.A(n_3050),
.B(n_2862),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_SL g3209 ( 
.A(n_3167),
.B(n_2862),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_3054),
.B(n_2950),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_SL g3211 ( 
.A(n_2993),
.B(n_2721),
.Y(n_3211)
);

NAND2xp33_ASAP7_75t_SL g3212 ( 
.A(n_3019),
.B(n_2936),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_SL g3213 ( 
.A(n_2995),
.B(n_2725),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_SL g3214 ( 
.A(n_3092),
.B(n_2759),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_3092),
.B(n_2675),
.Y(n_3215)
);

NAND2xp33_ASAP7_75t_SL g3216 ( 
.A(n_3129),
.B(n_2898),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_SL g3217 ( 
.A(n_2987),
.B(n_2676),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_SL g3218 ( 
.A(n_2989),
.B(n_2937),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_SL g3219 ( 
.A(n_3020),
.B(n_2716),
.Y(n_3219)
);

NAND2x1p5_ASAP7_75t_L g3220 ( 
.A(n_3009),
.B(n_2707),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_SL g3221 ( 
.A(n_3006),
.B(n_2724),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_3018),
.B(n_2799),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_SL g3223 ( 
.A(n_3014),
.B(n_2731),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_SL g3224 ( 
.A(n_3009),
.B(n_2731),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_SL g3225 ( 
.A(n_3149),
.B(n_2988),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_SL g3226 ( 
.A(n_2988),
.B(n_2790),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2990),
.B(n_2668),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_SL g3228 ( 
.A(n_3028),
.B(n_2790),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_3036),
.B(n_2668),
.Y(n_3229)
);

NAND2xp33_ASAP7_75t_SL g3230 ( 
.A(n_2973),
.B(n_2727),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_SL g3231 ( 
.A(n_3116),
.B(n_2814),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_SL g3232 ( 
.A(n_3024),
.B(n_2814),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_SL g3233 ( 
.A(n_3134),
.B(n_2886),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_SL g3234 ( 
.A(n_3148),
.B(n_2845),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_3089),
.B(n_2671),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_SL g3236 ( 
.A(n_2991),
.B(n_2911),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_SL g3237 ( 
.A(n_2991),
.B(n_2917),
.Y(n_3237)
);

AND2x4_ASAP7_75t_L g3238 ( 
.A(n_2974),
.B(n_2708),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_SL g3239 ( 
.A(n_3100),
.B(n_2741),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_SL g3240 ( 
.A(n_3133),
.B(n_2780),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_SL g3241 ( 
.A(n_3055),
.B(n_2913),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_SL g3242 ( 
.A(n_3010),
.B(n_2926),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_SL g3243 ( 
.A(n_3010),
.B(n_2671),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_SL g3244 ( 
.A(n_3180),
.B(n_2865),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_SL g3245 ( 
.A(n_3072),
.B(n_2763),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_SL g3246 ( 
.A(n_3072),
.B(n_2763),
.Y(n_3246)
);

AND2x2_ASAP7_75t_L g3247 ( 
.A(n_3106),
.B(n_2861),
.Y(n_3247)
);

AND2x4_ASAP7_75t_L g3248 ( 
.A(n_2974),
.B(n_2815),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_SL g3249 ( 
.A(n_3163),
.B(n_3013),
.Y(n_3249)
);

NAND2xp33_ASAP7_75t_SL g3250 ( 
.A(n_2971),
.B(n_2690),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_SL g3251 ( 
.A(n_3163),
.B(n_2803),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_SL g3252 ( 
.A(n_3013),
.B(n_2792),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_SL g3253 ( 
.A(n_2977),
.B(n_2793),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_SL g3254 ( 
.A(n_2977),
.B(n_2677),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_SL g3255 ( 
.A(n_2977),
.B(n_2686),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_SL g3256 ( 
.A(n_3177),
.B(n_2839),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_SL g3257 ( 
.A(n_3177),
.B(n_3091),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_SL g3258 ( 
.A(n_3157),
.B(n_2696),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_SL g3259 ( 
.A(n_3157),
.B(n_2667),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_SL g3260 ( 
.A(n_3192),
.B(n_2667),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_SL g3261 ( 
.A(n_3034),
.B(n_2760),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_3118),
.B(n_2922),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_SL g3263 ( 
.A(n_3186),
.B(n_3102),
.Y(n_3263)
);

NAND2xp33_ASAP7_75t_SL g3264 ( 
.A(n_2971),
.B(n_2342),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_SL g3265 ( 
.A(n_3102),
.B(n_2857),
.Y(n_3265)
);

NAND2xp33_ASAP7_75t_SL g3266 ( 
.A(n_3001),
.B(n_2342),
.Y(n_3266)
);

NAND2xp33_ASAP7_75t_SL g3267 ( 
.A(n_3119),
.B(n_2342),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_SL g3268 ( 
.A(n_3074),
.B(n_2776),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_3121),
.B(n_2922),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_SL g3270 ( 
.A(n_3074),
.B(n_2776),
.Y(n_3270)
);

NAND2xp33_ASAP7_75t_SL g3271 ( 
.A(n_3109),
.B(n_2342),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_2992),
.B(n_2853),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_SL g3273 ( 
.A(n_3183),
.B(n_2757),
.Y(n_3273)
);

AND2x2_ASAP7_75t_L g3274 ( 
.A(n_3032),
.B(n_2924),
.Y(n_3274)
);

NAND2xp33_ASAP7_75t_SL g3275 ( 
.A(n_3030),
.B(n_2350),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_SL g3276 ( 
.A(n_3183),
.B(n_2757),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_SL g3277 ( 
.A(n_3172),
.B(n_2916),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_SL g3278 ( 
.A(n_3184),
.B(n_2916),
.Y(n_3278)
);

OR2x2_ASAP7_75t_L g3279 ( 
.A(n_3061),
.B(n_2854),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_SL g3280 ( 
.A(n_3104),
.B(n_2855),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_SL g3281 ( 
.A(n_3032),
.B(n_2856),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_3154),
.B(n_2858),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_2992),
.B(n_2887),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_SL g3284 ( 
.A(n_3159),
.B(n_2864),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_SL g3285 ( 
.A(n_3107),
.B(n_2868),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_SL g3286 ( 
.A(n_3115),
.B(n_2869),
.Y(n_3286)
);

NAND2xp33_ASAP7_75t_SL g3287 ( 
.A(n_3131),
.B(n_2350),
.Y(n_3287)
);

NAND2xp33_ASAP7_75t_SL g3288 ( 
.A(n_3132),
.B(n_2350),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_SL g3289 ( 
.A(n_3078),
.B(n_3081),
.Y(n_3289)
);

NAND2xp33_ASAP7_75t_SL g3290 ( 
.A(n_3139),
.B(n_2350),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_SL g3291 ( 
.A(n_3195),
.B(n_2870),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_SL g3292 ( 
.A(n_3090),
.B(n_2871),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3053),
.B(n_2887),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_SL g3294 ( 
.A(n_3090),
.B(n_2872),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_SL g3295 ( 
.A(n_3099),
.B(n_3101),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_SL g3296 ( 
.A(n_3077),
.B(n_2945),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3053),
.B(n_2951),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_SL g3298 ( 
.A(n_3093),
.B(n_2949),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_SL g3299 ( 
.A(n_3147),
.B(n_2876),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_2986),
.B(n_2951),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_SL g3301 ( 
.A(n_3162),
.B(n_2878),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_SL g3302 ( 
.A(n_3166),
.B(n_2880),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_SL g3303 ( 
.A(n_3174),
.B(n_2881),
.Y(n_3303)
);

NAND2xp33_ASAP7_75t_SL g3304 ( 
.A(n_3026),
.B(n_2415),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3088),
.B(n_1187),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3031),
.B(n_2723),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3088),
.B(n_2723),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_SL g3308 ( 
.A(n_3182),
.B(n_3191),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_SL g3309 ( 
.A(n_3111),
.B(n_2873),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3179),
.B(n_2939),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_SL g3311 ( 
.A(n_3111),
.B(n_2882),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_SL g3312 ( 
.A(n_3117),
.B(n_3135),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3179),
.B(n_2940),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_SL g3314 ( 
.A(n_3117),
.B(n_2828),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_SL g3315 ( 
.A(n_3135),
.B(n_2832),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_SL g3316 ( 
.A(n_2997),
.B(n_2894),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_SL g3317 ( 
.A(n_2997),
.B(n_2896),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3142),
.B(n_2943),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_SL g3319 ( 
.A(n_3045),
.B(n_2903),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_SL g3320 ( 
.A(n_3045),
.B(n_2904),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_SL g3321 ( 
.A(n_3070),
.B(n_2907),
.Y(n_3321)
);

NAND2xp33_ASAP7_75t_SL g3322 ( 
.A(n_3178),
.B(n_2415),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_SL g3323 ( 
.A(n_3070),
.B(n_2909),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_3086),
.B(n_2912),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_SL g3325 ( 
.A(n_3086),
.B(n_2927),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_SL g3326 ( 
.A(n_3155),
.B(n_2929),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_SL g3327 ( 
.A(n_2972),
.B(n_3165),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_SL g3328 ( 
.A(n_2975),
.B(n_2824),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_SL g3329 ( 
.A(n_2980),
.B(n_2956),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_SL g3330 ( 
.A(n_2981),
.B(n_3175),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_SL g3331 ( 
.A(n_2994),
.B(n_2957),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3142),
.B(n_2665),
.Y(n_3332)
);

NAND2xp33_ASAP7_75t_SL g3333 ( 
.A(n_2983),
.B(n_2415),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3143),
.B(n_2967),
.Y(n_3334)
);

AND2x4_ASAP7_75t_L g3335 ( 
.A(n_2983),
.B(n_2843),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_SL g3336 ( 
.A(n_2996),
.B(n_2835),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_SL g3337 ( 
.A(n_3000),
.B(n_2775),
.Y(n_3337)
);

NAND2xp33_ASAP7_75t_SL g3338 ( 
.A(n_3027),
.B(n_2415),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_SL g3339 ( 
.A(n_3012),
.B(n_2519),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_SL g3340 ( 
.A(n_3015),
.B(n_2519),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_SL g3341 ( 
.A(n_3025),
.B(n_2519),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_SL g3342 ( 
.A(n_3038),
.B(n_2519),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_3042),
.B(n_3188),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_SL g3344 ( 
.A(n_3051),
.B(n_2565),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_SL g3345 ( 
.A(n_3052),
.B(n_2565),
.Y(n_3345)
);

NAND2xp33_ASAP7_75t_SL g3346 ( 
.A(n_3027),
.B(n_2450),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_SL g3347 ( 
.A(n_3058),
.B(n_2565),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_SL g3348 ( 
.A(n_3064),
.B(n_2565),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_SL g3349 ( 
.A(n_3066),
.B(n_2577),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_SL g3350 ( 
.A(n_3158),
.B(n_2577),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_SL g3351 ( 
.A(n_3161),
.B(n_2577),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_SL g3352 ( 
.A(n_3176),
.B(n_2577),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3152),
.B(n_2866),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_SL g3354 ( 
.A(n_3189),
.B(n_3193),
.Y(n_3354)
);

NAND2xp33_ASAP7_75t_SL g3355 ( 
.A(n_3130),
.B(n_2450),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3160),
.B(n_2440),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_SL g3357 ( 
.A(n_3130),
.B(n_2590),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_SL g3358 ( 
.A(n_3138),
.B(n_2590),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_SL g3359 ( 
.A(n_3138),
.B(n_2590),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_SL g3360 ( 
.A(n_3073),
.B(n_2590),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_SL g3361 ( 
.A(n_3073),
.B(n_2593),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3057),
.B(n_2453),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_SL g3363 ( 
.A(n_2978),
.B(n_3067),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_SL g3364 ( 
.A(n_2978),
.B(n_2593),
.Y(n_3364)
);

NAND2xp33_ASAP7_75t_SL g3365 ( 
.A(n_3041),
.B(n_3060),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_2982),
.B(n_2453),
.Y(n_3366)
);

NAND2xp33_ASAP7_75t_SL g3367 ( 
.A(n_3041),
.B(n_2450),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_3067),
.B(n_2593),
.Y(n_3368)
);

NAND2xp33_ASAP7_75t_SL g3369 ( 
.A(n_3041),
.B(n_2450),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_SL g3370 ( 
.A(n_3039),
.B(n_2593),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_SL g3371 ( 
.A(n_3039),
.B(n_2639),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_SL g3372 ( 
.A(n_3048),
.B(n_3127),
.Y(n_3372)
);

NAND2xp33_ASAP7_75t_SL g3373 ( 
.A(n_3060),
.B(n_2459),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_SL g3374 ( 
.A(n_3137),
.B(n_2639),
.Y(n_3374)
);

AND2x4_ASAP7_75t_L g3375 ( 
.A(n_3173),
.B(n_2319),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_SL g3376 ( 
.A(n_3151),
.B(n_2639),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_SL g3377 ( 
.A(n_3151),
.B(n_2639),
.Y(n_3377)
);

NAND2xp33_ASAP7_75t_SL g3378 ( 
.A(n_3060),
.B(n_2459),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_SL g3379 ( 
.A(n_2998),
.B(n_2652),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_SL g3380 ( 
.A(n_2998),
.B(n_2652),
.Y(n_3380)
);

AND2x2_ASAP7_75t_L g3381 ( 
.A(n_3145),
.B(n_1188),
.Y(n_3381)
);

NAND2xp33_ASAP7_75t_SL g3382 ( 
.A(n_3076),
.B(n_2459),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_SL g3383 ( 
.A(n_3122),
.B(n_2652),
.Y(n_3383)
);

NAND2xp33_ASAP7_75t_SL g3384 ( 
.A(n_3076),
.B(n_2459),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_SL g3385 ( 
.A(n_3122),
.B(n_2652),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_SL g3386 ( 
.A(n_3122),
.B(n_2653),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_2999),
.B(n_2454),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_SL g3388 ( 
.A(n_3128),
.B(n_2653),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3002),
.B(n_2454),
.Y(n_3389)
);

AND2x4_ASAP7_75t_L g3390 ( 
.A(n_3145),
.B(n_2319),
.Y(n_3390)
);

NAND2xp33_ASAP7_75t_SL g3391 ( 
.A(n_3076),
.B(n_2479),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_SL g3392 ( 
.A(n_3128),
.B(n_2653),
.Y(n_3392)
);

AND2x2_ASAP7_75t_L g3393 ( 
.A(n_3145),
.B(n_3023),
.Y(n_3393)
);

NAND2xp33_ASAP7_75t_SL g3394 ( 
.A(n_3085),
.B(n_2479),
.Y(n_3394)
);

AND2x4_ASAP7_75t_L g3395 ( 
.A(n_3046),
.B(n_3187),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_SL g3396 ( 
.A(n_3128),
.B(n_2653),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_SL g3397 ( 
.A(n_3171),
.B(n_2837),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_SL g3398 ( 
.A(n_3108),
.B(n_2837),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3037),
.B(n_2461),
.Y(n_3399)
);

NAND2xp33_ASAP7_75t_SL g3400 ( 
.A(n_3085),
.B(n_2479),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3043),
.B(n_2461),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_SL g3402 ( 
.A(n_3108),
.B(n_2948),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_3268),
.A2(n_3029),
.B(n_3008),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3327),
.Y(n_3404)
);

A2O1A1Ixp33_ASAP7_75t_L g3405 ( 
.A1(n_3216),
.A2(n_3123),
.B(n_3016),
.C(n_3156),
.Y(n_3405)
);

INVx3_ASAP7_75t_L g3406 ( 
.A(n_3395),
.Y(n_3406)
);

AOI21xp5_ASAP7_75t_L g3407 ( 
.A1(n_3270),
.A2(n_3197),
.B(n_3047),
.Y(n_3407)
);

OR2x6_ASAP7_75t_L g3408 ( 
.A(n_3249),
.B(n_3007),
.Y(n_3408)
);

AOI22xp33_ASAP7_75t_SL g3409 ( 
.A1(n_3283),
.A2(n_3011),
.B1(n_2976),
.B2(n_2985),
.Y(n_3409)
);

A2O1A1Ixp33_ASAP7_75t_L g3410 ( 
.A1(n_3207),
.A2(n_3208),
.B(n_3231),
.C(n_3197),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3330),
.Y(n_3411)
);

INVx1_ASAP7_75t_SL g3412 ( 
.A(n_3210),
.Y(n_3412)
);

INVx2_ASAP7_75t_SL g3413 ( 
.A(n_3305),
.Y(n_3413)
);

INVx3_ASAP7_75t_L g3414 ( 
.A(n_3395),
.Y(n_3414)
);

BUFx6f_ASAP7_75t_L g3415 ( 
.A(n_3395),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_L g3416 ( 
.A(n_3272),
.B(n_3022),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3200),
.B(n_3204),
.Y(n_3417)
);

BUFx12f_ASAP7_75t_L g3418 ( 
.A(n_3381),
.Y(n_3418)
);

AOI22xp33_ASAP7_75t_L g3419 ( 
.A1(n_3232),
.A2(n_3112),
.B1(n_3168),
.B2(n_3185),
.Y(n_3419)
);

AOI22xp33_ASAP7_75t_SL g3420 ( 
.A1(n_3203),
.A2(n_3011),
.B1(n_2976),
.B2(n_3082),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3196),
.B(n_3140),
.Y(n_3421)
);

OAI21x1_ASAP7_75t_L g3422 ( 
.A1(n_3372),
.A2(n_3164),
.B(n_2684),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3343),
.Y(n_3423)
);

AND2x4_ASAP7_75t_L g3424 ( 
.A(n_3393),
.B(n_3046),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3354),
.Y(n_3425)
);

INVx3_ASAP7_75t_L g3426 ( 
.A(n_3390),
.Y(n_3426)
);

AND2x4_ASAP7_75t_L g3427 ( 
.A(n_3390),
.B(n_3248),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_3308),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3336),
.Y(n_3429)
);

O2A1O1Ixp33_ASAP7_75t_L g3430 ( 
.A1(n_3234),
.A2(n_778),
.B(n_779),
.C(n_775),
.Y(n_3430)
);

CKINVDCx6p67_ASAP7_75t_R g3431 ( 
.A(n_3244),
.Y(n_3431)
);

AOI22xp33_ASAP7_75t_L g3432 ( 
.A1(n_3196),
.A2(n_3063),
.B1(n_859),
.B2(n_3098),
.Y(n_3432)
);

BUFx6f_ASAP7_75t_L g3433 ( 
.A(n_3247),
.Y(n_3433)
);

A2O1A1Ixp33_ASAP7_75t_SL g3434 ( 
.A1(n_3362),
.A2(n_3136),
.B(n_2884),
.C(n_3113),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_SL g3435 ( 
.A(n_3252),
.B(n_3141),
.Y(n_3435)
);

O2A1O1Ixp33_ASAP7_75t_L g3436 ( 
.A1(n_3209),
.A2(n_782),
.B(n_783),
.C(n_779),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3280),
.B(n_3084),
.Y(n_3437)
);

INVx1_ASAP7_75t_SL g3438 ( 
.A(n_3198),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3279),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3257),
.Y(n_3440)
);

BUFx6f_ASAP7_75t_L g3441 ( 
.A(n_3289),
.Y(n_3441)
);

BUFx6f_ASAP7_75t_L g3442 ( 
.A(n_3375),
.Y(n_3442)
);

NOR2x1_ASAP7_75t_L g3443 ( 
.A(n_3233),
.B(n_3265),
.Y(n_3443)
);

O2A1O1Ixp33_ASAP7_75t_L g3444 ( 
.A1(n_3218),
.A2(n_783),
.B(n_785),
.C(n_782),
.Y(n_3444)
);

AND2x4_ASAP7_75t_L g3445 ( 
.A(n_3390),
.B(n_3096),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3306),
.B(n_3094),
.Y(n_3446)
);

CKINVDCx20_ASAP7_75t_R g3447 ( 
.A(n_3201),
.Y(n_3447)
);

OAI22xp5_ASAP7_75t_L g3448 ( 
.A1(n_3206),
.A2(n_3033),
.B1(n_3156),
.B2(n_3022),
.Y(n_3448)
);

O2A1O1Ixp33_ASAP7_75t_L g3449 ( 
.A1(n_3239),
.A2(n_788),
.B(n_792),
.C(n_785),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3227),
.B(n_3103),
.Y(n_3450)
);

INVx2_ASAP7_75t_SL g3451 ( 
.A(n_3368),
.Y(n_3451)
);

BUFx6f_ASAP7_75t_L g3452 ( 
.A(n_3375),
.Y(n_3452)
);

OAI22xp5_ASAP7_75t_SL g3453 ( 
.A1(n_3297),
.A2(n_3056),
.B1(n_792),
.B2(n_793),
.Y(n_3453)
);

AOI22xp33_ASAP7_75t_SL g3454 ( 
.A1(n_3274),
.A2(n_3004),
.B1(n_3007),
.B2(n_3098),
.Y(n_3454)
);

BUFx2_ASAP7_75t_L g3455 ( 
.A(n_3230),
.Y(n_3455)
);

HB1xp67_ASAP7_75t_L g3456 ( 
.A(n_3243),
.Y(n_3456)
);

AOI21xp5_ASAP7_75t_L g3457 ( 
.A1(n_3398),
.A2(n_3226),
.B(n_3261),
.Y(n_3457)
);

AOI21xp5_ASAP7_75t_L g3458 ( 
.A1(n_3398),
.A2(n_3361),
.B(n_3360),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_R g3459 ( 
.A(n_3266),
.B(n_3007),
.Y(n_3459)
);

A2O1A1Ixp33_ASAP7_75t_L g3460 ( 
.A1(n_3224),
.A2(n_2682),
.B(n_2703),
.C(n_793),
.Y(n_3460)
);

HB1xp67_ASAP7_75t_L g3461 ( 
.A(n_3307),
.Y(n_3461)
);

HAxp5_ASAP7_75t_L g3462 ( 
.A(n_3205),
.B(n_720),
.CON(n_3462),
.SN(n_3462)
);

NOR2xp33_ASAP7_75t_L g3463 ( 
.A(n_3222),
.B(n_3035),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3219),
.B(n_3105),
.Y(n_3464)
);

BUFx2_ASAP7_75t_L g3465 ( 
.A(n_3365),
.Y(n_3465)
);

AOI222xp33_ASAP7_75t_L g3466 ( 
.A1(n_3223),
.A2(n_788),
.B1(n_818),
.B2(n_837),
.C1(n_835),
.C2(n_803),
.Y(n_3466)
);

BUFx2_ASAP7_75t_L g3467 ( 
.A(n_3212),
.Y(n_3467)
);

BUFx3_ASAP7_75t_L g3468 ( 
.A(n_3375),
.Y(n_3468)
);

A2O1A1Ixp33_ASAP7_75t_L g3469 ( 
.A1(n_3225),
.A2(n_3263),
.B(n_3260),
.C(n_3228),
.Y(n_3469)
);

BUFx2_ASAP7_75t_L g3470 ( 
.A(n_3275),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3221),
.B(n_3110),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3366),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3245),
.Y(n_3473)
);

OAI22xp5_ASAP7_75t_L g3474 ( 
.A1(n_3214),
.A2(n_2745),
.B1(n_2984),
.B2(n_3083),
.Y(n_3474)
);

BUFx6f_ASAP7_75t_L g3475 ( 
.A(n_3220),
.Y(n_3475)
);

INVx3_ASAP7_75t_L g3476 ( 
.A(n_3220),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3246),
.Y(n_3477)
);

INVx5_ASAP7_75t_L g3478 ( 
.A(n_3248),
.Y(n_3478)
);

INVxp67_ASAP7_75t_L g3479 ( 
.A(n_3242),
.Y(n_3479)
);

O2A1O1Ixp5_ASAP7_75t_L g3480 ( 
.A1(n_3402),
.A2(n_3397),
.B(n_3276),
.C(n_3273),
.Y(n_3480)
);

AND2x2_ASAP7_75t_SL g3481 ( 
.A(n_3235),
.B(n_3065),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3387),
.Y(n_3482)
);

AOI22xp5_ASAP7_75t_L g3483 ( 
.A1(n_3211),
.A2(n_3098),
.B1(n_733),
.B2(n_737),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3202),
.B(n_3120),
.Y(n_3484)
);

BUFx3_ASAP7_75t_L g3485 ( 
.A(n_3248),
.Y(n_3485)
);

INVx1_ASAP7_75t_SL g3486 ( 
.A(n_3312),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_3389),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3379),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_R g3489 ( 
.A(n_3267),
.B(n_3287),
.Y(n_3489)
);

INVx1_ASAP7_75t_SL g3490 ( 
.A(n_3293),
.Y(n_3490)
);

CKINVDCx16_ASAP7_75t_R g3491 ( 
.A(n_3288),
.Y(n_3491)
);

AOI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3397),
.A2(n_3286),
.B(n_3285),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3399),
.Y(n_3493)
);

OAI22xp5_ASAP7_75t_SL g3494 ( 
.A1(n_3300),
.A2(n_3229),
.B1(n_3269),
.B2(n_3262),
.Y(n_3494)
);

BUFx3_ASAP7_75t_L g3495 ( 
.A(n_3335),
.Y(n_3495)
);

AOI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_3402),
.A2(n_2831),
.B(n_2734),
.Y(n_3496)
);

INVx4_ASAP7_75t_L g3497 ( 
.A(n_3335),
.Y(n_3497)
);

OAI221xp5_ASAP7_75t_L g3498 ( 
.A1(n_3213),
.A2(n_1177),
.B1(n_818),
.B2(n_835),
.C(n_804),
.Y(n_3498)
);

AOI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_3202),
.A2(n_3371),
.B(n_3370),
.Y(n_3499)
);

INVx2_ASAP7_75t_SL g3500 ( 
.A(n_3309),
.Y(n_3500)
);

NOR2xp33_ASAP7_75t_L g3501 ( 
.A(n_3363),
.B(n_3125),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3295),
.B(n_3126),
.Y(n_3502)
);

CKINVDCx5p33_ASAP7_75t_R g3503 ( 
.A(n_3241),
.Y(n_3503)
);

INVx3_ASAP7_75t_L g3504 ( 
.A(n_3335),
.Y(n_3504)
);

NOR2x1_ASAP7_75t_L g3505 ( 
.A(n_3282),
.B(n_3169),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3401),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3334),
.B(n_3044),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3380),
.Y(n_3508)
);

INVx6_ASAP7_75t_L g3509 ( 
.A(n_3238),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_3299),
.Y(n_3510)
);

NOR2xp67_ASAP7_75t_L g3511 ( 
.A(n_3296),
.B(n_3049),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_3301),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3357),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3217),
.B(n_3291),
.Y(n_3514)
);

OAI21x1_ASAP7_75t_SL g3515 ( 
.A1(n_3353),
.A2(n_3190),
.B(n_3164),
.Y(n_3515)
);

NOR2xp67_ASAP7_75t_SL g3516 ( 
.A(n_3251),
.B(n_3146),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_SL g3517 ( 
.A(n_3215),
.B(n_3146),
.Y(n_3517)
);

NOR2xp33_ASAP7_75t_L g3518 ( 
.A(n_3240),
.B(n_3062),
.Y(n_3518)
);

BUFx6f_ASAP7_75t_L g3519 ( 
.A(n_3238),
.Y(n_3519)
);

AOI21xp5_ASAP7_75t_L g3520 ( 
.A1(n_3199),
.A2(n_2434),
.B(n_2359),
.Y(n_3520)
);

INVx3_ASAP7_75t_L g3521 ( 
.A(n_3238),
.Y(n_3521)
);

BUFx6f_ASAP7_75t_L g3522 ( 
.A(n_3258),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_SL g3523 ( 
.A(n_3250),
.B(n_3146),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3302),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_3303),
.Y(n_3525)
);

INVx2_ASAP7_75t_SL g3526 ( 
.A(n_3311),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3358),
.Y(n_3527)
);

AOI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_3199),
.A2(n_2434),
.B(n_2359),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3359),
.Y(n_3529)
);

CKINVDCx16_ASAP7_75t_R g3530 ( 
.A(n_3290),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3364),
.Y(n_3531)
);

INVx4_ASAP7_75t_L g3532 ( 
.A(n_3264),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3328),
.Y(n_3533)
);

OAI22xp5_ASAP7_75t_L g3534 ( 
.A1(n_3277),
.A2(n_2745),
.B1(n_3083),
.B2(n_2984),
.Y(n_3534)
);

BUFx6f_ASAP7_75t_L g3535 ( 
.A(n_3383),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3329),
.Y(n_3536)
);

OAI22xp5_ASAP7_75t_L g3537 ( 
.A1(n_3278),
.A2(n_3114),
.B1(n_3071),
.B2(n_3075),
.Y(n_3537)
);

AOI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_3236),
.A2(n_3098),
.B1(n_738),
.B2(n_739),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_SL g3539 ( 
.A(n_3253),
.B(n_3069),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3331),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3339),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_SL g3542 ( 
.A(n_3281),
.B(n_3080),
.Y(n_3542)
);

BUFx6f_ASAP7_75t_L g3543 ( 
.A(n_3385),
.Y(n_3543)
);

O2A1O1Ixp33_ASAP7_75t_L g3544 ( 
.A1(n_3254),
.A2(n_804),
.B(n_837),
.C(n_803),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3340),
.Y(n_3545)
);

OAI21xp5_ASAP7_75t_L g3546 ( 
.A1(n_3259),
.A2(n_3326),
.B(n_3256),
.Y(n_3546)
);

CKINVDCx16_ASAP7_75t_R g3547 ( 
.A(n_3322),
.Y(n_3547)
);

AO22x1_ASAP7_75t_L g3548 ( 
.A1(n_3318),
.A2(n_842),
.B1(n_848),
.B2(n_841),
.Y(n_3548)
);

AOI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_3310),
.A2(n_2434),
.B(n_2359),
.Y(n_3549)
);

BUFx6f_ASAP7_75t_L g3550 ( 
.A(n_3386),
.Y(n_3550)
);

AOI22xp33_ASAP7_75t_L g3551 ( 
.A1(n_3237),
.A2(n_2422),
.B1(n_2497),
.B2(n_2430),
.Y(n_3551)
);

INVx2_ASAP7_75t_SL g3552 ( 
.A(n_3388),
.Y(n_3552)
);

AOI22xp5_ASAP7_75t_L g3553 ( 
.A1(n_3255),
.A2(n_740),
.B1(n_742),
.B2(n_729),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_SL g3554 ( 
.A(n_3271),
.B(n_3095),
.Y(n_3554)
);

OR2x2_ASAP7_75t_L g3555 ( 
.A(n_3313),
.B(n_3096),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3341),
.Y(n_3556)
);

NOR2xp33_ASAP7_75t_L g3557 ( 
.A(n_3298),
.B(n_3113),
.Y(n_3557)
);

BUFx4f_ASAP7_75t_L g3558 ( 
.A(n_3304),
.Y(n_3558)
);

AND2x4_ASAP7_75t_L g3559 ( 
.A(n_3314),
.B(n_3124),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3342),
.Y(n_3560)
);

INVx5_ASAP7_75t_L g3561 ( 
.A(n_3367),
.Y(n_3561)
);

OAI22xp5_ASAP7_75t_L g3562 ( 
.A1(n_3292),
.A2(n_3114),
.B1(n_2944),
.B2(n_2494),
.Y(n_3562)
);

OAI22xp5_ASAP7_75t_L g3563 ( 
.A1(n_3294),
.A2(n_3284),
.B1(n_3315),
.B2(n_3376),
.Y(n_3563)
);

AND2x4_ASAP7_75t_L g3564 ( 
.A(n_3344),
.B(n_3124),
.Y(n_3564)
);

NOR2xp33_ASAP7_75t_L g3565 ( 
.A(n_3319),
.B(n_3170),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_3374),
.Y(n_3566)
);

INVx1_ASAP7_75t_SL g3567 ( 
.A(n_3392),
.Y(n_3567)
);

INVx5_ASAP7_75t_L g3568 ( 
.A(n_3369),
.Y(n_3568)
);

NOR2xp33_ASAP7_75t_L g3569 ( 
.A(n_3320),
.B(n_3170),
.Y(n_3569)
);

OAI22xp5_ASAP7_75t_L g3570 ( 
.A1(n_3377),
.A2(n_2944),
.B1(n_3194),
.B2(n_3187),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_3345),
.Y(n_3571)
);

BUFx3_ASAP7_75t_L g3572 ( 
.A(n_3332),
.Y(n_3572)
);

INVx1_ASAP7_75t_SL g3573 ( 
.A(n_3396),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3356),
.B(n_3194),
.Y(n_3574)
);

OR2x4_ASAP7_75t_L g3575 ( 
.A(n_3333),
.B(n_3085),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3321),
.B(n_3087),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3347),
.Y(n_3577)
);

BUFx6f_ASAP7_75t_L g3578 ( 
.A(n_3348),
.Y(n_3578)
);

INVx4_ASAP7_75t_L g3579 ( 
.A(n_3338),
.Y(n_3579)
);

AOI22xp5_ASAP7_75t_L g3580 ( 
.A1(n_3355),
.A2(n_747),
.B1(n_748),
.B2(n_745),
.Y(n_3580)
);

INVx2_ASAP7_75t_L g3581 ( 
.A(n_3349),
.Y(n_3581)
);

NOR2xp33_ASAP7_75t_L g3582 ( 
.A(n_3323),
.B(n_3087),
.Y(n_3582)
);

O2A1O1Ixp33_ASAP7_75t_L g3583 ( 
.A1(n_3316),
.A2(n_3317),
.B(n_3325),
.C(n_3324),
.Y(n_3583)
);

NOR2xp33_ASAP7_75t_L g3584 ( 
.A(n_3350),
.B(n_3087),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_3351),
.Y(n_3585)
);

OR2x2_ASAP7_75t_L g3586 ( 
.A(n_3337),
.B(n_3352),
.Y(n_3586)
);

INVx2_ASAP7_75t_L g3587 ( 
.A(n_3346),
.Y(n_3587)
);

A2O1A1Ixp33_ASAP7_75t_L g3588 ( 
.A1(n_3373),
.A2(n_842),
.B(n_848),
.C(n_841),
.Y(n_3588)
);

INVx4_ASAP7_75t_L g3589 ( 
.A(n_3378),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3382),
.Y(n_3590)
);

INVx5_ASAP7_75t_L g3591 ( 
.A(n_3384),
.Y(n_3591)
);

OR2x2_ASAP7_75t_L g3592 ( 
.A(n_3391),
.B(n_3097),
.Y(n_3592)
);

BUFx6f_ASAP7_75t_L g3593 ( 
.A(n_3394),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3400),
.Y(n_3594)
);

CKINVDCx6p67_ASAP7_75t_R g3595 ( 
.A(n_3244),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3200),
.B(n_3097),
.Y(n_3596)
);

OAI21xp33_ASAP7_75t_SL g3597 ( 
.A1(n_3197),
.A2(n_3169),
.B(n_3065),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3308),
.Y(n_3598)
);

INVx4_ASAP7_75t_L g3599 ( 
.A(n_3375),
.Y(n_3599)
);

BUFx3_ASAP7_75t_L g3600 ( 
.A(n_3247),
.Y(n_3600)
);

HB1xp67_ASAP7_75t_L g3601 ( 
.A(n_3257),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_3308),
.Y(n_3602)
);

OR2x6_ASAP7_75t_L g3603 ( 
.A(n_3249),
.B(n_3097),
.Y(n_3603)
);

BUFx2_ASAP7_75t_L g3604 ( 
.A(n_3393),
.Y(n_3604)
);

CKINVDCx5p33_ASAP7_75t_R g3605 ( 
.A(n_3201),
.Y(n_3605)
);

BUFx6f_ASAP7_75t_L g3606 ( 
.A(n_3395),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3200),
.B(n_3144),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3200),
.B(n_3144),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3268),
.A2(n_2434),
.B(n_2518),
.Y(n_3609)
);

INVx4_ASAP7_75t_L g3610 ( 
.A(n_3375),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3327),
.Y(n_3611)
);

AND2x4_ASAP7_75t_L g3612 ( 
.A(n_3393),
.B(n_3144),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3327),
.Y(n_3613)
);

AOI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_3268),
.A2(n_2518),
.B(n_2159),
.Y(n_3614)
);

AOI22xp5_ASAP7_75t_L g3615 ( 
.A1(n_3410),
.A2(n_753),
.B1(n_756),
.B2(n_752),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_3461),
.B(n_757),
.Y(n_3616)
);

NAND3xp33_ASAP7_75t_L g3617 ( 
.A(n_3469),
.B(n_857),
.C(n_855),
.Y(n_3617)
);

OAI21x1_ASAP7_75t_L g3618 ( 
.A1(n_3496),
.A2(n_2766),
.B(n_2335),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3417),
.B(n_760),
.Y(n_3619)
);

NOR2xp33_ASAP7_75t_L g3620 ( 
.A(n_3431),
.B(n_762),
.Y(n_3620)
);

AO31x2_ASAP7_75t_L g3621 ( 
.A1(n_3457),
.A2(n_2335),
.A3(n_2344),
.B(n_2328),
.Y(n_3621)
);

A2O1A1Ixp33_ASAP7_75t_L g3622 ( 
.A1(n_3480),
.A2(n_857),
.B(n_865),
.C(n_855),
.Y(n_3622)
);

AOI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_3403),
.A2(n_2344),
.B(n_2328),
.Y(n_3623)
);

NOR2xp33_ASAP7_75t_L g3624 ( 
.A(n_3595),
.B(n_764),
.Y(n_3624)
);

AND2x2_ASAP7_75t_L g3625 ( 
.A(n_3604),
.B(n_865),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3404),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3439),
.B(n_767),
.Y(n_3627)
);

A2O1A1Ixp33_ASAP7_75t_L g3628 ( 
.A1(n_3405),
.A2(n_870),
.B(n_876),
.C(n_866),
.Y(n_3628)
);

NAND3xp33_ASAP7_75t_L g3629 ( 
.A(n_3466),
.B(n_870),
.C(n_866),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3411),
.Y(n_3630)
);

AOI21x1_ASAP7_75t_L g3631 ( 
.A1(n_3548),
.A2(n_1306),
.B(n_1305),
.Y(n_3631)
);

NOR2xp67_ASAP7_75t_L g3632 ( 
.A(n_3479),
.B(n_1189),
.Y(n_3632)
);

OAI21x1_ASAP7_75t_L g3633 ( 
.A1(n_3422),
.A2(n_2351),
.B(n_2464),
.Y(n_3633)
);

A2O1A1Ixp33_ASAP7_75t_L g3634 ( 
.A1(n_3546),
.A2(n_879),
.B(n_880),
.C(n_876),
.Y(n_3634)
);

INVx2_ASAP7_75t_SL g3635 ( 
.A(n_3413),
.Y(n_3635)
);

AOI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_3407),
.A2(n_2351),
.B(n_2329),
.Y(n_3636)
);

O2A1O1Ixp33_ASAP7_75t_SL g3637 ( 
.A1(n_3523),
.A2(n_880),
.B(n_887),
.C(n_879),
.Y(n_3637)
);

AOI21xp5_ASAP7_75t_L g3638 ( 
.A1(n_3558),
.A2(n_2407),
.B(n_2355),
.Y(n_3638)
);

AOI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3558),
.A2(n_2407),
.B(n_2355),
.Y(n_3639)
);

HB1xp67_ASAP7_75t_L g3640 ( 
.A(n_3601),
.Y(n_3640)
);

O2A1O1Ixp5_ASAP7_75t_L g3641 ( 
.A1(n_3516),
.A2(n_898),
.B(n_900),
.C(n_887),
.Y(n_3641)
);

AND2x2_ASAP7_75t_L g3642 ( 
.A(n_3433),
.B(n_898),
.Y(n_3642)
);

INVx2_ASAP7_75t_SL g3643 ( 
.A(n_3600),
.Y(n_3643)
);

AO31x2_ASAP7_75t_L g3644 ( 
.A1(n_3609),
.A2(n_2468),
.A3(n_2476),
.B(n_2452),
.Y(n_3644)
);

AO32x2_ASAP7_75t_L g3645 ( 
.A1(n_3494),
.A2(n_3563),
.A3(n_3500),
.B1(n_3526),
.B2(n_3497),
.Y(n_3645)
);

A2O1A1Ixp33_ASAP7_75t_L g3646 ( 
.A1(n_3458),
.A2(n_901),
.B(n_908),
.C(n_900),
.Y(n_3646)
);

AO31x2_ASAP7_75t_L g3647 ( 
.A1(n_3520),
.A2(n_2468),
.A3(n_2476),
.B(n_2452),
.Y(n_3647)
);

AOI21xp5_ASAP7_75t_L g3648 ( 
.A1(n_3492),
.A2(n_2515),
.B(n_2509),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3423),
.Y(n_3649)
);

AOI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_3614),
.A2(n_2515),
.B(n_2509),
.Y(n_3650)
);

AOI22xp5_ASAP7_75t_L g3651 ( 
.A1(n_3443),
.A2(n_774),
.B1(n_781),
.B2(n_769),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3490),
.B(n_3572),
.Y(n_3652)
);

AOI221x1_ASAP7_75t_L g3653 ( 
.A1(n_3473),
.A2(n_915),
.B1(n_917),
.B2(n_908),
.C(n_901),
.Y(n_3653)
);

OAI22xp5_ASAP7_75t_L g3654 ( 
.A1(n_3420),
.A2(n_917),
.B1(n_931),
.B2(n_915),
.Y(n_3654)
);

INVx1_ASAP7_75t_SL g3655 ( 
.A(n_3438),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3425),
.Y(n_3656)
);

AO31x2_ASAP7_75t_L g3657 ( 
.A1(n_3528),
.A2(n_2527),
.A3(n_2548),
.B(n_2523),
.Y(n_3657)
);

OAI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_3432),
.A2(n_936),
.B(n_931),
.Y(n_3658)
);

OAI21x1_ASAP7_75t_L g3659 ( 
.A1(n_3549),
.A2(n_2469),
.B(n_2466),
.Y(n_3659)
);

OR2x2_ASAP7_75t_L g3660 ( 
.A(n_3412),
.B(n_1305),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3477),
.B(n_784),
.Y(n_3661)
);

OR2x2_ASAP7_75t_L g3662 ( 
.A(n_3433),
.B(n_1306),
.Y(n_3662)
);

OAI22xp5_ASAP7_75t_L g3663 ( 
.A1(n_3409),
.A2(n_3503),
.B1(n_3419),
.B2(n_3455),
.Y(n_3663)
);

BUFx3_ASAP7_75t_L g3664 ( 
.A(n_3418),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3611),
.Y(n_3665)
);

OAI21x1_ASAP7_75t_SL g3666 ( 
.A1(n_3583),
.A2(n_939),
.B(n_936),
.Y(n_3666)
);

INVx2_ASAP7_75t_SL g3667 ( 
.A(n_3433),
.Y(n_3667)
);

OAI21x1_ASAP7_75t_L g3668 ( 
.A1(n_3515),
.A2(n_2469),
.B(n_2466),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3613),
.Y(n_3669)
);

OAI21x1_ASAP7_75t_L g3670 ( 
.A1(n_3499),
.A2(n_2486),
.B(n_2478),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3456),
.B(n_789),
.Y(n_3671)
);

AO31x2_ASAP7_75t_L g3672 ( 
.A1(n_3429),
.A2(n_2527),
.A3(n_2548),
.B(n_2523),
.Y(n_3672)
);

INVx3_ASAP7_75t_L g3673 ( 
.A(n_3612),
.Y(n_3673)
);

AO31x2_ASAP7_75t_L g3674 ( 
.A1(n_3534),
.A2(n_940),
.A3(n_942),
.B(n_939),
.Y(n_3674)
);

AOI21xp5_ASAP7_75t_L g3675 ( 
.A1(n_3561),
.A2(n_2580),
.B(n_2563),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3428),
.Y(n_3676)
);

AOI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_3561),
.A2(n_2580),
.B(n_2563),
.Y(n_3677)
);

AO31x2_ASAP7_75t_L g3678 ( 
.A1(n_3474),
.A2(n_942),
.A3(n_943),
.B(n_940),
.Y(n_3678)
);

AOI22x1_ASAP7_75t_L g3679 ( 
.A1(n_3467),
.A2(n_794),
.B1(n_797),
.B2(n_790),
.Y(n_3679)
);

OAI21x1_ASAP7_75t_L g3680 ( 
.A1(n_3484),
.A2(n_2486),
.B(n_2478),
.Y(n_3680)
);

BUFx2_ASAP7_75t_L g3681 ( 
.A(n_3441),
.Y(n_3681)
);

AO31x2_ASAP7_75t_L g3682 ( 
.A1(n_3589),
.A2(n_943),
.A3(n_2621),
.B(n_2596),
.Y(n_3682)
);

INVx1_ASAP7_75t_SL g3683 ( 
.A(n_3463),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_SL g3684 ( 
.A(n_3481),
.B(n_3150),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3416),
.B(n_806),
.Y(n_3685)
);

O2A1O1Ixp33_ASAP7_75t_L g3686 ( 
.A1(n_3462),
.A2(n_1191),
.B(n_1192),
.C(n_1190),
.Y(n_3686)
);

A2O1A1Ixp33_ASAP7_75t_L g3687 ( 
.A1(n_3430),
.A2(n_812),
.B(n_813),
.C(n_808),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3514),
.B(n_814),
.Y(n_3688)
);

OAI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_3460),
.A2(n_1198),
.B(n_1194),
.Y(n_3689)
);

OAI21x1_ASAP7_75t_L g3690 ( 
.A1(n_3554),
.A2(n_2582),
.B(n_2570),
.Y(n_3690)
);

OAI21xp5_ASAP7_75t_L g3691 ( 
.A1(n_3483),
.A2(n_1201),
.B(n_1200),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3440),
.B(n_819),
.Y(n_3692)
);

AOI21xp5_ASAP7_75t_L g3693 ( 
.A1(n_3561),
.A2(n_2621),
.B(n_2596),
.Y(n_3693)
);

INVxp67_ASAP7_75t_SL g3694 ( 
.A(n_3421),
.Y(n_3694)
);

AOI221xp5_ASAP7_75t_SL g3695 ( 
.A1(n_3453),
.A2(n_1206),
.B1(n_1212),
.B2(n_1204),
.C(n_1202),
.Y(n_3695)
);

AOI22xp5_ASAP7_75t_L g3696 ( 
.A1(n_3448),
.A2(n_822),
.B1(n_825),
.B2(n_821),
.Y(n_3696)
);

AOI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_3568),
.A2(n_2479),
.B(n_2300),
.Y(n_3697)
);

CKINVDCx20_ASAP7_75t_R g3698 ( 
.A(n_3447),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3555),
.B(n_828),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3533),
.B(n_831),
.Y(n_3700)
);

AO32x2_ASAP7_75t_L g3701 ( 
.A1(n_3497),
.A2(n_5),
.A3(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3536),
.B(n_833),
.Y(n_3702)
);

A2O1A1Ixp33_ASAP7_75t_L g3703 ( 
.A1(n_3444),
.A2(n_3436),
.B(n_3449),
.C(n_3538),
.Y(n_3703)
);

INVx4_ASAP7_75t_L g3704 ( 
.A(n_3612),
.Y(n_3704)
);

A2O1A1Ixp33_ASAP7_75t_L g3705 ( 
.A1(n_3501),
.A2(n_3544),
.B(n_3580),
.C(n_3434),
.Y(n_3705)
);

CKINVDCx20_ASAP7_75t_R g3706 ( 
.A(n_3605),
.Y(n_3706)
);

AOI21xp5_ASAP7_75t_L g3707 ( 
.A1(n_3568),
.A2(n_2300),
.B(n_2537),
.Y(n_3707)
);

O2A1O1Ixp33_ASAP7_75t_SL g3708 ( 
.A1(n_3517),
.A2(n_1214),
.B(n_1215),
.C(n_1213),
.Y(n_3708)
);

INVx1_ASAP7_75t_SL g3709 ( 
.A(n_3424),
.Y(n_3709)
);

O2A1O1Ixp33_ASAP7_75t_L g3710 ( 
.A1(n_3588),
.A2(n_1220),
.B(n_1222),
.C(n_1216),
.Y(n_3710)
);

OR2x2_ASAP7_75t_L g3711 ( 
.A(n_3521),
.B(n_1224),
.Y(n_3711)
);

NAND3xp33_ASAP7_75t_L g3712 ( 
.A(n_3548),
.B(n_1230),
.C(n_1227),
.Y(n_3712)
);

AOI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_3568),
.A2(n_2560),
.B(n_2280),
.Y(n_3713)
);

OAI21xp33_ASAP7_75t_L g3714 ( 
.A1(n_3518),
.A2(n_836),
.B(n_834),
.Y(n_3714)
);

BUFx6f_ASAP7_75t_L g3715 ( 
.A(n_3415),
.Y(n_3715)
);

OAI21x1_ASAP7_75t_L g3716 ( 
.A1(n_3570),
.A2(n_2582),
.B(n_2570),
.Y(n_3716)
);

AOI21xp5_ASAP7_75t_L g3717 ( 
.A1(n_3591),
.A2(n_2560),
.B(n_2387),
.Y(n_3717)
);

AO31x2_ASAP7_75t_L g3718 ( 
.A1(n_3488),
.A2(n_2481),
.A3(n_2491),
.B(n_2480),
.Y(n_3718)
);

AOI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_3591),
.A2(n_2388),
.B(n_2380),
.Y(n_3719)
);

AO31x2_ASAP7_75t_L g3720 ( 
.A1(n_3508),
.A2(n_2481),
.A3(n_2491),
.B(n_2480),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3540),
.B(n_3596),
.Y(n_3721)
);

OAI21xp5_ASAP7_75t_L g3722 ( 
.A1(n_3597),
.A2(n_1234),
.B(n_1231),
.Y(n_3722)
);

INVxp67_ASAP7_75t_L g3723 ( 
.A(n_3607),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3513),
.Y(n_3724)
);

OAI21x1_ASAP7_75t_L g3725 ( 
.A1(n_3574),
.A2(n_3537),
.B(n_3529),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3608),
.B(n_839),
.Y(n_3726)
);

AOI21xp5_ASAP7_75t_L g3727 ( 
.A1(n_3591),
.A2(n_2418),
.B(n_2388),
.Y(n_3727)
);

BUFx10_ASAP7_75t_L g3728 ( 
.A(n_3424),
.Y(n_3728)
);

AO31x2_ASAP7_75t_L g3729 ( 
.A1(n_3527),
.A2(n_2505),
.A3(n_2510),
.B(n_2504),
.Y(n_3729)
);

O2A1O1Ixp33_ASAP7_75t_SL g3730 ( 
.A1(n_3435),
.A2(n_1272),
.B(n_1273),
.C(n_1262),
.Y(n_3730)
);

OAI21x1_ASAP7_75t_L g3731 ( 
.A1(n_3531),
.A2(n_2612),
.B(n_2585),
.Y(n_3731)
);

OAI21x1_ASAP7_75t_L g3732 ( 
.A1(n_3571),
.A2(n_2612),
.B(n_2585),
.Y(n_3732)
);

INVxp67_ASAP7_75t_SL g3733 ( 
.A(n_3586),
.Y(n_3733)
);

AOI31xp67_ASAP7_75t_L g3734 ( 
.A1(n_3590),
.A2(n_2505),
.A3(n_2510),
.B(n_2504),
.Y(n_3734)
);

NOR2xp33_ASAP7_75t_L g3735 ( 
.A(n_3441),
.B(n_840),
.Y(n_3735)
);

OAI21xp5_ASAP7_75t_L g3736 ( 
.A1(n_3505),
.A2(n_1277),
.B(n_1276),
.Y(n_3736)
);

CKINVDCx20_ASAP7_75t_R g3737 ( 
.A(n_3485),
.Y(n_3737)
);

AO31x2_ASAP7_75t_L g3738 ( 
.A1(n_3589),
.A2(n_1282),
.A3(n_1284),
.B(n_1279),
.Y(n_3738)
);

CKINVDCx5p33_ASAP7_75t_R g3739 ( 
.A(n_3415),
.Y(n_3739)
);

CKINVDCx20_ASAP7_75t_R g3740 ( 
.A(n_3495),
.Y(n_3740)
);

OAI21x1_ASAP7_75t_L g3741 ( 
.A1(n_3581),
.A2(n_2630),
.B(n_2614),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_3539),
.A2(n_2421),
.B(n_2418),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3450),
.B(n_845),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3521),
.B(n_3150),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3541),
.Y(n_3745)
);

OAI21x1_ASAP7_75t_L g3746 ( 
.A1(n_3585),
.A2(n_2630),
.B(n_2614),
.Y(n_3746)
);

BUFx6f_ASAP7_75t_L g3747 ( 
.A(n_3415),
.Y(n_3747)
);

O2A1O1Ixp33_ASAP7_75t_SL g3748 ( 
.A1(n_3451),
.A2(n_1287),
.B(n_1288),
.C(n_1285),
.Y(n_3748)
);

AOI22xp5_ASAP7_75t_L g3749 ( 
.A1(n_3408),
.A2(n_847),
.B1(n_849),
.B2(n_846),
.Y(n_3749)
);

A2O1A1Ixp33_ASAP7_75t_L g3750 ( 
.A1(n_3470),
.A2(n_853),
.B(n_858),
.C(n_850),
.Y(n_3750)
);

NOR2xp33_ASAP7_75t_L g3751 ( 
.A(n_3441),
.B(n_861),
.Y(n_3751)
);

AOI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_3579),
.A2(n_2421),
.B(n_2283),
.Y(n_3752)
);

CKINVDCx11_ASAP7_75t_R g3753 ( 
.A(n_3606),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3545),
.Y(n_3754)
);

CKINVDCx5p33_ASAP7_75t_R g3755 ( 
.A(n_3606),
.Y(n_3755)
);

AND2x4_ASAP7_75t_L g3756 ( 
.A(n_3406),
.B(n_3150),
.Y(n_3756)
);

INVx3_ASAP7_75t_L g3757 ( 
.A(n_3606),
.Y(n_3757)
);

NAND3xp33_ASAP7_75t_L g3758 ( 
.A(n_3565),
.B(n_1316),
.C(n_1315),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3556),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3560),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3577),
.Y(n_3761)
);

O2A1O1Ixp5_ASAP7_75t_L g3762 ( 
.A1(n_3532),
.A2(n_1319),
.B(n_1238),
.C(n_1239),
.Y(n_3762)
);

OAI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_3542),
.A2(n_2497),
.B(n_2430),
.Y(n_3763)
);

OA21x2_ASAP7_75t_L g3764 ( 
.A1(n_3594),
.A2(n_1238),
.B(n_1237),
.Y(n_3764)
);

BUFx3_ASAP7_75t_L g3765 ( 
.A(n_3445),
.Y(n_3765)
);

AOI22xp5_ASAP7_75t_L g3766 ( 
.A1(n_3408),
.A2(n_871),
.B1(n_873),
.B2(n_863),
.Y(n_3766)
);

OAI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_3553),
.A2(n_2497),
.B(n_2430),
.Y(n_3767)
);

OAI22x1_ASAP7_75t_L g3768 ( 
.A1(n_3478),
.A2(n_878),
.B1(n_881),
.B2(n_874),
.Y(n_3768)
);

O2A1O1Ixp33_ASAP7_75t_L g3769 ( 
.A1(n_3498),
.A2(n_1239),
.B(n_1240),
.C(n_1237),
.Y(n_3769)
);

AOI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3579),
.A2(n_2294),
.B(n_2277),
.Y(n_3770)
);

AOI21xp5_ASAP7_75t_L g3771 ( 
.A1(n_3532),
.A2(n_2637),
.B(n_2632),
.Y(n_3771)
);

AOI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3478),
.A2(n_2637),
.B(n_2632),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3504),
.B(n_1240),
.Y(n_3773)
);

BUFx6f_ASAP7_75t_L g3774 ( 
.A(n_3442),
.Y(n_3774)
);

AO31x2_ASAP7_75t_L g3775 ( 
.A1(n_3569),
.A2(n_2530),
.A3(n_2544),
.B(n_2521),
.Y(n_3775)
);

OAI21x1_ASAP7_75t_L g3776 ( 
.A1(n_3566),
.A2(n_2530),
.B(n_2521),
.Y(n_3776)
);

INVx2_ASAP7_75t_L g3777 ( 
.A(n_3598),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3478),
.A2(n_2545),
.B(n_2544),
.Y(n_3778)
);

NOR2xp33_ASAP7_75t_L g3779 ( 
.A(n_3522),
.B(n_884),
.Y(n_3779)
);

AO31x2_ASAP7_75t_L g3780 ( 
.A1(n_3582),
.A2(n_3562),
.A3(n_3584),
.B(n_3602),
.Y(n_3780)
);

AOI21xp5_ASAP7_75t_L g3781 ( 
.A1(n_3507),
.A2(n_2561),
.B(n_2545),
.Y(n_3781)
);

OAI22xp5_ASAP7_75t_L g3782 ( 
.A1(n_3491),
.A2(n_888),
.B1(n_889),
.B2(n_885),
.Y(n_3782)
);

OAI21xp5_ASAP7_75t_L g3783 ( 
.A1(n_3437),
.A2(n_2497),
.B(n_1242),
.Y(n_3783)
);

OAI21x1_ASAP7_75t_L g3784 ( 
.A1(n_3476),
.A2(n_2568),
.B(n_2561),
.Y(n_3784)
);

AO32x2_ASAP7_75t_L g3785 ( 
.A1(n_3552),
.A2(n_10),
.A3(n_3),
.B1(n_8),
.B2(n_11),
.Y(n_3785)
);

OR2x2_ASAP7_75t_L g3786 ( 
.A(n_3504),
.B(n_1241),
.Y(n_3786)
);

OAI21x1_ASAP7_75t_L g3787 ( 
.A1(n_3476),
.A2(n_2573),
.B(n_2568),
.Y(n_3787)
);

A2O1A1Ixp33_ASAP7_75t_L g3788 ( 
.A1(n_3454),
.A2(n_891),
.B(n_892),
.C(n_890),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3446),
.B(n_895),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3472),
.B(n_897),
.Y(n_3790)
);

AO31x2_ASAP7_75t_L g3791 ( 
.A1(n_3587),
.A2(n_2579),
.A3(n_2602),
.B(n_2573),
.Y(n_3791)
);

OAI21x1_ASAP7_75t_L g3792 ( 
.A1(n_3464),
.A2(n_2602),
.B(n_2579),
.Y(n_3792)
);

AO31x2_ASAP7_75t_L g3793 ( 
.A1(n_3510),
.A2(n_2611),
.A3(n_2606),
.B(n_2276),
.Y(n_3793)
);

BUFx10_ASAP7_75t_L g3794 ( 
.A(n_3557),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3512),
.Y(n_3795)
);

AO32x2_ASAP7_75t_L g3796 ( 
.A1(n_3599),
.A2(n_12),
.A3(n_8),
.B1(n_11),
.B2(n_13),
.Y(n_3796)
);

OAI21xp5_ASAP7_75t_L g3797 ( 
.A1(n_3511),
.A2(n_2497),
.B(n_1242),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3427),
.B(n_3519),
.Y(n_3798)
);

OR2x6_ASAP7_75t_L g3799 ( 
.A(n_3603),
.B(n_2606),
.Y(n_3799)
);

A2O1A1Ixp33_ASAP7_75t_L g3800 ( 
.A1(n_3465),
.A2(n_3486),
.B(n_3522),
.C(n_3524),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3525),
.Y(n_3801)
);

OAI21xp5_ASAP7_75t_L g3802 ( 
.A1(n_3471),
.A2(n_1243),
.B(n_1241),
.Y(n_3802)
);

OAI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_3502),
.A2(n_1245),
.B(n_1243),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3482),
.B(n_899),
.Y(n_3804)
);

AOI22xp33_ASAP7_75t_L g3805 ( 
.A1(n_3522),
.A2(n_904),
.B1(n_905),
.B2(n_903),
.Y(n_3805)
);

AOI21xp5_ASAP7_75t_L g3806 ( 
.A1(n_3530),
.A2(n_2611),
.B(n_2313),
.Y(n_3806)
);

AO21x1_ASAP7_75t_L g3807 ( 
.A1(n_3564),
.A2(n_1247),
.B(n_1245),
.Y(n_3807)
);

O2A1O1Ixp33_ASAP7_75t_SL g3808 ( 
.A1(n_3567),
.A2(n_3573),
.B(n_3592),
.C(n_3489),
.Y(n_3808)
);

OAI21xp5_ASAP7_75t_L g3809 ( 
.A1(n_3551),
.A2(n_1249),
.B(n_1247),
.Y(n_3809)
);

OAI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_3487),
.A2(n_1252),
.B(n_1249),
.Y(n_3810)
);

AND2x4_ASAP7_75t_L g3811 ( 
.A(n_3406),
.B(n_2319),
.Y(n_3811)
);

O2A1O1Ixp33_ASAP7_75t_L g3812 ( 
.A1(n_3603),
.A2(n_1257),
.B(n_1258),
.C(n_1252),
.Y(n_3812)
);

AOI21xp5_ASAP7_75t_L g3813 ( 
.A1(n_3575),
.A2(n_2310),
.B(n_2276),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3493),
.B(n_906),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_L g3815 ( 
.A(n_3506),
.B(n_907),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_3576),
.B(n_909),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3547),
.A2(n_2282),
.B(n_2268),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3578),
.Y(n_3818)
);

AOI21xp5_ASAP7_75t_L g3819 ( 
.A1(n_3593),
.A2(n_3559),
.B(n_3475),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3578),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3578),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_3414),
.B(n_910),
.Y(n_3822)
);

OAI21x1_ASAP7_75t_L g3823 ( 
.A1(n_3414),
.A2(n_2296),
.B(n_2285),
.Y(n_3823)
);

AOI221xp5_ASAP7_75t_SL g3824 ( 
.A1(n_3535),
.A2(n_1263),
.B1(n_1264),
.B2(n_1258),
.C(n_1257),
.Y(n_3824)
);

OAI21x1_ASAP7_75t_SL g3825 ( 
.A1(n_3599),
.A2(n_1264),
.B(n_1263),
.Y(n_3825)
);

OAI21x1_ASAP7_75t_L g3826 ( 
.A1(n_3426),
.A2(n_2296),
.B(n_2282),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3559),
.B(n_911),
.Y(n_3827)
);

OAI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3509),
.A2(n_918),
.B1(n_920),
.B2(n_913),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3593),
.A2(n_2286),
.B(n_2268),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3519),
.Y(n_3830)
);

OAI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_3564),
.A2(n_1270),
.B(n_1268),
.Y(n_3831)
);

A2O1A1Ixp33_ASAP7_75t_L g3832 ( 
.A1(n_3593),
.A2(n_923),
.B(n_925),
.C(n_922),
.Y(n_3832)
);

AO31x2_ASAP7_75t_L g3833 ( 
.A1(n_3610),
.A2(n_2291),
.A3(n_2308),
.B(n_2286),
.Y(n_3833)
);

OAI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3445),
.A2(n_1270),
.B(n_1268),
.Y(n_3834)
);

OAI22xp5_ASAP7_75t_L g3835 ( 
.A1(n_3509),
.A2(n_928),
.B1(n_930),
.B2(n_927),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3694),
.B(n_3519),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3733),
.B(n_3535),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3626),
.B(n_3535),
.Y(n_3838)
);

OAI21x1_ASAP7_75t_L g3839 ( 
.A1(n_3668),
.A2(n_3426),
.B(n_3459),
.Y(n_3839)
);

OAI21x1_ASAP7_75t_L g3840 ( 
.A1(n_3633),
.A2(n_2308),
.B(n_2291),
.Y(n_3840)
);

NAND2x1_ASAP7_75t_L g3841 ( 
.A(n_3630),
.B(n_3427),
.Y(n_3841)
);

OAI21x1_ASAP7_75t_L g3842 ( 
.A1(n_3680),
.A2(n_2230),
.B(n_1207),
.Y(n_3842)
);

BUFx8_ASAP7_75t_SL g3843 ( 
.A(n_3706),
.Y(n_3843)
);

OA21x2_ASAP7_75t_L g3844 ( 
.A1(n_3725),
.A2(n_3800),
.B(n_3731),
.Y(n_3844)
);

AOI22xp33_ASAP7_75t_L g3845 ( 
.A1(n_3663),
.A2(n_3475),
.B1(n_3550),
.B2(n_3543),
.Y(n_3845)
);

CKINVDCx16_ASAP7_75t_R g3846 ( 
.A(n_3698),
.Y(n_3846)
);

HB1xp67_ASAP7_75t_L g3847 ( 
.A(n_3640),
.Y(n_3847)
);

OAI21x1_ASAP7_75t_L g3848 ( 
.A1(n_3618),
.A2(n_1207),
.B(n_1203),
.Y(n_3848)
);

OA21x2_ASAP7_75t_L g3849 ( 
.A1(n_3690),
.A2(n_935),
.B(n_933),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3649),
.B(n_3543),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3669),
.Y(n_3851)
);

NAND2x1p5_ASAP7_75t_L g3852 ( 
.A(n_3684),
.B(n_3475),
.Y(n_3852)
);

A2O1A1Ixp33_ASAP7_75t_L g3853 ( 
.A1(n_3705),
.A2(n_3468),
.B(n_941),
.C(n_946),
.Y(n_3853)
);

O2A1O1Ixp33_ASAP7_75t_L g3854 ( 
.A1(n_3628),
.A2(n_1217),
.B(n_1221),
.C(n_1211),
.Y(n_3854)
);

HB1xp67_ASAP7_75t_L g3855 ( 
.A(n_3656),
.Y(n_3855)
);

AO21x2_ASAP7_75t_L g3856 ( 
.A1(n_3722),
.A2(n_1217),
.B(n_1211),
.Y(n_3856)
);

OAI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_3641),
.A2(n_3610),
.B(n_950),
.Y(n_3857)
);

AO31x2_ASAP7_75t_L g3858 ( 
.A1(n_3807),
.A2(n_1226),
.A3(n_1233),
.B(n_1221),
.Y(n_3858)
);

OAI21x1_ASAP7_75t_L g3859 ( 
.A1(n_3659),
.A2(n_1233),
.B(n_1226),
.Y(n_3859)
);

AND2x4_ASAP7_75t_L g3860 ( 
.A(n_3665),
.B(n_3543),
.Y(n_3860)
);

OA21x2_ASAP7_75t_L g3861 ( 
.A1(n_3819),
.A2(n_951),
.B(n_938),
.Y(n_3861)
);

A2O1A1Ixp33_ASAP7_75t_L g3862 ( 
.A1(n_3617),
.A2(n_3550),
.B(n_3442),
.C(n_3452),
.Y(n_3862)
);

NOR2xp33_ASAP7_75t_L g3863 ( 
.A(n_3683),
.B(n_3442),
.Y(n_3863)
);

CKINVDCx20_ASAP7_75t_R g3864 ( 
.A(n_3737),
.Y(n_3864)
);

CKINVDCx5p33_ASAP7_75t_R g3865 ( 
.A(n_3794),
.Y(n_3865)
);

AND2x4_ASAP7_75t_L g3866 ( 
.A(n_3724),
.B(n_3550),
.Y(n_3866)
);

AOI22xp33_ASAP7_75t_SL g3867 ( 
.A1(n_3658),
.A2(n_3452),
.B1(n_2581),
.B2(n_2599),
.Y(n_3867)
);

CKINVDCx5p33_ASAP7_75t_R g3868 ( 
.A(n_3753),
.Y(n_3868)
);

OAI21x1_ASAP7_75t_L g3869 ( 
.A1(n_3716),
.A2(n_1235),
.B(n_1659),
.Y(n_3869)
);

AOI221xp5_ASAP7_75t_L g3870 ( 
.A1(n_3654),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.C(n_16),
.Y(n_3870)
);

BUFx3_ASAP7_75t_L g3871 ( 
.A(n_3664),
.Y(n_3871)
);

OAI21x1_ASAP7_75t_L g3872 ( 
.A1(n_3792),
.A2(n_1235),
.B(n_1659),
.Y(n_3872)
);

NAND3xp33_ASAP7_75t_L g3873 ( 
.A(n_3634),
.B(n_3452),
.C(n_1311),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3745),
.Y(n_3874)
);

AO32x2_ASAP7_75t_L g3875 ( 
.A1(n_3667),
.A2(n_17),
.A3(n_14),
.B1(n_15),
.B2(n_19),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3754),
.Y(n_3876)
);

AOI22xp5_ASAP7_75t_L g3877 ( 
.A1(n_3695),
.A2(n_2564),
.B1(n_2599),
.B2(n_2581),
.Y(n_3877)
);

OAI21x1_ASAP7_75t_L g3878 ( 
.A1(n_3732),
.A2(n_1675),
.B(n_1659),
.Y(n_3878)
);

OAI22xp5_ASAP7_75t_L g3879 ( 
.A1(n_3615),
.A2(n_27),
.B1(n_20),
.B2(n_26),
.Y(n_3879)
);

AOI21xp33_ASAP7_75t_L g3880 ( 
.A1(n_3616),
.A2(n_20),
.B(n_28),
.Y(n_3880)
);

AOI22xp33_ASAP7_75t_L g3881 ( 
.A1(n_3629),
.A2(n_2581),
.B1(n_2599),
.B2(n_2564),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_3759),
.B(n_30),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3760),
.B(n_30),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3761),
.Y(n_3884)
);

OAI21xp5_ASAP7_75t_L g3885 ( 
.A1(n_3703),
.A2(n_2581),
.B(n_2564),
.Y(n_3885)
);

OAI21x1_ASAP7_75t_L g3886 ( 
.A1(n_3741),
.A2(n_1676),
.B(n_1675),
.Y(n_3886)
);

OAI21x1_ASAP7_75t_L g3887 ( 
.A1(n_3746),
.A2(n_1676),
.B(n_1675),
.Y(n_3887)
);

AOI22xp33_ASAP7_75t_SL g3888 ( 
.A1(n_3666),
.A2(n_2581),
.B1(n_2599),
.B2(n_2564),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3795),
.Y(n_3889)
);

INVx2_ASAP7_75t_L g3890 ( 
.A(n_3676),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3777),
.Y(n_3891)
);

AOI21xp5_ASAP7_75t_L g3892 ( 
.A1(n_3650),
.A2(n_2640),
.B(n_2599),
.Y(n_3892)
);

OAI21x1_ASAP7_75t_L g3893 ( 
.A1(n_3670),
.A2(n_1676),
.B(n_1743),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3801),
.Y(n_3894)
);

AND2x4_ASAP7_75t_L g3895 ( 
.A(n_3681),
.B(n_2546),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3818),
.Y(n_3896)
);

OAI22xp5_ASAP7_75t_L g3897 ( 
.A1(n_3696),
.A2(n_3655),
.B1(n_3652),
.B2(n_3622),
.Y(n_3897)
);

NAND2x1p5_ASAP7_75t_L g3898 ( 
.A(n_3764),
.B(n_1091),
.Y(n_3898)
);

OAI22xp33_ASAP7_75t_L g3899 ( 
.A1(n_3653),
.A2(n_1769),
.B1(n_1821),
.B2(n_1783),
.Y(n_3899)
);

AO21x1_ASAP7_75t_L g3900 ( 
.A1(n_3821),
.A2(n_31),
.B(n_33),
.Y(n_3900)
);

AOI221xp5_ASAP7_75t_L g3901 ( 
.A1(n_3646),
.A2(n_34),
.B1(n_31),
.B2(n_33),
.C(n_35),
.Y(n_3901)
);

OAI21x1_ASAP7_75t_L g3902 ( 
.A1(n_3636),
.A2(n_2649),
.B(n_2546),
.Y(n_3902)
);

OAI21xp5_ASAP7_75t_L g3903 ( 
.A1(n_3631),
.A2(n_2646),
.B(n_2640),
.Y(n_3903)
);

INVx8_ASAP7_75t_L g3904 ( 
.A(n_3799),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3721),
.Y(n_3905)
);

AOI21xp5_ASAP7_75t_L g3906 ( 
.A1(n_3806),
.A2(n_2646),
.B(n_2640),
.Y(n_3906)
);

OAI21x1_ASAP7_75t_L g3907 ( 
.A1(n_3823),
.A2(n_2649),
.B(n_2546),
.Y(n_3907)
);

NAND2x1p5_ASAP7_75t_L g3908 ( 
.A(n_3764),
.B(n_1311),
.Y(n_3908)
);

OAI21x1_ASAP7_75t_L g3909 ( 
.A1(n_3826),
.A2(n_3623),
.B(n_3778),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_3820),
.Y(n_3910)
);

O2A1O1Ixp33_ASAP7_75t_L g3911 ( 
.A1(n_3788),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_3911)
);

INVx2_ASAP7_75t_L g3912 ( 
.A(n_3830),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3723),
.Y(n_3913)
);

CKINVDCx20_ASAP7_75t_R g3914 ( 
.A(n_3740),
.Y(n_3914)
);

OAI21x1_ASAP7_75t_L g3915 ( 
.A1(n_3784),
.A2(n_2649),
.B(n_2646),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3798),
.B(n_38),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3718),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3718),
.Y(n_3918)
);

AOI21xp5_ASAP7_75t_L g3919 ( 
.A1(n_3797),
.A2(n_2646),
.B(n_2640),
.Y(n_3919)
);

OAI21x1_ASAP7_75t_L g3920 ( 
.A1(n_3787),
.A2(n_2646),
.B(n_2640),
.Y(n_3920)
);

OAI21x1_ASAP7_75t_L g3921 ( 
.A1(n_3776),
.A2(n_400),
.B(n_399),
.Y(n_3921)
);

BUFx2_ASAP7_75t_L g3922 ( 
.A(n_3673),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3718),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3720),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3720),
.Y(n_3925)
);

OAI21x1_ASAP7_75t_L g3926 ( 
.A1(n_3648),
.A2(n_408),
.B(n_405),
.Y(n_3926)
);

OAI21x1_ASAP7_75t_L g3927 ( 
.A1(n_3762),
.A2(n_411),
.B(n_410),
.Y(n_3927)
);

NAND2x1p5_ASAP7_75t_L g3928 ( 
.A(n_3773),
.B(n_1311),
.Y(n_3928)
);

OAI21x1_ASAP7_75t_L g3929 ( 
.A1(n_3817),
.A2(n_414),
.B(n_413),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3720),
.Y(n_3930)
);

OAI21x1_ASAP7_75t_L g3931 ( 
.A1(n_3825),
.A2(n_3752),
.B(n_3770),
.Y(n_3931)
);

OAI21x1_ASAP7_75t_L g3932 ( 
.A1(n_3763),
.A2(n_419),
.B(n_418),
.Y(n_3932)
);

AOI221xp5_ASAP7_75t_L g3933 ( 
.A1(n_3686),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.C(n_42),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3729),
.Y(n_3934)
);

A2O1A1Ixp33_ASAP7_75t_L g3935 ( 
.A1(n_3620),
.A2(n_43),
.B(n_40),
.C(n_41),
.Y(n_3935)
);

AO31x2_ASAP7_75t_L g3936 ( 
.A1(n_3768),
.A2(n_1664),
.A3(n_46),
.B(n_44),
.Y(n_3936)
);

OAI21x1_ASAP7_75t_L g3937 ( 
.A1(n_3771),
.A2(n_422),
.B(n_421),
.Y(n_3937)
);

NAND2x1p5_ASAP7_75t_L g3938 ( 
.A(n_3709),
.B(n_1311),
.Y(n_3938)
);

OAI21x1_ASAP7_75t_L g3939 ( 
.A1(n_3767),
.A2(n_3781),
.B(n_3697),
.Y(n_3939)
);

OAI22xp5_ASAP7_75t_L g3940 ( 
.A1(n_3651),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3729),
.Y(n_3941)
);

BUFx12f_ASAP7_75t_L g3942 ( 
.A(n_3662),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3729),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3780),
.Y(n_3944)
);

OAI21x1_ASAP7_75t_L g3945 ( 
.A1(n_3717),
.A2(n_425),
.B(n_423),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3643),
.B(n_48),
.Y(n_3946)
);

AOI22x1_ASAP7_75t_L g3947 ( 
.A1(n_3660),
.A2(n_1311),
.B1(n_52),
.B2(n_48),
.Y(n_3947)
);

OAI21x1_ASAP7_75t_L g3948 ( 
.A1(n_3713),
.A2(n_3707),
.B(n_3813),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3780),
.B(n_51),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3780),
.Y(n_3950)
);

AO31x2_ASAP7_75t_L g3951 ( 
.A1(n_3734),
.A2(n_1664),
.A3(n_56),
.B(n_53),
.Y(n_3951)
);

OAI21x1_ASAP7_75t_L g3952 ( 
.A1(n_3772),
.A2(n_427),
.B(n_426),
.Y(n_3952)
);

NOR2xp33_ASAP7_75t_SL g3953 ( 
.A(n_3739),
.B(n_1769),
.Y(n_3953)
);

AOI22xp33_ASAP7_75t_L g3954 ( 
.A1(n_3685),
.A2(n_1821),
.B1(n_1829),
.B2(n_1783),
.Y(n_3954)
);

AO31x2_ASAP7_75t_L g3955 ( 
.A1(n_3675),
.A2(n_58),
.A3(n_54),
.B(n_57),
.Y(n_3955)
);

NOR2xp33_ASAP7_75t_L g3956 ( 
.A(n_3688),
.B(n_3735),
.Y(n_3956)
);

NAND2x1p5_ASAP7_75t_L g3957 ( 
.A(n_3757),
.B(n_1783),
.Y(n_3957)
);

AOI21xp5_ASAP7_75t_L g3958 ( 
.A1(n_3783),
.A2(n_1821),
.B(n_1783),
.Y(n_3958)
);

OAI21x1_ASAP7_75t_L g3959 ( 
.A1(n_3786),
.A2(n_429),
.B(n_428),
.Y(n_3959)
);

OAI21x1_ASAP7_75t_L g3960 ( 
.A1(n_3831),
.A2(n_433),
.B(n_431),
.Y(n_3960)
);

OAI21x1_ASAP7_75t_L g3961 ( 
.A1(n_3677),
.A2(n_435),
.B(n_434),
.Y(n_3961)
);

OAI21x1_ASAP7_75t_L g3962 ( 
.A1(n_3693),
.A2(n_440),
.B(n_436),
.Y(n_3962)
);

OAI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3687),
.A2(n_57),
.B(n_59),
.Y(n_3963)
);

AO31x2_ASAP7_75t_L g3964 ( 
.A1(n_3719),
.A2(n_61),
.A3(n_59),
.B(n_60),
.Y(n_3964)
);

BUFx4f_ASAP7_75t_SL g3965 ( 
.A(n_3715),
.Y(n_3965)
);

OAI21xp5_ASAP7_75t_L g3966 ( 
.A1(n_3758),
.A2(n_62),
.B(n_63),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3642),
.Y(n_3967)
);

OA21x2_ASAP7_75t_L g3968 ( 
.A1(n_3824),
.A2(n_62),
.B(n_63),
.Y(n_3968)
);

OAI21x1_ASAP7_75t_L g3969 ( 
.A1(n_3727),
.A2(n_443),
.B(n_441),
.Y(n_3969)
);

AOI21xp5_ASAP7_75t_L g3970 ( 
.A1(n_3638),
.A2(n_1829),
.B(n_1821),
.Y(n_3970)
);

OAI21x1_ASAP7_75t_L g3971 ( 
.A1(n_3812),
.A2(n_448),
.B(n_447),
.Y(n_3971)
);

OAI21x1_ASAP7_75t_L g3972 ( 
.A1(n_3711),
.A2(n_452),
.B(n_449),
.Y(n_3972)
);

BUFx6f_ASAP7_75t_L g3973 ( 
.A(n_3774),
.Y(n_3973)
);

INVx3_ASAP7_75t_L g3974 ( 
.A(n_3728),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_SL g3975 ( 
.A(n_3704),
.B(n_1829),
.Y(n_3975)
);

A2O1A1Ixp33_ASAP7_75t_L g3976 ( 
.A1(n_3624),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_3976)
);

BUFx2_ASAP7_75t_L g3977 ( 
.A(n_3755),
.Y(n_3977)
);

OA21x2_ASAP7_75t_L g3978 ( 
.A1(n_3802),
.A2(n_64),
.B(n_65),
.Y(n_3978)
);

OAI21x1_ASAP7_75t_L g3979 ( 
.A1(n_3829),
.A2(n_3810),
.B(n_3803),
.Y(n_3979)
);

BUFx2_ASAP7_75t_L g3980 ( 
.A(n_3765),
.Y(n_3980)
);

OAI22x1_ASAP7_75t_L g3981 ( 
.A1(n_3635),
.A2(n_3751),
.B1(n_3766),
.B2(n_3749),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3775),
.Y(n_3982)
);

OAI21x1_ASAP7_75t_L g3983 ( 
.A1(n_3742),
.A2(n_455),
.B(n_454),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3674),
.B(n_66),
.Y(n_3984)
);

BUFx3_ASAP7_75t_L g3985 ( 
.A(n_3715),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_3672),
.Y(n_3986)
);

OAI21x1_ASAP7_75t_L g3987 ( 
.A1(n_3809),
.A2(n_458),
.B(n_457),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_3672),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_3775),
.Y(n_3989)
);

INVx4_ASAP7_75t_L g3990 ( 
.A(n_3774),
.Y(n_3990)
);

OAI21x1_ASAP7_75t_L g3991 ( 
.A1(n_3639),
.A2(n_460),
.B(n_459),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3672),
.Y(n_3992)
);

OAI21x1_ASAP7_75t_L g3993 ( 
.A1(n_3834),
.A2(n_462),
.B(n_461),
.Y(n_3993)
);

OAI21x1_ASAP7_75t_L g3994 ( 
.A1(n_3736),
.A2(n_464),
.B(n_463),
.Y(n_3994)
);

INVx2_ASAP7_75t_SL g3995 ( 
.A(n_3747),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3775),
.Y(n_3996)
);

BUFx2_ASAP7_75t_L g3997 ( 
.A(n_3744),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3625),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3674),
.B(n_67),
.Y(n_3999)
);

NAND2x1p5_ASAP7_75t_L g4000 ( 
.A(n_3747),
.B(n_1829),
.Y(n_4000)
);

AOI22xp33_ASAP7_75t_L g4001 ( 
.A1(n_3714),
.A2(n_1837),
.B1(n_1840),
.B2(n_1830),
.Y(n_4001)
);

OAI21x1_ASAP7_75t_L g4002 ( 
.A1(n_3822),
.A2(n_466),
.B(n_465),
.Y(n_4002)
);

OR2x2_ASAP7_75t_L g4003 ( 
.A(n_3678),
.B(n_67),
.Y(n_4003)
);

OAI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_3632),
.A2(n_68),
.B(n_69),
.Y(n_4004)
);

OAI21x1_ASAP7_75t_L g4005 ( 
.A1(n_3689),
.A2(n_469),
.B(n_468),
.Y(n_4005)
);

NOR2xp33_ASAP7_75t_L g4006 ( 
.A(n_3816),
.B(n_70),
.Y(n_4006)
);

OA21x2_ASAP7_75t_L g4007 ( 
.A1(n_3661),
.A2(n_71),
.B(n_72),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3645),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3678),
.B(n_72),
.Y(n_4009)
);

INVx1_ASAP7_75t_SL g4010 ( 
.A(n_3827),
.Y(n_4010)
);

OA21x2_ASAP7_75t_L g4011 ( 
.A1(n_3671),
.A2(n_73),
.B(n_75),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3645),
.Y(n_4012)
);

BUFx2_ASAP7_75t_L g4013 ( 
.A(n_3974),
.Y(n_4013)
);

AND2x4_ASAP7_75t_L g4014 ( 
.A(n_3860),
.B(n_3644),
.Y(n_4014)
);

OR2x2_ASAP7_75t_L g4015 ( 
.A(n_3847),
.B(n_3699),
.Y(n_4015)
);

NAND2xp33_ASAP7_75t_R g4016 ( 
.A(n_3868),
.B(n_3779),
.Y(n_4016)
);

CKINVDCx5p33_ASAP7_75t_R g4017 ( 
.A(n_3843),
.Y(n_4017)
);

AOI22xp33_ASAP7_75t_L g4018 ( 
.A1(n_3963),
.A2(n_3933),
.B1(n_3956),
.B2(n_3879),
.Y(n_4018)
);

OAI21x1_ASAP7_75t_L g4019 ( 
.A1(n_3948),
.A2(n_3692),
.B(n_3700),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3997),
.B(n_3645),
.Y(n_4020)
);

OR2x2_ASAP7_75t_L g4021 ( 
.A(n_3855),
.B(n_3644),
.Y(n_4021)
);

OR2x6_ASAP7_75t_L g4022 ( 
.A(n_3904),
.B(n_3799),
.Y(n_4022)
);

AOI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_3958),
.A2(n_3808),
.B(n_3637),
.Y(n_4023)
);

OAI22xp5_ASAP7_75t_L g4024 ( 
.A1(n_3845),
.A2(n_3805),
.B1(n_3750),
.B2(n_3789),
.Y(n_4024)
);

OR2x2_ASAP7_75t_L g4025 ( 
.A(n_3836),
.B(n_3837),
.Y(n_4025)
);

INVx3_ASAP7_75t_L g4026 ( 
.A(n_3841),
.Y(n_4026)
);

AOI221xp5_ASAP7_75t_L g4027 ( 
.A1(n_3880),
.A2(n_3782),
.B1(n_3748),
.B2(n_3702),
.C(n_3619),
.Y(n_4027)
);

AOI22xp33_ASAP7_75t_L g4028 ( 
.A1(n_3963),
.A2(n_3679),
.B1(n_3828),
.B2(n_3712),
.Y(n_4028)
);

AOI21x1_ASAP7_75t_L g4029 ( 
.A1(n_3949),
.A2(n_3743),
.B(n_3627),
.Y(n_4029)
);

BUFx2_ASAP7_75t_L g4030 ( 
.A(n_3974),
.Y(n_4030)
);

INVx3_ASAP7_75t_L g4031 ( 
.A(n_3860),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3874),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3905),
.B(n_3726),
.Y(n_4033)
);

OAI21x1_ASAP7_75t_L g4034 ( 
.A1(n_3839),
.A2(n_3804),
.B(n_3790),
.Y(n_4034)
);

AOI22xp5_ASAP7_75t_L g4035 ( 
.A1(n_3933),
.A2(n_3708),
.B1(n_3815),
.B2(n_3814),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3876),
.Y(n_4036)
);

INVx3_ASAP7_75t_L g4037 ( 
.A(n_3866),
.Y(n_4037)
);

AOI21xp5_ASAP7_75t_L g4038 ( 
.A1(n_3958),
.A2(n_3730),
.B(n_3691),
.Y(n_4038)
);

AOI22xp33_ASAP7_75t_L g4039 ( 
.A1(n_3879),
.A2(n_3835),
.B1(n_3811),
.B2(n_3756),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3884),
.Y(n_4040)
);

AND2x4_ASAP7_75t_L g4041 ( 
.A(n_3866),
.B(n_3644),
.Y(n_4041)
);

OR2x2_ASAP7_75t_L g4042 ( 
.A(n_3836),
.B(n_3621),
.Y(n_4042)
);

AOI32xp33_ASAP7_75t_L g4043 ( 
.A1(n_3940),
.A2(n_3785),
.A3(n_3796),
.B1(n_3701),
.B2(n_78),
.Y(n_4043)
);

A2O1A1Ixp33_ASAP7_75t_L g4044 ( 
.A1(n_3853),
.A2(n_3832),
.B(n_3785),
.C(n_3796),
.Y(n_4044)
);

NOR3xp33_ASAP7_75t_SL g4045 ( 
.A(n_3865),
.B(n_3710),
.C(n_3769),
.Y(n_4045)
);

INVx1_ASAP7_75t_SL g4046 ( 
.A(n_4010),
.Y(n_4046)
);

NAND2x1_ASAP7_75t_L g4047 ( 
.A(n_3844),
.B(n_3701),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3922),
.B(n_3647),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3889),
.Y(n_4049)
);

OR2x2_ASAP7_75t_L g4050 ( 
.A(n_3837),
.B(n_3621),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3891),
.Y(n_4051)
);

AND2x2_ASAP7_75t_L g4052 ( 
.A(n_3980),
.B(n_3647),
.Y(n_4052)
);

BUFx2_ASAP7_75t_L g4053 ( 
.A(n_3942),
.Y(n_4053)
);

INVx3_ASAP7_75t_L g4054 ( 
.A(n_3896),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3851),
.Y(n_4055)
);

HB1xp67_ASAP7_75t_L g4056 ( 
.A(n_3944),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3913),
.B(n_3647),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3890),
.Y(n_4058)
);

AND2x4_ASAP7_75t_L g4059 ( 
.A(n_3910),
.B(n_3657),
.Y(n_4059)
);

BUFx2_ASAP7_75t_L g4060 ( 
.A(n_3990),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3894),
.B(n_3657),
.Y(n_4061)
);

CKINVDCx6p67_ASAP7_75t_R g4062 ( 
.A(n_3871),
.Y(n_4062)
);

INVx2_ASAP7_75t_SL g4063 ( 
.A(n_3977),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_4010),
.B(n_3657),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3838),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_3912),
.B(n_3701),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_3838),
.Y(n_4067)
);

OAI22xp5_ASAP7_75t_L g4068 ( 
.A1(n_3862),
.A2(n_3785),
.B1(n_3796),
.B2(n_3682),
.Y(n_4068)
);

O2A1O1Ixp5_ASAP7_75t_L g4069 ( 
.A1(n_3900),
.A2(n_3738),
.B(n_3682),
.C(n_78),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3850),
.B(n_3738),
.Y(n_4070)
);

INVxp33_ASAP7_75t_L g4071 ( 
.A(n_3863),
.Y(n_4071)
);

A2O1A1Ixp33_ASAP7_75t_L g4072 ( 
.A1(n_3911),
.A2(n_80),
.B(n_73),
.C(n_77),
.Y(n_4072)
);

OAI22xp5_ASAP7_75t_L g4073 ( 
.A1(n_3873),
.A2(n_3833),
.B1(n_3621),
.B2(n_3791),
.Y(n_4073)
);

OAI22xp5_ASAP7_75t_L g4074 ( 
.A1(n_3873),
.A2(n_3833),
.B1(n_3791),
.B2(n_3793),
.Y(n_4074)
);

NOR3xp33_ASAP7_75t_SL g4075 ( 
.A(n_3949),
.B(n_77),
.C(n_81),
.Y(n_4075)
);

INVx4_ASAP7_75t_SL g4076 ( 
.A(n_3965),
.Y(n_4076)
);

INVx4_ASAP7_75t_L g4077 ( 
.A(n_3973),
.Y(n_4077)
);

BUFx12f_ASAP7_75t_L g4078 ( 
.A(n_3946),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_3850),
.Y(n_4079)
);

BUFx12f_ASAP7_75t_L g4080 ( 
.A(n_3916),
.Y(n_4080)
);

BUFx2_ASAP7_75t_L g4081 ( 
.A(n_3990),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3950),
.Y(n_4082)
);

OAI22xp5_ASAP7_75t_L g4083 ( 
.A1(n_3901),
.A2(n_3833),
.B1(n_3793),
.B2(n_1837),
.Y(n_4083)
);

OAI221xp5_ASAP7_75t_L g4084 ( 
.A1(n_3935),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.C(n_84),
.Y(n_4084)
);

AOI21x1_ASAP7_75t_L g4085 ( 
.A1(n_3882),
.A2(n_3793),
.B(n_82),
.Y(n_4085)
);

AOI22xp33_ASAP7_75t_L g4086 ( 
.A1(n_3940),
.A2(n_1837),
.B1(n_1840),
.B2(n_1830),
.Y(n_4086)
);

AND2x2_ASAP7_75t_L g4087 ( 
.A(n_3998),
.B(n_83),
.Y(n_4087)
);

AOI21xp33_ASAP7_75t_L g4088 ( 
.A1(n_3861),
.A2(n_84),
.B(n_85),
.Y(n_4088)
);

BUFx6f_ASAP7_75t_L g4089 ( 
.A(n_3973),
.Y(n_4089)
);

OAI221xp5_ASAP7_75t_SL g4090 ( 
.A1(n_3976),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.C(n_92),
.Y(n_4090)
);

AOI21xp5_ASAP7_75t_L g4091 ( 
.A1(n_3857),
.A2(n_1837),
.B(n_1830),
.Y(n_4091)
);

INVx2_ASAP7_75t_L g4092 ( 
.A(n_3852),
.Y(n_4092)
);

AOI22xp33_ASAP7_75t_L g4093 ( 
.A1(n_3870),
.A2(n_1840),
.B1(n_1842),
.B2(n_1830),
.Y(n_4093)
);

OAI22xp5_ASAP7_75t_L g4094 ( 
.A1(n_3901),
.A2(n_1842),
.B1(n_1861),
.B2(n_1840),
.Y(n_4094)
);

OAI22xp5_ASAP7_75t_L g4095 ( 
.A1(n_3867),
.A2(n_1861),
.B1(n_1842),
.B2(n_95),
.Y(n_4095)
);

OR2x2_ASAP7_75t_L g4096 ( 
.A(n_3967),
.B(n_90),
.Y(n_4096)
);

OAI21x1_ASAP7_75t_L g4097 ( 
.A1(n_3939),
.A2(n_94),
.B(n_96),
.Y(n_4097)
);

INVx4_ASAP7_75t_L g4098 ( 
.A(n_3973),
.Y(n_4098)
);

AOI21xp5_ASAP7_75t_SL g4099 ( 
.A1(n_3861),
.A2(n_3978),
.B(n_4011),
.Y(n_4099)
);

AND2x2_ASAP7_75t_L g4100 ( 
.A(n_3846),
.B(n_94),
.Y(n_4100)
);

AND2x2_ASAP7_75t_L g4101 ( 
.A(n_3985),
.B(n_97),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3852),
.Y(n_4102)
);

HB1xp67_ASAP7_75t_L g4103 ( 
.A(n_4008),
.Y(n_4103)
);

NOR3xp33_ASAP7_75t_SL g4104 ( 
.A(n_3897),
.B(n_98),
.C(n_100),
.Y(n_4104)
);

AOI22xp33_ASAP7_75t_SL g4105 ( 
.A1(n_3947),
.A2(n_4011),
.B1(n_4007),
.B2(n_3966),
.Y(n_4105)
);

NAND3xp33_ASAP7_75t_SL g4106 ( 
.A(n_4004),
.B(n_101),
.C(n_102),
.Y(n_4106)
);

BUFx3_ASAP7_75t_L g4107 ( 
.A(n_3864),
.Y(n_4107)
);

AOI221xp5_ASAP7_75t_L g4108 ( 
.A1(n_3880),
.A2(n_3870),
.B1(n_4004),
.B2(n_4006),
.C(n_3966),
.Y(n_4108)
);

INVx2_ASAP7_75t_L g4109 ( 
.A(n_3986),
.Y(n_4109)
);

AOI22xp33_ASAP7_75t_L g4110 ( 
.A1(n_3885),
.A2(n_1861),
.B1(n_1842),
.B2(n_1695),
.Y(n_4110)
);

NAND3xp33_ASAP7_75t_SL g4111 ( 
.A(n_3885),
.B(n_103),
.C(n_104),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_3988),
.Y(n_4112)
);

AOI211xp5_ASAP7_75t_L g4113 ( 
.A1(n_3897),
.A2(n_106),
.B(n_103),
.C(n_105),
.Y(n_4113)
);

AO21x2_ASAP7_75t_L g4114 ( 
.A1(n_3992),
.A2(n_107),
.B(n_108),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_4012),
.Y(n_4115)
);

AOI22xp5_ASAP7_75t_L g4116 ( 
.A1(n_4007),
.A2(n_1861),
.B1(n_112),
.B2(n_109),
.Y(n_4116)
);

AOI22xp33_ASAP7_75t_L g4117 ( 
.A1(n_3981),
.A2(n_3857),
.B1(n_3978),
.B2(n_4003),
.Y(n_4117)
);

AND2x4_ASAP7_75t_L g4118 ( 
.A(n_3995),
.B(n_109),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_3844),
.Y(n_4119)
);

AND2x4_ASAP7_75t_L g4120 ( 
.A(n_3895),
.B(n_110),
.Y(n_4120)
);

OAI22xp5_ASAP7_75t_L g4121 ( 
.A1(n_3968),
.A2(n_113),
.B1(n_110),
.B2(n_112),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3882),
.Y(n_4122)
);

HB1xp67_ASAP7_75t_L g4123 ( 
.A(n_3883),
.Y(n_4123)
);

OAI22xp5_ASAP7_75t_L g4124 ( 
.A1(n_3877),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3883),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_SL g4126 ( 
.A(n_3914),
.B(n_1691),
.Y(n_4126)
);

OR2x2_ASAP7_75t_L g4127 ( 
.A(n_3982),
.B(n_116),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3917),
.Y(n_4128)
);

INVxp67_ASAP7_75t_SL g4129 ( 
.A(n_3938),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3918),
.Y(n_4130)
);

AND2x4_ASAP7_75t_L g4131 ( 
.A(n_3895),
.B(n_117),
.Y(n_4131)
);

NAND2xp33_ASAP7_75t_R g4132 ( 
.A(n_3968),
.B(n_119),
.Y(n_4132)
);

O2A1O1Ixp33_ASAP7_75t_L g4133 ( 
.A1(n_3984),
.A2(n_123),
.B(n_119),
.C(n_120),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3984),
.B(n_124),
.Y(n_4134)
);

NAND2x1p5_ASAP7_75t_L g4135 ( 
.A(n_3975),
.B(n_1636),
.Y(n_4135)
);

CKINVDCx16_ASAP7_75t_R g4136 ( 
.A(n_3953),
.Y(n_4136)
);

INVx4_ASAP7_75t_L g4137 ( 
.A(n_3938),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3923),
.Y(n_4138)
);

AOI22xp5_ASAP7_75t_L g4139 ( 
.A1(n_3999),
.A2(n_4009),
.B1(n_3899),
.B2(n_3877),
.Y(n_4139)
);

OAI22xp5_ASAP7_75t_L g4140 ( 
.A1(n_3888),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3999),
.B(n_126),
.Y(n_4141)
);

CKINVDCx8_ASAP7_75t_R g4142 ( 
.A(n_3904),
.Y(n_4142)
);

OR2x2_ASAP7_75t_L g4143 ( 
.A(n_3989),
.B(n_127),
.Y(n_4143)
);

AOI22xp33_ASAP7_75t_SL g4144 ( 
.A1(n_4009),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_4144)
);

AOI21x1_ASAP7_75t_L g4145 ( 
.A1(n_3970),
.A2(n_128),
.B(n_129),
.Y(n_4145)
);

AND2x4_ASAP7_75t_L g4146 ( 
.A(n_3924),
.B(n_130),
.Y(n_4146)
);

CKINVDCx8_ASAP7_75t_R g4147 ( 
.A(n_3904),
.Y(n_4147)
);

AOI222xp33_ASAP7_75t_L g4148 ( 
.A1(n_4001),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.C1(n_135),
.C2(n_137),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_4082),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_L g4150 ( 
.A(n_4046),
.B(n_3955),
.Y(n_4150)
);

AOI21xp5_ASAP7_75t_L g4151 ( 
.A1(n_4091),
.A2(n_3906),
.B(n_3970),
.Y(n_4151)
);

AOI222xp33_ASAP7_75t_L g4152 ( 
.A1(n_4108),
.A2(n_3954),
.B1(n_4002),
.B2(n_3875),
.C1(n_3994),
.C2(n_4005),
.Y(n_4152)
);

AOI22xp33_ASAP7_75t_L g4153 ( 
.A1(n_4018),
.A2(n_3849),
.B1(n_3979),
.B2(n_3919),
.Y(n_4153)
);

AOI22xp33_ASAP7_75t_L g4154 ( 
.A1(n_4106),
.A2(n_3849),
.B1(n_3906),
.B2(n_3856),
.Y(n_4154)
);

OAI22xp5_ASAP7_75t_L g4155 ( 
.A1(n_4044),
.A2(n_3928),
.B1(n_3957),
.B2(n_3881),
.Y(n_4155)
);

OR2x6_ASAP7_75t_L g4156 ( 
.A(n_4099),
.B(n_3928),
.Y(n_4156)
);

CKINVDCx9p33_ASAP7_75t_R g4157 ( 
.A(n_4053),
.Y(n_4157)
);

AOI221xp5_ASAP7_75t_L g4158 ( 
.A1(n_4113),
.A2(n_3996),
.B1(n_3925),
.B2(n_3941),
.C(n_3934),
.Y(n_4158)
);

OAI221xp5_ASAP7_75t_L g4159 ( 
.A1(n_4117),
.A2(n_3953),
.B1(n_3903),
.B2(n_3957),
.C(n_3892),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_4032),
.Y(n_4160)
);

INVx2_ASAP7_75t_L g4161 ( 
.A(n_4092),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4036),
.Y(n_4162)
);

OAI21xp33_ASAP7_75t_L g4163 ( 
.A1(n_4075),
.A2(n_3971),
.B(n_3991),
.Y(n_4163)
);

INVx5_ASAP7_75t_L g4164 ( 
.A(n_4137),
.Y(n_4164)
);

BUFx2_ASAP7_75t_L g4165 ( 
.A(n_4013),
.Y(n_4165)
);

OAI21x1_ASAP7_75t_L g4166 ( 
.A1(n_4119),
.A2(n_3943),
.B(n_3930),
.Y(n_4166)
);

AND2x4_ASAP7_75t_L g4167 ( 
.A(n_4026),
.B(n_3931),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_4040),
.Y(n_4168)
);

OAI22xp33_ASAP7_75t_L g4169 ( 
.A1(n_4116),
.A2(n_3892),
.B1(n_3908),
.B2(n_3898),
.Y(n_4169)
);

AOI22xp33_ASAP7_75t_L g4170 ( 
.A1(n_4084),
.A2(n_3856),
.B1(n_3987),
.B2(n_3960),
.Y(n_4170)
);

A2O1A1Ixp33_ASAP7_75t_L g4171 ( 
.A1(n_4113),
.A2(n_3929),
.B(n_3993),
.C(n_3926),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_4102),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_4046),
.B(n_3955),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4049),
.Y(n_4174)
);

NOR2xp33_ASAP7_75t_L g4175 ( 
.A(n_4017),
.B(n_3972),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_4054),
.Y(n_4176)
);

OAI22xp5_ASAP7_75t_L g4177 ( 
.A1(n_4043),
.A2(n_3908),
.B1(n_3898),
.B2(n_3903),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_4123),
.B(n_3955),
.Y(n_4178)
);

AOI22xp33_ASAP7_75t_L g4179 ( 
.A1(n_4105),
.A2(n_3932),
.B1(n_3962),
.B2(n_3961),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_4065),
.B(n_3964),
.Y(n_4180)
);

OAI22xp5_ASAP7_75t_L g4181 ( 
.A1(n_4043),
.A2(n_3875),
.B1(n_4000),
.B2(n_3936),
.Y(n_4181)
);

BUFx6f_ASAP7_75t_L g4182 ( 
.A(n_4089),
.Y(n_4182)
);

NOR2x1_ASAP7_75t_SL g4183 ( 
.A(n_4020),
.B(n_3875),
.Y(n_4183)
);

HB1xp67_ASAP7_75t_L g4184 ( 
.A(n_4064),
.Y(n_4184)
);

OA21x2_ASAP7_75t_L g4185 ( 
.A1(n_4130),
.A2(n_3909),
.B(n_3886),
.Y(n_4185)
);

AOI22xp5_ASAP7_75t_L g4186 ( 
.A1(n_4104),
.A2(n_3959),
.B1(n_3945),
.B2(n_3937),
.Y(n_4186)
);

OAI221xp5_ASAP7_75t_L g4187 ( 
.A1(n_4133),
.A2(n_3854),
.B1(n_4000),
.B2(n_3936),
.C(n_3964),
.Y(n_4187)
);

OAI321xp33_ASAP7_75t_L g4188 ( 
.A1(n_4090),
.A2(n_3936),
.A3(n_3964),
.B1(n_141),
.B2(n_142),
.C(n_143),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_4051),
.Y(n_4189)
);

AOI22xp5_ASAP7_75t_L g4190 ( 
.A1(n_4111),
.A2(n_3952),
.B1(n_3969),
.B2(n_3983),
.Y(n_4190)
);

A2O1A1Ixp33_ASAP7_75t_L g4191 ( 
.A1(n_4072),
.A2(n_4116),
.B(n_4088),
.C(n_4023),
.Y(n_4191)
);

OAI22xp33_ASAP7_75t_L g4192 ( 
.A1(n_4132),
.A2(n_3902),
.B1(n_3858),
.B2(n_3927),
.Y(n_4192)
);

BUFx12f_ASAP7_75t_L g4193 ( 
.A(n_4100),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4056),
.Y(n_4194)
);

AOI22xp33_ASAP7_75t_L g4195 ( 
.A1(n_4028),
.A2(n_4094),
.B1(n_4024),
.B2(n_4027),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_4054),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_4025),
.Y(n_4197)
);

AOI22xp33_ASAP7_75t_SL g4198 ( 
.A1(n_4068),
.A2(n_3921),
.B1(n_3869),
.B2(n_3842),
.Y(n_4198)
);

HB1xp67_ASAP7_75t_L g4199 ( 
.A(n_4057),
.Y(n_4199)
);

INVx2_ASAP7_75t_SL g4200 ( 
.A(n_4062),
.Y(n_4200)
);

AOI21xp33_ASAP7_75t_L g4201 ( 
.A1(n_4019),
.A2(n_4047),
.B(n_4034),
.Y(n_4201)
);

AOI22xp33_ASAP7_75t_L g4202 ( 
.A1(n_4038),
.A2(n_3872),
.B1(n_3859),
.B2(n_3893),
.Y(n_4202)
);

AOI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_4121),
.A2(n_3887),
.B(n_3878),
.Y(n_4203)
);

BUFx3_ASAP7_75t_L g4204 ( 
.A(n_4107),
.Y(n_4204)
);

BUFx2_ASAP7_75t_L g4205 ( 
.A(n_4030),
.Y(n_4205)
);

AND2x4_ASAP7_75t_L g4206 ( 
.A(n_4026),
.B(n_3920),
.Y(n_4206)
);

BUFx8_ASAP7_75t_SL g4207 ( 
.A(n_4120),
.Y(n_4207)
);

AOI22xp33_ASAP7_75t_L g4208 ( 
.A1(n_4148),
.A2(n_3907),
.B1(n_3848),
.B2(n_3915),
.Y(n_4208)
);

INVx2_ASAP7_75t_SL g4209 ( 
.A(n_4063),
.Y(n_4209)
);

OR2x2_ASAP7_75t_L g4210 ( 
.A(n_4050),
.B(n_3951),
.Y(n_4210)
);

OA21x2_ASAP7_75t_L g4211 ( 
.A1(n_4138),
.A2(n_3840),
.B(n_3951),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_4031),
.Y(n_4212)
);

INVx4_ASAP7_75t_L g4213 ( 
.A(n_4076),
.Y(n_4213)
);

NOR2xp33_ASAP7_75t_L g4214 ( 
.A(n_4033),
.B(n_137),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_4067),
.B(n_3951),
.Y(n_4215)
);

OAI211xp5_ASAP7_75t_L g4216 ( 
.A1(n_4144),
.A2(n_146),
.B(n_140),
.C(n_142),
.Y(n_4216)
);

AOI21x1_ASAP7_75t_L g4217 ( 
.A1(n_4029),
.A2(n_3858),
.B(n_140),
.Y(n_4217)
);

AND2x2_ASAP7_75t_L g4218 ( 
.A(n_4031),
.B(n_3858),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4055),
.Y(n_4219)
);

A2O1A1Ixp33_ASAP7_75t_L g4220 ( 
.A1(n_4035),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4058),
.Y(n_4221)
);

INVxp67_ASAP7_75t_SL g4222 ( 
.A(n_4070),
.Y(n_4222)
);

AOI222xp33_ASAP7_75t_L g4223 ( 
.A1(n_4134),
.A2(n_149),
.B1(n_150),
.B2(n_155),
.C1(n_156),
.C2(n_157),
.Y(n_4223)
);

OAI22xp5_ASAP7_75t_L g4224 ( 
.A1(n_4139),
.A2(n_155),
.B1(n_149),
.B2(n_150),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_4079),
.B(n_157),
.Y(n_4225)
);

AOI22xp33_ASAP7_75t_L g4226 ( 
.A1(n_4148),
.A2(n_1695),
.B1(n_1691),
.B2(n_1641),
.Y(n_4226)
);

OAI221xp5_ASAP7_75t_L g4227 ( 
.A1(n_4035),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.C(n_161),
.Y(n_4227)
);

AOI221xp5_ASAP7_75t_L g4228 ( 
.A1(n_4141),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.C(n_162),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_4122),
.B(n_162),
.Y(n_4229)
);

AOI22xp33_ASAP7_75t_SL g4230 ( 
.A1(n_4121),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_4230)
);

AOI22xp33_ASAP7_75t_L g4231 ( 
.A1(n_4071),
.A2(n_1695),
.B1(n_1691),
.B2(n_1641),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_4125),
.B(n_167),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_4115),
.Y(n_4233)
);

OAI22xp33_ASAP7_75t_L g4234 ( 
.A1(n_4139),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_4234)
);

AOI22xp33_ASAP7_75t_SL g4235 ( 
.A1(n_4136),
.A2(n_4124),
.B1(n_4095),
.B2(n_4140),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4103),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_4015),
.B(n_169),
.Y(n_4237)
);

OAI22xp33_ASAP7_75t_L g4238 ( 
.A1(n_4022),
.A2(n_173),
.B1(n_170),
.B2(n_171),
.Y(n_4238)
);

AND2x2_ASAP7_75t_L g4239 ( 
.A(n_4037),
.B(n_4060),
.Y(n_4239)
);

NAND2x1_ASAP7_75t_L g4240 ( 
.A(n_4014),
.B(n_4041),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4128),
.Y(n_4241)
);

AOI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_4093),
.A2(n_1695),
.B1(n_1641),
.B2(n_1652),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_4066),
.B(n_174),
.Y(n_4243)
);

OAI221xp5_ASAP7_75t_L g4244 ( 
.A1(n_4142),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.C(n_179),
.Y(n_4244)
);

INVx2_ASAP7_75t_L g4245 ( 
.A(n_4037),
.Y(n_4245)
);

OA21x2_ASAP7_75t_L g4246 ( 
.A1(n_4109),
.A2(n_179),
.B(n_180),
.Y(n_4246)
);

OAI21x1_ASAP7_75t_L g4247 ( 
.A1(n_4061),
.A2(n_180),
.B(n_182),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_4081),
.Y(n_4248)
);

OAI221xp5_ASAP7_75t_SL g4249 ( 
.A1(n_4086),
.A2(n_182),
.B1(n_183),
.B2(n_185),
.C(n_186),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4052),
.B(n_187),
.Y(n_4250)
);

AND2x2_ASAP7_75t_L g4251 ( 
.A(n_4048),
.B(n_187),
.Y(n_4251)
);

OR2x2_ASAP7_75t_SL g4252 ( 
.A(n_4096),
.B(n_188),
.Y(n_4252)
);

AOI22xp5_ASAP7_75t_L g4253 ( 
.A1(n_4045),
.A2(n_191),
.B1(n_188),
.B2(n_189),
.Y(n_4253)
);

CKINVDCx20_ASAP7_75t_R g4254 ( 
.A(n_4076),
.Y(n_4254)
);

AOI22xp5_ASAP7_75t_L g4255 ( 
.A1(n_4120),
.A2(n_194),
.B1(n_191),
.B2(n_193),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4021),
.Y(n_4256)
);

AOI211xp5_ASAP7_75t_L g4257 ( 
.A1(n_4097),
.A2(n_199),
.B(n_196),
.C(n_197),
.Y(n_4257)
);

BUFx2_ASAP7_75t_L g4258 ( 
.A(n_4077),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4127),
.Y(n_4259)
);

INVxp67_ASAP7_75t_SL g4260 ( 
.A(n_4129),
.Y(n_4260)
);

INVx2_ASAP7_75t_SL g4261 ( 
.A(n_4089),
.Y(n_4261)
);

AOI222xp33_ASAP7_75t_L g4262 ( 
.A1(n_4087),
.A2(n_196),
.B1(n_199),
.B2(n_200),
.C1(n_201),
.C2(n_202),
.Y(n_4262)
);

BUFx6f_ASAP7_75t_L g4263 ( 
.A(n_4089),
.Y(n_4263)
);

INVx6_ASAP7_75t_L g4264 ( 
.A(n_4078),
.Y(n_4264)
);

AOI221xp5_ASAP7_75t_L g4265 ( 
.A1(n_4069),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.C(n_206),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_4059),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4042),
.B(n_205),
.Y(n_4267)
);

NOR2xp33_ASAP7_75t_SL g4268 ( 
.A(n_4147),
.B(n_4077),
.Y(n_4268)
);

OAI21xp33_ASAP7_75t_L g4269 ( 
.A1(n_4143),
.A2(n_206),
.B(n_209),
.Y(n_4269)
);

BUFx2_ASAP7_75t_L g4270 ( 
.A(n_4098),
.Y(n_4270)
);

OR2x2_ASAP7_75t_L g4271 ( 
.A(n_4014),
.B(n_209),
.Y(n_4271)
);

AO31x2_ASAP7_75t_L g4272 ( 
.A1(n_4112),
.A2(n_210),
.A3(n_212),
.B(n_213),
.Y(n_4272)
);

AOI221xp5_ASAP7_75t_L g4273 ( 
.A1(n_4146),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.C(n_216),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4267),
.B(n_4146),
.Y(n_4274)
);

INVxp67_ASAP7_75t_L g4275 ( 
.A(n_4271),
.Y(n_4275)
);

BUFx3_ASAP7_75t_L g4276 ( 
.A(n_4254),
.Y(n_4276)
);

AND2x2_ASAP7_75t_L g4277 ( 
.A(n_4239),
.B(n_4041),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4189),
.Y(n_4278)
);

NAND2xp33_ASAP7_75t_R g4279 ( 
.A(n_4258),
.B(n_4118),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4160),
.Y(n_4280)
);

AND2x4_ASAP7_75t_L g4281 ( 
.A(n_4164),
.B(n_4022),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_4260),
.B(n_4101),
.Y(n_4282)
);

AND2x2_ASAP7_75t_L g4283 ( 
.A(n_4197),
.B(n_4098),
.Y(n_4283)
);

NOR2xp33_ASAP7_75t_R g4284 ( 
.A(n_4213),
.B(n_4016),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4182),
.Y(n_4285)
);

XNOR2xp5_ASAP7_75t_L g4286 ( 
.A(n_4200),
.B(n_4252),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_4250),
.B(n_4118),
.Y(n_4287)
);

NOR2xp67_ASAP7_75t_L g4288 ( 
.A(n_4213),
.B(n_4137),
.Y(n_4288)
);

NAND2xp33_ASAP7_75t_R g4289 ( 
.A(n_4270),
.B(n_4246),
.Y(n_4289)
);

NAND2xp33_ASAP7_75t_R g4290 ( 
.A(n_4246),
.B(n_4131),
.Y(n_4290)
);

OR2x6_ASAP7_75t_L g4291 ( 
.A(n_4264),
.B(n_4022),
.Y(n_4291)
);

AND2x2_ASAP7_75t_L g4292 ( 
.A(n_4248),
.B(n_4059),
.Y(n_4292)
);

XNOR2xp5_ASAP7_75t_L g4293 ( 
.A(n_4204),
.B(n_4131),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4162),
.Y(n_4294)
);

XNOR2xp5_ASAP7_75t_L g4295 ( 
.A(n_4253),
.B(n_4039),
.Y(n_4295)
);

NAND2xp33_ASAP7_75t_R g4296 ( 
.A(n_4157),
.B(n_214),
.Y(n_4296)
);

NOR2xp33_ASAP7_75t_R g4297 ( 
.A(n_4268),
.B(n_4080),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4168),
.Y(n_4298)
);

AND2x4_ASAP7_75t_L g4299 ( 
.A(n_4164),
.B(n_4114),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4182),
.Y(n_4300)
);

NAND2xp33_ASAP7_75t_R g4301 ( 
.A(n_4251),
.B(n_217),
.Y(n_4301)
);

INVx2_ASAP7_75t_L g4302 ( 
.A(n_4182),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_4263),
.Y(n_4303)
);

XOR2xp5_ASAP7_75t_L g4304 ( 
.A(n_4235),
.B(n_4126),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_SL g4305 ( 
.A(n_4164),
.B(n_4085),
.Y(n_4305)
);

NAND2xp33_ASAP7_75t_R g4306 ( 
.A(n_4243),
.B(n_217),
.Y(n_4306)
);

NOR2xp33_ASAP7_75t_L g4307 ( 
.A(n_4264),
.B(n_4145),
.Y(n_4307)
);

OR2x6_ASAP7_75t_L g4308 ( 
.A(n_4193),
.B(n_4135),
.Y(n_4308)
);

NOR2xp33_ASAP7_75t_R g4309 ( 
.A(n_4175),
.B(n_218),
.Y(n_4309)
);

CKINVDCx5p33_ASAP7_75t_R g4310 ( 
.A(n_4207),
.Y(n_4310)
);

NAND2xp33_ASAP7_75t_R g4311 ( 
.A(n_4156),
.B(n_219),
.Y(n_4311)
);

XNOR2xp5_ASAP7_75t_L g4312 ( 
.A(n_4253),
.B(n_4255),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_4195),
.B(n_4114),
.Y(n_4313)
);

CKINVDCx20_ASAP7_75t_R g4314 ( 
.A(n_4209),
.Y(n_4314)
);

AND2x4_ASAP7_75t_L g4315 ( 
.A(n_4165),
.B(n_4205),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_L g4316 ( 
.A(n_4259),
.B(n_4083),
.Y(n_4316)
);

BUFx3_ASAP7_75t_L g4317 ( 
.A(n_4261),
.Y(n_4317)
);

INVxp67_ASAP7_75t_L g4318 ( 
.A(n_4178),
.Y(n_4318)
);

NOR2xp33_ASAP7_75t_L g4319 ( 
.A(n_4214),
.B(n_219),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4174),
.Y(n_4320)
);

AND2x2_ASAP7_75t_L g4321 ( 
.A(n_4212),
.B(n_4074),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_4222),
.B(n_4110),
.Y(n_4322)
);

NOR2xp33_ASAP7_75t_R g4323 ( 
.A(n_4237),
.B(n_220),
.Y(n_4323)
);

NAND2xp33_ASAP7_75t_R g4324 ( 
.A(n_4156),
.B(n_220),
.Y(n_4324)
);

INVxp67_ASAP7_75t_L g4325 ( 
.A(n_4247),
.Y(n_4325)
);

BUFx10_ASAP7_75t_L g4326 ( 
.A(n_4263),
.Y(n_4326)
);

NAND2xp33_ASAP7_75t_R g4327 ( 
.A(n_4225),
.B(n_222),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_4263),
.Y(n_4328)
);

INVx2_ASAP7_75t_L g4329 ( 
.A(n_4245),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_4229),
.B(n_4073),
.Y(n_4330)
);

INVxp67_ASAP7_75t_L g4331 ( 
.A(n_4232),
.Y(n_4331)
);

NAND2xp33_ASAP7_75t_R g4332 ( 
.A(n_4150),
.B(n_222),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4149),
.Y(n_4333)
);

AND2x4_ASAP7_75t_L g4334 ( 
.A(n_4236),
.B(n_223),
.Y(n_4334)
);

XNOR2xp5_ASAP7_75t_L g4335 ( 
.A(n_4255),
.B(n_223),
.Y(n_4335)
);

BUFx3_ASAP7_75t_L g4336 ( 
.A(n_4240),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_4173),
.B(n_225),
.Y(n_4337)
);

AND2x4_ASAP7_75t_L g4338 ( 
.A(n_4194),
.B(n_226),
.Y(n_4338)
);

AND2x4_ASAP7_75t_L g4339 ( 
.A(n_4167),
.B(n_227),
.Y(n_4339)
);

NAND2xp33_ASAP7_75t_R g4340 ( 
.A(n_4167),
.B(n_4180),
.Y(n_4340)
);

XNOR2xp5_ASAP7_75t_L g4341 ( 
.A(n_4224),
.B(n_228),
.Y(n_4341)
);

INVx3_ASAP7_75t_L g4342 ( 
.A(n_4266),
.Y(n_4342)
);

NOR2xp33_ASAP7_75t_R g4343 ( 
.A(n_4217),
.B(n_229),
.Y(n_4343)
);

NOR2xp33_ASAP7_75t_L g4344 ( 
.A(n_4163),
.B(n_230),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_SL g4345 ( 
.A(n_4163),
.B(n_1636),
.Y(n_4345)
);

OR2x2_ASAP7_75t_L g4346 ( 
.A(n_4219),
.B(n_230),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4233),
.Y(n_4347)
);

AND2x4_ASAP7_75t_L g4348 ( 
.A(n_4206),
.B(n_232),
.Y(n_4348)
);

AND2x4_ASAP7_75t_L g4349 ( 
.A(n_4206),
.B(n_233),
.Y(n_4349)
);

INVxp67_ASAP7_75t_L g4350 ( 
.A(n_4183),
.Y(n_4350)
);

NAND2xp33_ASAP7_75t_R g4351 ( 
.A(n_4210),
.B(n_233),
.Y(n_4351)
);

NOR2x1_ASAP7_75t_L g4352 ( 
.A(n_4191),
.B(n_235),
.Y(n_4352)
);

NOR2xp33_ASAP7_75t_R g4353 ( 
.A(n_4179),
.B(n_235),
.Y(n_4353)
);

CKINVDCx5p33_ASAP7_75t_R g4354 ( 
.A(n_4155),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_4221),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_L g4356 ( 
.A(n_4161),
.B(n_236),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_4172),
.B(n_236),
.Y(n_4357)
);

NOR2xp33_ASAP7_75t_R g4358 ( 
.A(n_4153),
.B(n_237),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_4152),
.B(n_237),
.Y(n_4359)
);

NAND2xp33_ASAP7_75t_R g4360 ( 
.A(n_4188),
.B(n_4215),
.Y(n_4360)
);

NAND2xp33_ASAP7_75t_R g4361 ( 
.A(n_4218),
.B(n_238),
.Y(n_4361)
);

NAND2xp33_ASAP7_75t_R g4362 ( 
.A(n_4223),
.B(n_238),
.Y(n_4362)
);

AND2x4_ASAP7_75t_L g4363 ( 
.A(n_4256),
.B(n_239),
.Y(n_4363)
);

NAND2xp33_ASAP7_75t_R g4364 ( 
.A(n_4176),
.B(n_239),
.Y(n_4364)
);

OR2x6_ASAP7_75t_L g4365 ( 
.A(n_4269),
.B(n_240),
.Y(n_4365)
);

INVxp67_ASAP7_75t_L g4366 ( 
.A(n_4196),
.Y(n_4366)
);

HB1xp67_ASAP7_75t_L g4367 ( 
.A(n_4199),
.Y(n_4367)
);

INVxp67_ASAP7_75t_L g4368 ( 
.A(n_4184),
.Y(n_4368)
);

AND2x4_ASAP7_75t_L g4369 ( 
.A(n_4241),
.B(n_241),
.Y(n_4369)
);

AND2x4_ASAP7_75t_L g4370 ( 
.A(n_4272),
.B(n_241),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_4299),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4278),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4313),
.B(n_4158),
.Y(n_4373)
);

BUFx3_ASAP7_75t_L g4374 ( 
.A(n_4276),
.Y(n_4374)
);

AND2x2_ASAP7_75t_L g4375 ( 
.A(n_4350),
.B(n_4201),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4280),
.Y(n_4376)
);

HB1xp67_ASAP7_75t_L g4377 ( 
.A(n_4367),
.Y(n_4377)
);

AOI22xp33_ASAP7_75t_L g4378 ( 
.A1(n_4352),
.A2(n_4227),
.B1(n_4265),
.B2(n_4234),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4294),
.Y(n_4379)
);

HB1xp67_ASAP7_75t_L g4380 ( 
.A(n_4289),
.Y(n_4380)
);

AND2x2_ASAP7_75t_L g4381 ( 
.A(n_4321),
.B(n_4166),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4298),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_4299),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4320),
.Y(n_4384)
);

INVx2_ASAP7_75t_SL g4385 ( 
.A(n_4326),
.Y(n_4385)
);

INVxp67_ASAP7_75t_L g4386 ( 
.A(n_4351),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4333),
.Y(n_4387)
);

AND2x2_ASAP7_75t_L g4388 ( 
.A(n_4336),
.B(n_4198),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_4315),
.B(n_4185),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_4347),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4355),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4370),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4315),
.B(n_4185),
.Y(n_4393)
);

BUFx2_ASAP7_75t_SL g4394 ( 
.A(n_4288),
.Y(n_4394)
);

INVx2_ASAP7_75t_L g4395 ( 
.A(n_4339),
.Y(n_4395)
);

OR2x2_ASAP7_75t_L g4396 ( 
.A(n_4318),
.B(n_4181),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4370),
.Y(n_4397)
);

INVx2_ASAP7_75t_L g4398 ( 
.A(n_4339),
.Y(n_4398)
);

OR2x2_ASAP7_75t_L g4399 ( 
.A(n_4368),
.B(n_4272),
.Y(n_4399)
);

HB1xp67_ASAP7_75t_L g4400 ( 
.A(n_4290),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4275),
.Y(n_4401)
);

INVx2_ASAP7_75t_L g4402 ( 
.A(n_4348),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_4281),
.B(n_4272),
.Y(n_4403)
);

INVx2_ASAP7_75t_L g4404 ( 
.A(n_4348),
.Y(n_4404)
);

AND2x2_ASAP7_75t_L g4405 ( 
.A(n_4281),
.B(n_4151),
.Y(n_4405)
);

AND2x2_ASAP7_75t_L g4406 ( 
.A(n_4277),
.B(n_4171),
.Y(n_4406)
);

NAND2x1_ASAP7_75t_L g4407 ( 
.A(n_4291),
.B(n_4190),
.Y(n_4407)
);

NOR2xp33_ASAP7_75t_L g4408 ( 
.A(n_4310),
.B(n_4244),
.Y(n_4408)
);

AND2x2_ASAP7_75t_L g4409 ( 
.A(n_4292),
.B(n_4211),
.Y(n_4409)
);

OR2x2_ASAP7_75t_L g4410 ( 
.A(n_4316),
.B(n_4211),
.Y(n_4410)
);

AND2x2_ASAP7_75t_L g4411 ( 
.A(n_4291),
.B(n_4285),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4346),
.Y(n_4412)
);

INVx2_ASAP7_75t_SL g4413 ( 
.A(n_4326),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4349),
.Y(n_4414)
);

HB1xp67_ASAP7_75t_L g4415 ( 
.A(n_4279),
.Y(n_4415)
);

OR2x2_ASAP7_75t_L g4416 ( 
.A(n_4322),
.B(n_4177),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_4349),
.Y(n_4417)
);

HB1xp67_ASAP7_75t_L g4418 ( 
.A(n_4325),
.Y(n_4418)
);

AND2x4_ASAP7_75t_L g4419 ( 
.A(n_4329),
.B(n_4203),
.Y(n_4419)
);

INVx2_ASAP7_75t_L g4420 ( 
.A(n_4363),
.Y(n_4420)
);

BUFx6f_ASAP7_75t_L g4421 ( 
.A(n_4359),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4331),
.B(n_4269),
.Y(n_4422)
);

AND2x2_ASAP7_75t_L g4423 ( 
.A(n_4300),
.B(n_4154),
.Y(n_4423)
);

OR2x2_ASAP7_75t_L g4424 ( 
.A(n_4337),
.B(n_4187),
.Y(n_4424)
);

HB1xp67_ASAP7_75t_L g4425 ( 
.A(n_4360),
.Y(n_4425)
);

AND2x2_ASAP7_75t_L g4426 ( 
.A(n_4302),
.B(n_4190),
.Y(n_4426)
);

HB1xp67_ASAP7_75t_L g4427 ( 
.A(n_4332),
.Y(n_4427)
);

AND2x2_ASAP7_75t_L g4428 ( 
.A(n_4303),
.B(n_4186),
.Y(n_4428)
);

BUFx2_ASAP7_75t_L g4429 ( 
.A(n_4284),
.Y(n_4429)
);

AND2x2_ASAP7_75t_L g4430 ( 
.A(n_4328),
.B(n_4186),
.Y(n_4430)
);

INVx2_ASAP7_75t_L g4431 ( 
.A(n_4363),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4283),
.B(n_4170),
.Y(n_4432)
);

OR2x2_ASAP7_75t_L g4433 ( 
.A(n_4305),
.B(n_4330),
.Y(n_4433)
);

INVx2_ASAP7_75t_L g4434 ( 
.A(n_4369),
.Y(n_4434)
);

OR2x2_ASAP7_75t_L g4435 ( 
.A(n_4345),
.B(n_4192),
.Y(n_4435)
);

HB1xp67_ASAP7_75t_L g4436 ( 
.A(n_4361),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_4369),
.Y(n_4437)
);

INVx2_ASAP7_75t_L g4438 ( 
.A(n_4334),
.Y(n_4438)
);

AND2x2_ASAP7_75t_L g4439 ( 
.A(n_4342),
.B(n_4208),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_4334),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_4307),
.B(n_4202),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_4427),
.B(n_4312),
.Y(n_4442)
);

NAND3xp33_ASAP7_75t_L g4443 ( 
.A(n_4425),
.B(n_4362),
.C(n_4296),
.Y(n_4443)
);

NAND3xp33_ASAP7_75t_L g4444 ( 
.A(n_4425),
.B(n_4373),
.C(n_4380),
.Y(n_4444)
);

AND2x4_ASAP7_75t_L g4445 ( 
.A(n_4385),
.B(n_4317),
.Y(n_4445)
);

NAND4xp25_ASAP7_75t_L g4446 ( 
.A(n_4373),
.B(n_4306),
.C(n_4327),
.D(n_4301),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4427),
.B(n_4295),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_L g4448 ( 
.A(n_4436),
.B(n_4344),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_4429),
.B(n_4286),
.Y(n_4449)
);

AND2x2_ASAP7_75t_L g4450 ( 
.A(n_4429),
.B(n_4297),
.Y(n_4450)
);

AND2x2_ASAP7_75t_L g4451 ( 
.A(n_4411),
.B(n_4366),
.Y(n_4451)
);

OAI22xp5_ASAP7_75t_L g4452 ( 
.A1(n_4415),
.A2(n_4354),
.B1(n_4304),
.B2(n_4365),
.Y(n_4452)
);

OAI21xp33_ASAP7_75t_L g4453 ( 
.A1(n_4400),
.A2(n_4358),
.B(n_4353),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_4436),
.B(n_4338),
.Y(n_4454)
);

AND2x2_ASAP7_75t_L g4455 ( 
.A(n_4411),
.B(n_4308),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_SL g4456 ( 
.A(n_4386),
.B(n_4309),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_4386),
.B(n_4438),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_SL g4458 ( 
.A(n_4380),
.B(n_4400),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_4438),
.B(n_4338),
.Y(n_4459)
);

AND2x2_ASAP7_75t_L g4460 ( 
.A(n_4411),
.B(n_4374),
.Y(n_4460)
);

NAND4xp25_ASAP7_75t_L g4461 ( 
.A(n_4378),
.B(n_4364),
.C(n_4228),
.D(n_4324),
.Y(n_4461)
);

NAND2xp33_ASAP7_75t_SL g4462 ( 
.A(n_4415),
.B(n_4311),
.Y(n_4462)
);

NOR2xp33_ASAP7_75t_L g4463 ( 
.A(n_4374),
.B(n_4314),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_4438),
.B(n_4440),
.Y(n_4464)
);

NAND3xp33_ASAP7_75t_L g4465 ( 
.A(n_4421),
.B(n_4433),
.C(n_4424),
.Y(n_4465)
);

OAI21xp5_ASAP7_75t_SL g4466 ( 
.A1(n_4421),
.A2(n_4335),
.B(n_4341),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4440),
.B(n_4319),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_L g4468 ( 
.A(n_4440),
.B(n_4274),
.Y(n_4468)
);

AND2x2_ASAP7_75t_L g4469 ( 
.A(n_4374),
.B(n_4308),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_4395),
.B(n_4282),
.Y(n_4470)
);

NOR3xp33_ASAP7_75t_SL g4471 ( 
.A(n_4401),
.B(n_4220),
.C(n_4216),
.Y(n_4471)
);

AOI221xp5_ASAP7_75t_L g4472 ( 
.A1(n_4421),
.A2(n_4343),
.B1(n_4238),
.B2(n_4323),
.C(n_4273),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_L g4473 ( 
.A(n_4395),
.B(n_4356),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_4395),
.B(n_4357),
.Y(n_4474)
);

AOI22xp33_ASAP7_75t_L g4475 ( 
.A1(n_4421),
.A2(n_4365),
.B1(n_4230),
.B2(n_4262),
.Y(n_4475)
);

NAND4xp25_ASAP7_75t_L g4476 ( 
.A(n_4433),
.B(n_4257),
.C(n_4340),
.D(n_4249),
.Y(n_4476)
);

NAND3xp33_ASAP7_75t_L g4477 ( 
.A(n_4421),
.B(n_4226),
.C(n_4159),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_4398),
.B(n_4287),
.Y(n_4478)
);

AOI21xp5_ASAP7_75t_SL g4479 ( 
.A1(n_4385),
.A2(n_4413),
.B(n_4422),
.Y(n_4479)
);

OAI21xp33_ASAP7_75t_L g4480 ( 
.A1(n_4416),
.A2(n_4293),
.B(n_4169),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_L g4481 ( 
.A(n_4398),
.B(n_4231),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_4398),
.B(n_4402),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_4402),
.B(n_4242),
.Y(n_4483)
);

AND2x2_ASAP7_75t_L g4484 ( 
.A(n_4420),
.B(n_242),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_L g4485 ( 
.A(n_4402),
.B(n_242),
.Y(n_4485)
);

OAI221xp5_ASAP7_75t_L g4486 ( 
.A1(n_4421),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.C(n_249),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4457),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4482),
.Y(n_4488)
);

AND2x4_ASAP7_75t_L g4489 ( 
.A(n_4460),
.B(n_4385),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4450),
.B(n_4394),
.Y(n_4490)
);

AND2x2_ASAP7_75t_L g4491 ( 
.A(n_4449),
.B(n_4394),
.Y(n_4491)
);

AND2x2_ASAP7_75t_L g4492 ( 
.A(n_4445),
.B(n_4413),
.Y(n_4492)
);

NAND3xp33_ASAP7_75t_L g4493 ( 
.A(n_4444),
.B(n_4443),
.C(n_4465),
.Y(n_4493)
);

NAND2x1p5_ASAP7_75t_L g4494 ( 
.A(n_4456),
.B(n_4407),
.Y(n_4494)
);

HB1xp67_ASAP7_75t_L g4495 ( 
.A(n_4454),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_SL g4496 ( 
.A(n_4462),
.B(n_4420),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_L g4497 ( 
.A(n_4442),
.B(n_4421),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4464),
.Y(n_4498)
);

INVx2_ASAP7_75t_L g4499 ( 
.A(n_4458),
.Y(n_4499)
);

NOR3xp33_ASAP7_75t_SL g4500 ( 
.A(n_4462),
.B(n_4401),
.C(n_4408),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4445),
.B(n_4413),
.Y(n_4501)
);

AND2x2_ASAP7_75t_L g4502 ( 
.A(n_4455),
.B(n_4404),
.Y(n_4502)
);

AOI211xp5_ASAP7_75t_SL g4503 ( 
.A1(n_4479),
.A2(n_4453),
.B(n_4486),
.C(n_4452),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_4466),
.B(n_4420),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4469),
.B(n_4404),
.Y(n_4505)
);

AND2x4_ASAP7_75t_L g4506 ( 
.A(n_4458),
.B(n_4371),
.Y(n_4506)
);

AO21x2_ASAP7_75t_L g4507 ( 
.A1(n_4447),
.A2(n_4418),
.B(n_4375),
.Y(n_4507)
);

OAI22xp5_ASAP7_75t_SL g4508 ( 
.A1(n_4475),
.A2(n_4422),
.B1(n_4407),
.B2(n_4424),
.Y(n_4508)
);

INVx2_ASAP7_75t_L g4509 ( 
.A(n_4456),
.Y(n_4509)
);

AND2x2_ASAP7_75t_L g4510 ( 
.A(n_4451),
.B(n_4404),
.Y(n_4510)
);

OR2x2_ASAP7_75t_L g4511 ( 
.A(n_4478),
.B(n_4377),
.Y(n_4511)
);

INVx1_ASAP7_75t_L g4512 ( 
.A(n_4484),
.Y(n_4512)
);

AND2x2_ASAP7_75t_L g4513 ( 
.A(n_4463),
.B(n_4417),
.Y(n_4513)
);

AND2x2_ASAP7_75t_L g4514 ( 
.A(n_4463),
.B(n_4417),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_4475),
.B(n_4377),
.Y(n_4515)
);

NAND4xp25_ASAP7_75t_L g4516 ( 
.A(n_4503),
.B(n_4446),
.C(n_4448),
.D(n_4461),
.Y(n_4516)
);

HB1xp67_ASAP7_75t_L g4517 ( 
.A(n_4506),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4490),
.B(n_4417),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4506),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4513),
.B(n_4431),
.Y(n_4520)
);

AND2x2_ASAP7_75t_L g4521 ( 
.A(n_4490),
.B(n_4432),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_4491),
.B(n_4432),
.Y(n_4522)
);

AND2x2_ASAP7_75t_L g4523 ( 
.A(n_4491),
.B(n_4432),
.Y(n_4523)
);

OR2x2_ASAP7_75t_L g4524 ( 
.A(n_4499),
.B(n_4470),
.Y(n_4524)
);

AND2x2_ASAP7_75t_L g4525 ( 
.A(n_4492),
.B(n_4431),
.Y(n_4525)
);

INVx4_ASAP7_75t_L g4526 ( 
.A(n_4489),
.Y(n_4526)
);

AND2x2_ASAP7_75t_L g4527 ( 
.A(n_4492),
.B(n_4431),
.Y(n_4527)
);

AND2x2_ASAP7_75t_L g4528 ( 
.A(n_4501),
.B(n_4434),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_4513),
.B(n_4414),
.Y(n_4529)
);

INVx2_ASAP7_75t_L g4530 ( 
.A(n_4506),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_4514),
.B(n_4414),
.Y(n_4531)
);

NAND5xp2_ASAP7_75t_L g4532 ( 
.A(n_4503),
.B(n_4472),
.C(n_4480),
.D(n_4468),
.E(n_4471),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_4501),
.B(n_4434),
.Y(n_4533)
);

OR2x2_ASAP7_75t_L g4534 ( 
.A(n_4504),
.B(n_4467),
.Y(n_4534)
);

NAND2xp5_ASAP7_75t_L g4535 ( 
.A(n_4514),
.B(n_4434),
.Y(n_4535)
);

HB1xp67_ASAP7_75t_L g4536 ( 
.A(n_4506),
.Y(n_4536)
);

AND2x4_ASAP7_75t_L g4537 ( 
.A(n_4489),
.B(n_4371),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4517),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_4526),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4536),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4530),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4530),
.Y(n_4542)
);

INVx1_ASAP7_75t_SL g4543 ( 
.A(n_4522),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4519),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_L g4545 ( 
.A(n_4522),
.B(n_4505),
.Y(n_4545)
);

OR2x2_ASAP7_75t_L g4546 ( 
.A(n_4516),
.B(n_4499),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_4523),
.B(n_4489),
.Y(n_4547)
);

OR2x2_ASAP7_75t_L g4548 ( 
.A(n_4520),
.B(n_4509),
.Y(n_4548)
);

AND2x2_ASAP7_75t_L g4549 ( 
.A(n_4523),
.B(n_4489),
.Y(n_4549)
);

OAI21xp5_ASAP7_75t_SL g4550 ( 
.A1(n_4521),
.A2(n_4493),
.B(n_4515),
.Y(n_4550)
);

AOI321xp33_ASAP7_75t_L g4551 ( 
.A1(n_4521),
.A2(n_4515),
.A3(n_4496),
.B1(n_4509),
.B2(n_4499),
.C(n_4497),
.Y(n_4551)
);

CKINVDCx16_ASAP7_75t_R g4552 ( 
.A(n_4547),
.Y(n_4552)
);

AO221x2_ASAP7_75t_L g4553 ( 
.A1(n_4550),
.A2(n_4493),
.B1(n_4509),
.B2(n_4508),
.C(n_4512),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_4547),
.B(n_4525),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_4549),
.B(n_4525),
.Y(n_4555)
);

AO221x2_ASAP7_75t_L g4556 ( 
.A1(n_4545),
.A2(n_4508),
.B1(n_4512),
.B2(n_4529),
.C(n_4531),
.Y(n_4556)
);

NOR2xp33_ASAP7_75t_R g4557 ( 
.A(n_4543),
.B(n_4549),
.Y(n_4557)
);

CKINVDCx5p33_ASAP7_75t_R g4558 ( 
.A(n_4546),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4538),
.B(n_4527),
.Y(n_4559)
);

INVxp33_ASAP7_75t_SL g4560 ( 
.A(n_4546),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4552),
.B(n_4502),
.Y(n_4561)
);

OR2x2_ASAP7_75t_L g4562 ( 
.A(n_4554),
.B(n_4535),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4555),
.B(n_4502),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4557),
.B(n_4518),
.Y(n_4564)
);

OAI211xp5_ASAP7_75t_L g4565 ( 
.A1(n_4558),
.A2(n_4551),
.B(n_4500),
.C(n_4540),
.Y(n_4565)
);

BUFx3_ASAP7_75t_L g4566 ( 
.A(n_4559),
.Y(n_4566)
);

OAI22xp33_ASAP7_75t_L g4567 ( 
.A1(n_4560),
.A2(n_4494),
.B1(n_4476),
.B2(n_4435),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_4553),
.B(n_4527),
.Y(n_4568)
);

AND2x4_ASAP7_75t_SL g4569 ( 
.A(n_4556),
.B(n_4505),
.Y(n_4569)
);

OR2x2_ASAP7_75t_L g4570 ( 
.A(n_4552),
.B(n_4497),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_4552),
.Y(n_4571)
);

INVxp67_ASAP7_75t_L g4572 ( 
.A(n_4554),
.Y(n_4572)
);

AOI222xp33_ASAP7_75t_L g4573 ( 
.A1(n_4565),
.A2(n_4487),
.B1(n_4495),
.B2(n_4498),
.C1(n_4488),
.C2(n_4518),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_4561),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4570),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4564),
.Y(n_4576)
);

INVx2_ASAP7_75t_SL g4577 ( 
.A(n_4571),
.Y(n_4577)
);

NAND2x1_ASAP7_75t_L g4578 ( 
.A(n_4563),
.B(n_4526),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4562),
.Y(n_4579)
);

INVx3_ASAP7_75t_L g4580 ( 
.A(n_4566),
.Y(n_4580)
);

NAND2xp5_ASAP7_75t_L g4581 ( 
.A(n_4569),
.B(n_4528),
.Y(n_4581)
);

AND2x2_ASAP7_75t_L g4582 ( 
.A(n_4574),
.B(n_4528),
.Y(n_4582)
);

OAI21xp5_ASAP7_75t_L g4583 ( 
.A1(n_4581),
.A2(n_4565),
.B(n_4568),
.Y(n_4583)
);

AOI21xp33_ASAP7_75t_L g4584 ( 
.A1(n_4578),
.A2(n_4567),
.B(n_4507),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4575),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_4577),
.B(n_4533),
.Y(n_4586)
);

A2O1A1Ixp33_ASAP7_75t_L g4587 ( 
.A1(n_4578),
.A2(n_4568),
.B(n_4524),
.C(n_4471),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4576),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4573),
.B(n_4533),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4582),
.Y(n_4590)
);

AOI22xp5_ASAP7_75t_L g4591 ( 
.A1(n_4588),
.A2(n_4572),
.B1(n_4580),
.B2(n_4507),
.Y(n_4591)
);

O2A1O1Ixp33_ASAP7_75t_L g4592 ( 
.A1(n_4587),
.A2(n_4539),
.B(n_4532),
.C(n_4541),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4586),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4585),
.Y(n_4594)
);

AOI22xp5_ASAP7_75t_L g4595 ( 
.A1(n_4589),
.A2(n_4507),
.B1(n_4526),
.B2(n_4510),
.Y(n_4595)
);

AOI22xp5_ASAP7_75t_L g4596 ( 
.A1(n_4583),
.A2(n_4507),
.B1(n_4510),
.B2(n_4537),
.Y(n_4596)
);

AOI221xp5_ASAP7_75t_L g4597 ( 
.A1(n_4592),
.A2(n_4584),
.B1(n_4544),
.B2(n_4542),
.C(n_4539),
.Y(n_4597)
);

AND2x2_ASAP7_75t_L g4598 ( 
.A(n_4590),
.B(n_4579),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4596),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_4593),
.B(n_4548),
.Y(n_4600)
);

NAND3xp33_ASAP7_75t_L g4601 ( 
.A(n_4595),
.B(n_4487),
.C(n_4524),
.Y(n_4601)
);

AOI222xp33_ASAP7_75t_L g4602 ( 
.A1(n_4594),
.A2(n_4488),
.B1(n_4498),
.B2(n_4537),
.C1(n_4418),
.C2(n_4477),
.Y(n_4602)
);

XOR2xp5_ASAP7_75t_L g4603 ( 
.A(n_4591),
.B(n_4534),
.Y(n_4603)
);

O2A1O1Ixp33_ASAP7_75t_L g4604 ( 
.A1(n_4592),
.A2(n_4494),
.B(n_4511),
.C(n_4485),
.Y(n_4604)
);

AOI21xp5_ASAP7_75t_L g4605 ( 
.A1(n_4592),
.A2(n_4511),
.B(n_4537),
.Y(n_4605)
);

NAND2xp5_ASAP7_75t_L g4606 ( 
.A(n_4595),
.B(n_4459),
.Y(n_4606)
);

INVxp67_ASAP7_75t_L g4607 ( 
.A(n_4590),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4595),
.B(n_4392),
.Y(n_4608)
);

INVx1_ASAP7_75t_SL g4609 ( 
.A(n_4590),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_4595),
.B(n_4392),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4592),
.Y(n_4611)
);

HB1xp67_ASAP7_75t_L g4612 ( 
.A(n_4600),
.Y(n_4612)
);

INVx2_ASAP7_75t_L g4613 ( 
.A(n_4598),
.Y(n_4613)
);

CKINVDCx5p33_ASAP7_75t_R g4614 ( 
.A(n_4609),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4608),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_4610),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4606),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_4604),
.Y(n_4618)
);

INVx2_ASAP7_75t_L g4619 ( 
.A(n_4607),
.Y(n_4619)
);

INVx1_ASAP7_75t_SL g4620 ( 
.A(n_4605),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4601),
.Y(n_4621)
);

INVx2_ASAP7_75t_L g4622 ( 
.A(n_4611),
.Y(n_4622)
);

INVx2_ASAP7_75t_L g4623 ( 
.A(n_4599),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4603),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4602),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4597),
.Y(n_4626)
);

INVxp67_ASAP7_75t_SL g4627 ( 
.A(n_4600),
.Y(n_4627)
);

INVx1_ASAP7_75t_SL g4628 ( 
.A(n_4600),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4598),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4602),
.B(n_4473),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4598),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4598),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4598),
.Y(n_4633)
);

INVx1_ASAP7_75t_SL g4634 ( 
.A(n_4600),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4598),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4598),
.Y(n_4636)
);

A2O1A1Ixp33_ASAP7_75t_L g4637 ( 
.A1(n_4627),
.A2(n_4383),
.B(n_4371),
.C(n_4375),
.Y(n_4637)
);

OAI21xp33_ASAP7_75t_L g4638 ( 
.A1(n_4614),
.A2(n_4494),
.B(n_4474),
.Y(n_4638)
);

NOR2x1_ASAP7_75t_L g4639 ( 
.A(n_4613),
.B(n_4416),
.Y(n_4639)
);

NAND5xp2_ASAP7_75t_L g4640 ( 
.A(n_4624),
.B(n_4375),
.C(n_4388),
.D(n_4397),
.E(n_4481),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4612),
.Y(n_4641)
);

AOI211xp5_ASAP7_75t_L g4642 ( 
.A1(n_4620),
.A2(n_4383),
.B(n_4397),
.C(n_4483),
.Y(n_4642)
);

AOI21xp33_ASAP7_75t_L g4643 ( 
.A1(n_4627),
.A2(n_4383),
.B(n_4441),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4612),
.B(n_4437),
.Y(n_4644)
);

OAI21xp33_ASAP7_75t_L g4645 ( 
.A1(n_4628),
.A2(n_4441),
.B(n_4388),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4613),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4629),
.Y(n_4647)
);

AOI221xp5_ASAP7_75t_L g4648 ( 
.A1(n_4625),
.A2(n_4412),
.B1(n_4441),
.B2(n_4437),
.C(n_4428),
.Y(n_4648)
);

OAI22xp33_ASAP7_75t_SL g4649 ( 
.A1(n_4630),
.A2(n_4435),
.B1(n_4410),
.B2(n_4399),
.Y(n_4649)
);

AOI211xp5_ASAP7_75t_L g4650 ( 
.A1(n_4634),
.A2(n_4435),
.B(n_4428),
.C(n_4430),
.Y(n_4650)
);

NOR2xp33_ASAP7_75t_L g4651 ( 
.A(n_4629),
.B(n_4412),
.Y(n_4651)
);

XNOR2x1_ASAP7_75t_L g4652 ( 
.A(n_4622),
.B(n_4388),
.Y(n_4652)
);

OAI21xp5_ASAP7_75t_L g4653 ( 
.A1(n_4631),
.A2(n_4437),
.B(n_4430),
.Y(n_4653)
);

INVxp67_ASAP7_75t_L g4654 ( 
.A(n_4632),
.Y(n_4654)
);

AOI322xp5_ASAP7_75t_L g4655 ( 
.A1(n_4636),
.A2(n_4430),
.A3(n_4428),
.B1(n_4426),
.B2(n_4403),
.C1(n_4423),
.C2(n_4405),
.Y(n_4655)
);

AOI21xp5_ASAP7_75t_L g4656 ( 
.A1(n_4633),
.A2(n_4399),
.B(n_4410),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4635),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4618),
.Y(n_4658)
);

XOR2x2_ASAP7_75t_L g4659 ( 
.A(n_4626),
.B(n_4396),
.Y(n_4659)
);

OAI221xp5_ASAP7_75t_L g4660 ( 
.A1(n_4621),
.A2(n_4396),
.B1(n_4372),
.B2(n_4390),
.C(n_4376),
.Y(n_4660)
);

AOI22xp5_ASAP7_75t_L g4661 ( 
.A1(n_4623),
.A2(n_4426),
.B1(n_4423),
.B2(n_4405),
.Y(n_4661)
);

AOI21xp5_ASAP7_75t_SL g4662 ( 
.A1(n_4623),
.A2(n_4616),
.B(n_4619),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4616),
.Y(n_4663)
);

AOI22xp5_ASAP7_75t_L g4664 ( 
.A1(n_4617),
.A2(n_4426),
.B1(n_4423),
.B2(n_4405),
.Y(n_4664)
);

OAI21xp5_ASAP7_75t_L g4665 ( 
.A1(n_4639),
.A2(n_4615),
.B(n_4403),
.Y(n_4665)
);

NAND4xp75_ASAP7_75t_L g4666 ( 
.A(n_4641),
.B(n_4403),
.C(n_4389),
.D(n_4393),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_4644),
.Y(n_4667)
);

NOR4xp25_ASAP7_75t_L g4668 ( 
.A(n_4646),
.B(n_4387),
.C(n_4376),
.D(n_4379),
.Y(n_4668)
);

NAND2xp33_ASAP7_75t_R g4669 ( 
.A(n_4647),
.B(n_246),
.Y(n_4669)
);

OAI21xp5_ASAP7_75t_L g4670 ( 
.A1(n_4643),
.A2(n_4645),
.B(n_4652),
.Y(n_4670)
);

AOI221xp5_ASAP7_75t_L g4671 ( 
.A1(n_4649),
.A2(n_4372),
.B1(n_4379),
.B2(n_4382),
.C(n_4384),
.Y(n_4671)
);

OAI221xp5_ASAP7_75t_L g4672 ( 
.A1(n_4638),
.A2(n_4390),
.B1(n_4382),
.B2(n_4384),
.C(n_4387),
.Y(n_4672)
);

AOI211xp5_ASAP7_75t_L g4673 ( 
.A1(n_4662),
.A2(n_4391),
.B(n_4389),
.C(n_4393),
.Y(n_4673)
);

AOI322xp5_ASAP7_75t_L g4674 ( 
.A1(n_4648),
.A2(n_4419),
.A3(n_4406),
.B1(n_4393),
.B2(n_4389),
.C1(n_4391),
.C2(n_4439),
.Y(n_4674)
);

OAI211xp5_ASAP7_75t_SL g4675 ( 
.A1(n_4654),
.A2(n_247),
.B(n_250),
.C(n_251),
.Y(n_4675)
);

NAND4xp25_ASAP7_75t_L g4676 ( 
.A(n_4642),
.B(n_4406),
.C(n_4439),
.D(n_4419),
.Y(n_4676)
);

NAND4xp25_ASAP7_75t_L g4677 ( 
.A(n_4640),
.B(n_4406),
.C(n_4439),
.D(n_4419),
.Y(n_4677)
);

AOI222xp33_ASAP7_75t_L g4678 ( 
.A1(n_4653),
.A2(n_4419),
.B1(n_4381),
.B2(n_4409),
.C1(n_257),
.C2(n_258),
.Y(n_4678)
);

NAND3xp33_ASAP7_75t_L g4679 ( 
.A(n_4657),
.B(n_4419),
.C(n_4381),
.Y(n_4679)
);

NAND2xp5_ASAP7_75t_L g4680 ( 
.A(n_4661),
.B(n_4381),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4659),
.Y(n_4681)
);

AND2x2_ASAP7_75t_L g4682 ( 
.A(n_4664),
.B(n_4409),
.Y(n_4682)
);

AOI211xp5_ASAP7_75t_SL g4683 ( 
.A1(n_4658),
.A2(n_4409),
.B(n_254),
.C(n_255),
.Y(n_4683)
);

O2A1O1Ixp33_ASAP7_75t_L g4684 ( 
.A1(n_4663),
.A2(n_252),
.B(n_258),
.C(n_259),
.Y(n_4684)
);

OAI211xp5_ASAP7_75t_SL g4685 ( 
.A1(n_4651),
.A2(n_260),
.B(n_261),
.C(n_262),
.Y(n_4685)
);

AOI221x1_ASAP7_75t_L g4686 ( 
.A1(n_4656),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.C(n_264),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_SL g4687 ( 
.A(n_4637),
.B(n_264),
.Y(n_4687)
);

INVx2_ASAP7_75t_SL g4688 ( 
.A(n_4650),
.Y(n_4688)
);

AOI21xp33_ASAP7_75t_SL g4689 ( 
.A1(n_4660),
.A2(n_265),
.B(n_266),
.Y(n_4689)
);

AOI221xp5_ASAP7_75t_L g4690 ( 
.A1(n_4689),
.A2(n_4655),
.B1(n_267),
.B2(n_268),
.C(n_269),
.Y(n_4690)
);

AOI22xp5_ASAP7_75t_L g4691 ( 
.A1(n_4688),
.A2(n_266),
.B1(n_267),
.B2(n_270),
.Y(n_4691)
);

AOI221xp5_ASAP7_75t_L g4692 ( 
.A1(n_4668),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.C(n_277),
.Y(n_4692)
);

NOR3xp33_ASAP7_75t_L g4693 ( 
.A(n_4670),
.B(n_273),
.C(n_274),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4680),
.Y(n_4694)
);

OAI32xp33_ASAP7_75t_L g4695 ( 
.A1(n_4669),
.A2(n_277),
.A3(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_4695)
);

BUFx6f_ASAP7_75t_L g4696 ( 
.A(n_4667),
.Y(n_4696)
);

OAI22xp5_ASAP7_75t_L g4697 ( 
.A1(n_4679),
.A2(n_4673),
.B1(n_4666),
.B2(n_4681),
.Y(n_4697)
);

OAI21xp33_ASAP7_75t_L g4698 ( 
.A1(n_4677),
.A2(n_280),
.B(n_282),
.Y(n_4698)
);

AOI211xp5_ASAP7_75t_L g4699 ( 
.A1(n_4665),
.A2(n_283),
.B(n_284),
.C(n_285),
.Y(n_4699)
);

NOR2x1_ASAP7_75t_L g4700 ( 
.A(n_4675),
.B(n_283),
.Y(n_4700)
);

AOI221xp5_ASAP7_75t_L g4701 ( 
.A1(n_4682),
.A2(n_284),
.B1(n_285),
.B2(n_287),
.C(n_289),
.Y(n_4701)
);

NAND3xp33_ASAP7_75t_L g4702 ( 
.A(n_4683),
.B(n_291),
.C(n_292),
.Y(n_4702)
);

NAND4xp75_ASAP7_75t_L g4703 ( 
.A(n_4686),
.B(n_291),
.C(n_292),
.D(n_293),
.Y(n_4703)
);

AND4x1_ASAP7_75t_L g4704 ( 
.A(n_4684),
.B(n_294),
.C(n_295),
.D(n_297),
.Y(n_4704)
);

AOI221xp5_ASAP7_75t_L g4705 ( 
.A1(n_4687),
.A2(n_294),
.B1(n_295),
.B2(n_297),
.C(n_298),
.Y(n_4705)
);

OAI211xp5_ASAP7_75t_L g4706 ( 
.A1(n_4685),
.A2(n_299),
.B(n_300),
.C(n_301),
.Y(n_4706)
);

NAND3x1_ASAP7_75t_L g4707 ( 
.A(n_4671),
.B(n_299),
.C(n_302),
.Y(n_4707)
);

NOR2x1_ASAP7_75t_L g4708 ( 
.A(n_4703),
.B(n_4676),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4702),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_4707),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4704),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4692),
.B(n_4678),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4700),
.Y(n_4713)
);

INVx2_ASAP7_75t_L g4714 ( 
.A(n_4696),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_SL g4715 ( 
.A(n_4690),
.B(n_4674),
.Y(n_4715)
);

NOR2xp33_ASAP7_75t_L g4716 ( 
.A(n_4698),
.B(n_4672),
.Y(n_4716)
);

NOR2xp67_ASAP7_75t_L g4717 ( 
.A(n_4706),
.B(n_302),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4695),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4696),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4691),
.Y(n_4720)
);

INVx1_ASAP7_75t_SL g4721 ( 
.A(n_4694),
.Y(n_4721)
);

AOI22xp5_ASAP7_75t_L g4722 ( 
.A1(n_4693),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4717),
.B(n_4699),
.Y(n_4723)
);

NAND3xp33_ASAP7_75t_L g4724 ( 
.A(n_4715),
.B(n_4697),
.C(n_4701),
.Y(n_4724)
);

AOI221xp5_ASAP7_75t_L g4725 ( 
.A1(n_4721),
.A2(n_4705),
.B1(n_306),
.B2(n_307),
.C(n_310),
.Y(n_4725)
);

NOR2x1_ASAP7_75t_L g4726 ( 
.A(n_4713),
.B(n_304),
.Y(n_4726)
);

NAND2x1_ASAP7_75t_L g4727 ( 
.A(n_4711),
.B(n_307),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4708),
.Y(n_4728)
);

NOR3xp33_ASAP7_75t_L g4729 ( 
.A(n_4714),
.B(n_310),
.C(n_311),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4718),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4722),
.B(n_311),
.Y(n_4731)
);

NOR3xp33_ASAP7_75t_L g4732 ( 
.A(n_4719),
.B(n_313),
.C(n_315),
.Y(n_4732)
);

NAND4xp25_ASAP7_75t_L g4733 ( 
.A(n_4716),
.B(n_315),
.C(n_317),
.D(n_319),
.Y(n_4733)
);

OR2x2_ASAP7_75t_L g4734 ( 
.A(n_4710),
.B(n_317),
.Y(n_4734)
);

NOR2x1_ASAP7_75t_L g4735 ( 
.A(n_4709),
.B(n_319),
.Y(n_4735)
);

NOR2xp33_ASAP7_75t_R g4736 ( 
.A(n_4730),
.B(n_4720),
.Y(n_4736)
);

XNOR2xp5_ASAP7_75t_L g4737 ( 
.A(n_4724),
.B(n_4712),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_SL g4738 ( 
.A(n_4725),
.B(n_320),
.Y(n_4738)
);

NOR2xp33_ASAP7_75t_R g4739 ( 
.A(n_4728),
.B(n_320),
.Y(n_4739)
);

NOR2xp33_ASAP7_75t_R g4740 ( 
.A(n_4734),
.B(n_321),
.Y(n_4740)
);

NAND3xp33_ASAP7_75t_L g4741 ( 
.A(n_4726),
.B(n_321),
.C(n_322),
.Y(n_4741)
);

NAND3xp33_ASAP7_75t_L g4742 ( 
.A(n_4735),
.B(n_322),
.C(n_323),
.Y(n_4742)
);

NAND2x1_ASAP7_75t_SL g4743 ( 
.A(n_4727),
.B(n_323),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_SL g4744 ( 
.A(n_4729),
.B(n_326),
.Y(n_4744)
);

AND4x1_ASAP7_75t_L g4745 ( 
.A(n_4732),
.B(n_327),
.C(n_328),
.D(n_329),
.Y(n_4745)
);

A2O1A1Ixp33_ASAP7_75t_L g4746 ( 
.A1(n_4743),
.A2(n_4731),
.B(n_4723),
.C(n_4733),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4741),
.Y(n_4747)
);

NOR4xp75_ASAP7_75t_L g4748 ( 
.A(n_4738),
.B(n_329),
.C(n_330),
.D(n_331),
.Y(n_4748)
);

INVx2_ASAP7_75t_L g4749 ( 
.A(n_4737),
.Y(n_4749)
);

INVx1_ASAP7_75t_SL g4750 ( 
.A(n_4739),
.Y(n_4750)
);

NOR3xp33_ASAP7_75t_L g4751 ( 
.A(n_4744),
.B(n_330),
.C(n_331),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_L g4752 ( 
.A(n_4745),
.B(n_332),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4752),
.Y(n_4753)
);

CKINVDCx5p33_ASAP7_75t_R g4754 ( 
.A(n_4750),
.Y(n_4754)
);

INVx1_ASAP7_75t_SL g4755 ( 
.A(n_4748),
.Y(n_4755)
);

OR2x2_ASAP7_75t_L g4756 ( 
.A(n_4755),
.B(n_4742),
.Y(n_4756)
);

OAI21xp5_ASAP7_75t_L g4757 ( 
.A1(n_4753),
.A2(n_4746),
.B(n_4749),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4756),
.Y(n_4758)
);

HB1xp67_ASAP7_75t_L g4759 ( 
.A(n_4757),
.Y(n_4759)
);

OAI22xp5_ASAP7_75t_L g4760 ( 
.A1(n_4759),
.A2(n_4754),
.B1(n_4747),
.B2(n_4751),
.Y(n_4760)
);

AND2x4_ASAP7_75t_L g4761 ( 
.A(n_4758),
.B(n_4736),
.Y(n_4761)
);

INVx2_ASAP7_75t_L g4762 ( 
.A(n_4758),
.Y(n_4762)
);

AOI31xp33_ASAP7_75t_L g4763 ( 
.A1(n_4760),
.A2(n_4740),
.A3(n_333),
.B(n_334),
.Y(n_4763)
);

AOI22xp33_ASAP7_75t_L g4764 ( 
.A1(n_4762),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_4764)
);

AOI22xp33_ASAP7_75t_L g4765 ( 
.A1(n_4761),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_4765)
);

AOI31xp33_ASAP7_75t_L g4766 ( 
.A1(n_4760),
.A2(n_336),
.A3(n_338),
.B(n_339),
.Y(n_4766)
);

HB1xp67_ASAP7_75t_L g4767 ( 
.A(n_4763),
.Y(n_4767)
);

INVx1_ASAP7_75t_SL g4768 ( 
.A(n_4766),
.Y(n_4768)
);

AOI222xp33_ASAP7_75t_SL g4769 ( 
.A1(n_4765),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.C1(n_341),
.C2(n_342),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4764),
.Y(n_4770)
);

AOI21xp5_ASAP7_75t_L g4771 ( 
.A1(n_4763),
.A2(n_340),
.B(n_341),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_SL g4772 ( 
.A(n_4771),
.B(n_344),
.Y(n_4772)
);

AOI21xp33_ASAP7_75t_SL g4773 ( 
.A1(n_4770),
.A2(n_345),
.B(n_346),
.Y(n_4773)
);

AOI21xp5_ASAP7_75t_L g4774 ( 
.A1(n_4768),
.A2(n_4767),
.B(n_4769),
.Y(n_4774)
);

AOI21xp5_ASAP7_75t_L g4775 ( 
.A1(n_4768),
.A2(n_346),
.B(n_348),
.Y(n_4775)
);

OAI21x1_ASAP7_75t_SL g4776 ( 
.A1(n_4771),
.A2(n_348),
.B(n_349),
.Y(n_4776)
);

OA22x2_ASAP7_75t_L g4777 ( 
.A1(n_4768),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_4771),
.B(n_350),
.Y(n_4778)
);

AOI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_4768),
.A2(n_352),
.B(n_353),
.Y(n_4779)
);

AOI21xp5_ASAP7_75t_L g4780 ( 
.A1(n_4768),
.A2(n_355),
.B(n_357),
.Y(n_4780)
);

AOI222xp33_ASAP7_75t_L g4781 ( 
.A1(n_4768),
.A2(n_355),
.B1(n_359),
.B2(n_360),
.C1(n_362),
.C2(n_363),
.Y(n_4781)
);

AOI22xp33_ASAP7_75t_R g4782 ( 
.A1(n_4776),
.A2(n_359),
.B1(n_362),
.B2(n_364),
.Y(n_4782)
);

INVxp67_ASAP7_75t_L g4783 ( 
.A(n_4778),
.Y(n_4783)
);

AOI22xp5_ASAP7_75t_L g4784 ( 
.A1(n_4772),
.A2(n_4774),
.B1(n_4780),
.B2(n_4779),
.Y(n_4784)
);

AOI222xp33_ASAP7_75t_L g4785 ( 
.A1(n_4775),
.A2(n_365),
.B1(n_366),
.B2(n_368),
.C1(n_369),
.C2(n_370),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4777),
.Y(n_4786)
);

OR2x6_ASAP7_75t_L g4787 ( 
.A(n_4773),
.B(n_1641),
.Y(n_4787)
);

AOI31xp33_ASAP7_75t_L g4788 ( 
.A1(n_4781),
.A2(n_368),
.A3(n_369),
.B(n_370),
.Y(n_4788)
);

AOI222xp33_ASAP7_75t_SL g4789 ( 
.A1(n_4776),
.A2(n_373),
.B1(n_374),
.B2(n_375),
.C1(n_376),
.C2(n_378),
.Y(n_4789)
);

OAI21xp5_ASAP7_75t_L g4790 ( 
.A1(n_4774),
.A2(n_373),
.B(n_374),
.Y(n_4790)
);

HB1xp67_ASAP7_75t_L g4791 ( 
.A(n_4786),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4787),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4790),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4788),
.Y(n_4794)
);

AOI21xp33_ASAP7_75t_L g4795 ( 
.A1(n_4783),
.A2(n_375),
.B(n_376),
.Y(n_4795)
);

XNOR2xp5_ASAP7_75t_L g4796 ( 
.A(n_4791),
.B(n_4784),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4794),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4793),
.Y(n_4798)
);

AOI22xp33_ASAP7_75t_L g4799 ( 
.A1(n_4792),
.A2(n_4785),
.B1(n_4782),
.B2(n_4789),
.Y(n_4799)
);

OAI221xp5_ASAP7_75t_R g4800 ( 
.A1(n_4796),
.A2(n_4795),
.B1(n_380),
.B2(n_381),
.C(n_382),
.Y(n_4800)
);

OAI221xp5_ASAP7_75t_R g4801 ( 
.A1(n_4799),
.A2(n_379),
.B1(n_380),
.B2(n_381),
.C(n_382),
.Y(n_4801)
);

OAI221xp5_ASAP7_75t_R g4802 ( 
.A1(n_4798),
.A2(n_4797),
.B1(n_384),
.B2(n_386),
.C(n_387),
.Y(n_4802)
);

OAI221xp5_ASAP7_75t_R g4803 ( 
.A1(n_4796),
.A2(n_383),
.B1(n_384),
.B2(n_386),
.C(n_389),
.Y(n_4803)
);

AOI21xp5_ASAP7_75t_L g4804 ( 
.A1(n_4800),
.A2(n_1679),
.B(n_1652),
.Y(n_4804)
);

AOI211xp5_ASAP7_75t_L g4805 ( 
.A1(n_4804),
.A2(n_4802),
.B(n_4801),
.C(n_4803),
.Y(n_4805)
);


endmodule