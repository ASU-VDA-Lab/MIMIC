module fake_jpeg_14073_n_176 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_33),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_12),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

CKINVDCx6p67_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_24),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_77),
.Y(n_82)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_78),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_25),
.B1(n_46),
.B2(n_43),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_71),
.B1(n_58),
.B2(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_26),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_89),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_94),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_55),
.Y(n_89)
);

OA22x2_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_71),
.B1(n_62),
.B2(n_64),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_69),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_70),
.Y(n_101)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_110),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_58),
.B1(n_60),
.B2(n_65),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_69),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_85),
.B1(n_89),
.B2(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_60),
.B1(n_63),
.B2(n_54),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_67),
.B1(n_59),
.B2(n_51),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_53),
.B1(n_64),
.B2(n_7),
.Y(n_130)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_114),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_54),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_0),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_113),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_116),
.B1(n_6),
.B2(n_7),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_1),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_28),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_118),
.B(n_122),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_69),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_126),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_2),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_128),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_97),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_16),
.B1(n_20),
.B2(n_22),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_64),
.C(n_53),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_133),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_4),
.B(n_6),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_108),
.B(n_11),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_4),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_8),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_99),
.B1(n_12),
.B2(n_13),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_140),
.B(n_146),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_123),
.B(n_118),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_144),
.Y(n_158)
);

INVxp33_ASAP7_75t_SL g144 ( 
.A(n_130),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_147),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_10),
.B(n_14),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_154),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_131),
.A2(n_23),
.B1(n_29),
.B2(n_31),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_47),
.B1(n_35),
.B2(n_36),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_137),
.B(n_125),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_132),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_157),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_117),
.C(n_129),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_117),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_149),
.B(n_146),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_164),
.A2(n_152),
.B1(n_150),
.B2(n_139),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_165),
.Y(n_170)
);

AOI321xp33_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_167),
.A3(n_160),
.B1(n_162),
.B2(n_163),
.C(n_164),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_143),
.B1(n_148),
.B2(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_169),
.B(n_168),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_170),
.B1(n_168),
.B2(n_161),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_161),
.B(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_34),
.C(n_37),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_38),
.Y(n_176)
);


endmodule