module fake_jpeg_31003_n_66 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_66);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_66;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_1),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_5),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_30),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_9),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_29),
.B1(n_15),
.B2(n_18),
.Y(n_34)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_31),
.B1(n_16),
.B2(n_19),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_13),
.B(n_6),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_7),
.B(n_16),
.C(n_21),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_14),
.A2(n_7),
.B1(n_15),
.B2(n_18),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_28),
.Y(n_42)
);

NOR2xp67_ASAP7_75t_R g47 ( 
.A(n_35),
.B(n_39),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_23),
.A2(n_31),
.B1(n_22),
.B2(n_26),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_23),
.B1(n_37),
.B2(n_40),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_28),
.C(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_43),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_23),
.Y(n_43)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_34),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_49),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_45),
.B(n_47),
.C(n_37),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_53),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_58),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_63),
.C(n_46),
.Y(n_64)
);

AOI221xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_56),
.B1(n_57),
.B2(n_55),
.C(n_32),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_36),
.B(n_40),
.Y(n_65)
);

INVxp33_ASAP7_75t_SL g66 ( 
.A(n_65),
.Y(n_66)
);


endmodule