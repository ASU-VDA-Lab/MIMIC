module fake_jpeg_2779_n_561 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_561);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_561;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_509;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_6),
.B(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_59),
.B(n_77),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_62),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_65),
.Y(n_135)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g202 ( 
.A(n_64),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_23),
.B(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_30),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_66),
.B(n_72),
.Y(n_150)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g127 ( 
.A(n_67),
.Y(n_127)
);

INVx11_ASAP7_75t_SL g68 ( 
.A(n_30),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_68),
.Y(n_130)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_70),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_71),
.B(n_74),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_25),
.B(n_1),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_75),
.B(n_78),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_1),
.C(n_3),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_79),
.B(n_101),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_83),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_81),
.B(n_98),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_82),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_3),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_85),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_86),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_87),
.B(n_97),
.Y(n_154)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_89),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_49),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_54),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_25),
.B(n_4),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_40),
.B(n_4),
.Y(n_106)
);

NAND2xp67_ASAP7_75t_SL g168 ( 
.A(n_106),
.B(n_32),
.Y(n_168)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_27),
.B(n_5),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_108),
.B(n_116),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_40),
.Y(n_112)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_29),
.B(n_32),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_34),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_118),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_34),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_40),
.Y(n_119)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_120),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_29),
.B(n_5),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_37),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_31),
.Y(n_125)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_33),
.B1(n_26),
.B2(n_23),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_132),
.A2(n_140),
.B1(n_166),
.B2(n_171),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_33),
.B1(n_26),
.B2(n_35),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_60),
.A2(n_42),
.B1(n_55),
.B2(n_53),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_142),
.A2(n_191),
.B1(n_198),
.B2(n_207),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_145),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_66),
.A2(n_39),
.B1(n_55),
.B2(n_53),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_149),
.A2(n_70),
.B1(n_111),
.B2(n_90),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_152),
.B(n_163),
.Y(n_243)
);

BUFx2_ASAP7_75t_R g161 ( 
.A(n_68),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_161),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_88),
.B(n_35),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_72),
.A2(n_101),
.B1(n_106),
.B2(n_97),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_168),
.B(n_192),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_125),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_170),
.B(n_172),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_79),
.A2(n_37),
.B1(n_51),
.B2(n_43),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_91),
.B(n_31),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_178),
.B(n_188),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_72),
.A2(n_39),
.B1(n_51),
.B2(n_43),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_185),
.B1(n_187),
.B2(n_193),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_76),
.A2(n_86),
.B1(n_82),
.B2(n_85),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_99),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_103),
.B(n_44),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_61),
.A2(n_41),
.B1(n_34),
.B2(n_45),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_69),
.B(n_5),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_101),
.A2(n_34),
.B1(n_48),
.B2(n_45),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_93),
.Y(n_194)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_74),
.B(n_5),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_197),
.B(n_206),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_73),
.A2(n_34),
.B1(n_48),
.B2(n_45),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_94),
.Y(n_199)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_107),
.A2(n_56),
.B1(n_48),
.B2(n_10),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_200),
.A2(n_109),
.B1(n_105),
.B2(n_11),
.Y(n_267)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_205),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_106),
.B(n_8),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_95),
.A2(n_56),
.B1(n_9),
.B2(n_10),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_191),
.A2(n_102),
.B1(n_64),
.B2(n_92),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_209),
.A2(n_278),
.B1(n_202),
.B2(n_203),
.Y(n_291)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_145),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_211),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_212),
.Y(n_299)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_215),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_120),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_216),
.B(n_221),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_217),
.Y(n_316)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_144),
.Y(n_218)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_218),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_153),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_219),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_135),
.B(n_89),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_222),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_138),
.B(n_119),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_223),
.B(n_236),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_136),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_224),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_173),
.A2(n_112),
.B(n_119),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_225),
.A2(n_176),
.B(n_182),
.Y(n_306)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_140),
.A2(n_100),
.B1(n_113),
.B2(n_110),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_230),
.A2(n_233),
.B1(n_267),
.B2(n_270),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_154),
.B(n_104),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_231),
.B(n_232),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_173),
.B(n_114),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_185),
.A2(n_115),
.B1(n_96),
.B2(n_121),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_139),
.B(n_84),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_238),
.B(n_251),
.Y(n_303)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_141),
.Y(n_239)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_239),
.Y(n_314)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_242),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_127),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_244),
.B(n_245),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_130),
.Y(n_245)
);

AO22x1_ASAP7_75t_L g246 ( 
.A1(n_150),
.A2(n_62),
.B1(n_111),
.B2(n_90),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_246),
.A2(n_208),
.B(n_156),
.Y(n_292)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_165),
.Y(n_247)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_247),
.Y(n_308)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_134),
.Y(n_248)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_249),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_136),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_250),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_147),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_127),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_252),
.B(n_255),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_196),
.Y(n_253)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_253),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_196),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_160),
.Y(n_256)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_150),
.B(n_8),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_176),
.Y(n_298)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_160),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_258),
.Y(n_293)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_169),
.Y(n_259)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_143),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_263),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_151),
.Y(n_261)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_261),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_151),
.Y(n_262)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_184),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_137),
.A2(n_122),
.B1(n_56),
.B2(n_124),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_264),
.A2(n_274),
.B1(n_208),
.B2(n_158),
.Y(n_279)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_175),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_269),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_129),
.B(n_8),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_266),
.B(n_273),
.Y(n_330)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_169),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_200),
.A2(n_131),
.B1(n_143),
.B2(n_133),
.Y(n_270)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_181),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_275),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_128),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_158),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_157),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_186),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_276),
.Y(n_296)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_204),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_189),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_159),
.B(n_10),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_279),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_213),
.A2(n_142),
.B1(n_207),
.B2(n_149),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_282),
.A2(n_305),
.B1(n_229),
.B2(n_210),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_201),
.B1(n_184),
.B2(n_195),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_287),
.A2(n_289),
.B1(n_328),
.B2(n_267),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_271),
.A2(n_195),
.B1(n_201),
.B2(n_203),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_291),
.A2(n_297),
.B1(n_323),
.B2(n_326),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_292),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_225),
.A2(n_182),
.B(n_156),
.Y(n_294)
);

OA21x2_ASAP7_75t_L g369 ( 
.A1(n_294),
.A2(n_211),
.B(n_259),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_214),
.A2(n_146),
.B1(n_202),
.B2(n_204),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_298),
.B(n_283),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_231),
.B(n_155),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_301),
.B(n_218),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_214),
.A2(n_126),
.B1(n_155),
.B2(n_128),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_306),
.Y(n_338)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_232),
.A2(n_182),
.B(n_157),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_246),
.C(n_238),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_246),
.B(n_126),
.Y(n_318)
);

XNOR2x1_ASAP7_75t_SL g354 ( 
.A(n_318),
.B(n_270),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_253),
.A2(n_189),
.B1(n_167),
.B2(n_13),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_253),
.A2(n_167),
.B1(n_12),
.B2(n_13),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_213),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_353),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_331),
.A2(n_237),
.B1(n_227),
.B2(n_222),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_335),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_312),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_336),
.B(n_337),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_312),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_280),
.Y(n_339)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_303),
.B(n_243),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_341),
.B(n_342),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_281),
.B(n_254),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_343),
.A2(n_357),
.B1(n_362),
.B2(n_370),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_309),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_356),
.Y(n_375)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_346),
.B(n_348),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_347),
.B(n_358),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_301),
.B(n_257),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_295),
.B(n_241),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_360),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_295),
.B(n_265),
.C(n_229),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_350),
.B(n_359),
.C(n_363),
.Y(n_390)
);

AOI31xp67_ASAP7_75t_L g376 ( 
.A1(n_354),
.A2(n_318),
.A3(n_292),
.B(n_304),
.Y(n_376)
);

INVx6_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_283),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_287),
.A2(n_240),
.B1(n_263),
.B2(n_224),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_283),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_294),
.B(n_217),
.C(n_212),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_307),
.B(n_268),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_210),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_289),
.A2(n_261),
.B1(n_262),
.B2(n_250),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_306),
.B(n_248),
.C(n_277),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_285),
.Y(n_364)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_365),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_321),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_366),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_304),
.A2(n_256),
.B1(n_258),
.B2(n_269),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_367),
.A2(n_369),
.B(n_220),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_317),
.B(n_234),
.C(n_272),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_372),
.C(n_308),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_328),
.A2(n_318),
.B1(n_305),
.B2(n_291),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_285),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_371),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_298),
.B(n_228),
.C(n_249),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_320),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_373),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_376),
.A2(n_397),
.B(n_401),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_338),
.A2(n_290),
.B1(n_300),
.B2(n_313),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_382),
.A2(n_389),
.B1(n_403),
.B2(n_406),
.Y(n_408)
);

AOI22x1_ASAP7_75t_SL g386 ( 
.A1(n_338),
.A2(n_300),
.B1(n_290),
.B2(n_293),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_386),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_311),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_388),
.B(n_395),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_353),
.A2(n_320),
.B1(n_310),
.B2(n_325),
.Y(n_389)
);

AO22x1_ASAP7_75t_L g391 ( 
.A1(n_340),
.A2(n_311),
.B1(n_310),
.B2(n_315),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_356),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_392),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_348),
.B(n_288),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_340),
.A2(n_286),
.B(n_322),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_308),
.C(n_315),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_402),
.C(n_333),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_363),
.B(n_359),
.C(n_368),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_346),
.A2(n_327),
.B1(n_325),
.B2(n_322),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_354),
.A2(n_327),
.B1(n_319),
.B2(n_302),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_324),
.B1(n_302),
.B2(n_319),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_407),
.A2(n_366),
.B1(n_367),
.B2(n_371),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_381),
.A2(n_343),
.B1(n_369),
.B2(n_357),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_409),
.A2(n_417),
.B1(n_424),
.B2(n_431),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_410),
.A2(n_415),
.B1(n_421),
.B2(n_435),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_412),
.A2(n_434),
.B(n_429),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_388),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_416),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_393),
.B(n_385),
.Y(n_414)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_414),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_381),
.A2(n_336),
.B1(n_337),
.B2(n_352),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_347),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_406),
.A2(n_369),
.B1(n_351),
.B2(n_362),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_375),
.Y(n_418)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_418),
.Y(n_445)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_377),
.Y(n_419)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_419),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_372),
.Y(n_420)
);

OAI21xp33_ASAP7_75t_L g443 ( 
.A1(n_420),
.A2(n_422),
.B(n_385),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_407),
.A2(n_358),
.B1(n_333),
.B2(n_342),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_393),
.B(n_344),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_402),
.C(n_390),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_389),
.A2(n_369),
.B1(n_364),
.B2(n_339),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_425),
.Y(n_444)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_378),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_427),
.Y(n_450)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_399),
.Y(n_428)
);

NAND4xp25_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_432),
.C(n_405),
.D(n_284),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_382),
.A2(n_345),
.B1(n_361),
.B2(n_373),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_399),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_403),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_433),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_384),
.A2(n_391),
.B1(n_376),
.B2(n_387),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_386),
.A2(n_365),
.B1(n_355),
.B2(n_341),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_384),
.A2(n_360),
.B1(n_319),
.B2(n_321),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_436),
.A2(n_387),
.B1(n_380),
.B2(n_397),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_390),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_440),
.B(n_457),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_464),
.C(n_430),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_451),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_415),
.A2(n_384),
.B1(n_401),
.B2(n_391),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_446),
.A2(n_448),
.B1(n_454),
.B2(n_456),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_447),
.A2(n_449),
.B1(n_424),
.B2(n_431),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_433),
.A2(n_396),
.B1(n_404),
.B2(n_392),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_409),
.A2(n_404),
.B1(n_396),
.B2(n_394),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_429),
.A2(n_380),
.B(n_374),
.Y(n_451)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_421),
.A2(n_435),
.B1(n_408),
.B2(n_411),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_455),
.B(n_410),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_408),
.A2(n_394),
.B1(n_398),
.B2(n_383),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_395),
.Y(n_457)
);

MAJx2_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_405),
.C(n_288),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_SL g473 ( 
.A(n_459),
.B(n_412),
.C(n_413),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_420),
.B(n_288),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_462),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_430),
.B(n_332),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_411),
.A2(n_383),
.B1(n_321),
.B2(n_324),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_463),
.A2(n_417),
.B1(n_436),
.B2(n_434),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_332),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_467),
.C(n_468),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_422),
.C(n_414),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_457),
.C(n_464),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_450),
.Y(n_469)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_459),
.C(n_456),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_470),
.B(n_487),
.C(n_444),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_481),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_477),
.Y(n_497)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_460),
.Y(n_474)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_448),
.B(n_434),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_479),
.A2(n_486),
.B1(n_439),
.B2(n_447),
.Y(n_493)
);

BUFx12f_ASAP7_75t_L g480 ( 
.A(n_451),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_480),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_444),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_461),
.B(n_416),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_299),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_445),
.B(n_418),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_484),
.Y(n_496)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_460),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_485),
.A2(n_438),
.B(n_463),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_439),
.A2(n_432),
.B1(n_428),
.B2(n_427),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_441),
.B(n_419),
.C(n_425),
.Y(n_487)
);

OAI322xp33_ASAP7_75t_L g491 ( 
.A1(n_478),
.A2(n_458),
.A3(n_452),
.B1(n_455),
.B2(n_449),
.C1(n_446),
.C2(n_438),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_491),
.B(n_494),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_454),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_470),
.C(n_465),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_493),
.A2(n_498),
.B1(n_316),
.B2(n_284),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_500),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_475),
.A2(n_458),
.B1(n_426),
.B2(n_286),
.Y(n_498)
);

NOR2xp67_ASAP7_75t_R g499 ( 
.A(n_480),
.B(n_314),
.Y(n_499)
);

O2A1O1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_499),
.A2(n_480),
.B(n_466),
.C(n_471),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_476),
.B(n_482),
.Y(n_500)
);

AOI221xp5_ASAP7_75t_L g502 ( 
.A1(n_487),
.A2(n_296),
.B1(n_299),
.B2(n_314),
.C(n_355),
.Y(n_502)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_502),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_504),
.B(n_505),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_467),
.B(n_316),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_506),
.B(n_497),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_496),
.Y(n_507)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_507),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_486),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_508),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_517),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_477),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_513),
.B(n_514),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_503),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_468),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_516),
.C(n_500),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_489),
.B(n_472),
.C(n_473),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_501),
.B(n_472),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_518),
.A2(n_498),
.B1(n_493),
.B2(n_504),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_488),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_521),
.B(n_524),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_506),
.B(n_489),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_510),
.A2(n_499),
.B1(n_497),
.B2(n_495),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_526),
.B(n_529),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_527),
.B(n_528),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_505),
.C(n_492),
.Y(n_528)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_530),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_519),
.B(n_275),
.C(n_316),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_531),
.B(n_518),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_509),
.B(n_514),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_532),
.A2(n_520),
.B1(n_226),
.B2(n_276),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_517),
.C(n_508),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_533),
.B(n_535),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_523),
.A2(n_522),
.B(n_528),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_523),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_536),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_525),
.A2(n_511),
.B(n_512),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_538),
.A2(n_536),
.B(n_537),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_540),
.B(n_525),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_539),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_543),
.A2(n_544),
.B1(n_546),
.B2(n_226),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_534),
.Y(n_544)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_545),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_547),
.B(n_215),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_541),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_549),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_548),
.B(n_538),
.C(n_228),
.Y(n_550)
);

AOI21x1_ASAP7_75t_L g555 ( 
.A1(n_550),
.A2(n_553),
.B(n_548),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_551),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_555),
.A2(n_234),
.B1(n_242),
.B2(n_239),
.Y(n_558)
);

MAJx2_ASAP7_75t_L g557 ( 
.A(n_554),
.B(n_552),
.C(n_550),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_557),
.A2(n_558),
.B(n_556),
.Y(n_559)
);

AOI221xp5_ASAP7_75t_L g560 ( 
.A1(n_559),
.A2(n_247),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_560),
.A2(n_15),
.B(n_18),
.Y(n_561)
);


endmodule