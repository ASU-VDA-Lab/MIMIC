module fake_jpeg_7743_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_0),
.B(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_2),
.C(n_3),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_2),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_32),
.B1(n_18),
.B2(n_31),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_58),
.B(n_68),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_33),
.B1(n_31),
.B2(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_57),
.B1(n_62),
.B2(n_21),
.Y(n_72)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_44),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_33),
.B1(n_30),
.B2(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_32),
.B1(n_18),
.B2(n_24),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_29),
.B1(n_22),
.B2(n_24),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_44),
.B1(n_4),
.B2(n_38),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_22),
.B1(n_27),
.B2(n_23),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_36),
.B(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_26),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_21),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_16),
.B1(n_25),
.B2(n_6),
.Y(n_68)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_81),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_85),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_43),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_47),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_40),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_79),
.B(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_3),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_3),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_43),
.B(n_25),
.C(n_38),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_53),
.B(n_61),
.C(n_55),
.Y(n_104)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_4),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_46),
.Y(n_95)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_101),
.B(n_104),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_4),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_65),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_97),
.C(n_112),
.Y(n_123)
);

BUFx24_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_55),
.B(n_46),
.C(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_83),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_55),
.B1(n_8),
.B2(n_9),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_113),
.A2(n_117),
.B1(n_89),
.B2(n_87),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_7),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_13),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_126),
.B1(n_71),
.B2(n_81),
.Y(n_154)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_76),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_124),
.C(n_117),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_75),
.C(n_94),
.Y(n_124)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_75),
.C(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_129),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_78),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_74),
.Y(n_128)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_84),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_107),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_133),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_70),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_137),
.C(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_101),
.B(n_104),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_127),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_146),
.C(n_149),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_101),
.C(n_114),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_108),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_126),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_130),
.B(n_133),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_83),
.B1(n_99),
.B2(n_90),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_105),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_105),
.B(n_98),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_129),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_162),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_131),
.C(n_136),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_159),
.C(n_161),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_119),
.C(n_118),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_150),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_167),
.Y(n_170)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_155),
.C(n_159),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_154),
.B1(n_140),
.B2(n_145),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_174),
.A2(n_177),
.B1(n_142),
.B2(n_158),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_150),
.B1(n_152),
.B2(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_184),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_180),
.C(n_169),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_155),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_161),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_183),
.B(n_168),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_148),
.B(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_170),
.B(n_137),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_185),
.A2(n_178),
.B(n_177),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_171),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.C(n_180),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_176),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_189),
.A2(n_183),
.B(n_173),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_191),
.B(n_193),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_SL g193 ( 
.A1(n_186),
.A2(n_175),
.B(n_181),
.C(n_146),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_130),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_189),
.B(n_134),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_198),
.B(n_195),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_91),
.C(n_90),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_14),
.Y(n_200)
);


endmodule