module fake_jpeg_3469_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_43;
wire n_37;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_6),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_21),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_8),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_20),
.B1(n_23),
.B2(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_16),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_11),
.A2(n_0),
.B1(n_3),
.B2(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_9),
.A2(n_12),
.B1(n_16),
.B2(n_10),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_20),
.B1(n_12),
.B2(n_14),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_16),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_18),
.B(n_19),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_39),
.C(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_22),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_44),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

FAx1_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_38),
.CI(n_37),
.CON(n_44),
.SN(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_49),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_39),
.B1(n_40),
.B2(n_29),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_42),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_53),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_44),
.B1(n_45),
.B2(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

AOI322xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_52),
.A3(n_53),
.B1(n_14),
.B2(n_50),
.C1(n_15),
.C2(n_29),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_50),
.C(n_55),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_55),
.C(n_15),
.Y(n_59)
);


endmodule