module fake_jpeg_28575_n_387 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_387);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_387;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_41),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_42),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_20),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_56),
.Y(n_85)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_51),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_58),
.Y(n_87)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_57),
.Y(n_95)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

NOR2xp67_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_37),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_34),
.CON(n_94),
.SN(n_94)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_60),
.Y(n_66)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_63),
.B(n_30),
.Y(n_72)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_27),
.B(n_0),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_65),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_21),
.B1(n_25),
.B2(n_36),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_67),
.A2(n_70),
.B1(n_78),
.B2(n_44),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_27),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_76),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_21),
.B1(n_25),
.B2(n_36),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_72),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_27),
.B1(n_37),
.B2(n_26),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_35),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_17),
.B(n_22),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_89),
.C(n_85),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_19),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_34),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_77),
.B(n_32),
.Y(n_107)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_36),
.B1(n_21),
.B2(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_38),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_39),
.B(n_0),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_43),
.A2(n_29),
.B1(n_36),
.B2(n_25),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_91),
.B1(n_39),
.B2(n_30),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_29),
.B1(n_30),
.B2(n_17),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_38),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_46),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_15),
.Y(n_116)
);

CKINVDCx6p67_ASAP7_75t_R g102 ( 
.A(n_100),
.Y(n_102)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_49),
.B(n_40),
.C(n_51),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_105),
.B(n_111),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_41),
.A3(n_42),
.B1(n_17),
.B2(n_32),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_109),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_107),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_65),
.A3(n_42),
.B1(n_22),
.B2(n_60),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_35),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_116),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_115),
.B(n_125),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_33),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_121),
.Y(n_163)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_75),
.B(n_15),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_123),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_33),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_126),
.B1(n_70),
.B2(n_89),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_67),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_46),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_130),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_62),
.B1(n_47),
.B2(n_53),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_46),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_77),
.B(n_14),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_132),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_98),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_134),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_114),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_66),
.B(n_33),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_100),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_165),
.B1(n_168),
.B2(n_95),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_85),
.B(n_95),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_143),
.A2(n_88),
.B(n_82),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_144),
.B(n_131),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_145),
.B(n_156),
.C(n_159),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_112),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_103),
.Y(n_180)
);

OR2x4_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_113),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g204 ( 
.A1(n_154),
.A2(n_98),
.B(n_30),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_89),
.C(n_85),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_95),
.C(n_66),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_102),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_78),
.B1(n_96),
.B2(n_62),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_115),
.A2(n_78),
.B1(n_74),
.B2(n_69),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_185),
.B1(n_191),
.B2(n_192),
.Y(n_222)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_103),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_176),
.Y(n_225)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_179),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_195),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_190),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_121),
.B1(n_117),
.B2(n_106),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_182),
.A2(n_183),
.B1(n_188),
.B2(n_196),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_105),
.B1(n_135),
.B2(n_129),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_127),
.B1(n_125),
.B2(n_138),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_130),
.B1(n_74),
.B2(n_69),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_163),
.B(n_111),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_140),
.A2(n_57),
.B1(n_50),
.B2(n_44),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_50),
.B1(n_57),
.B2(n_136),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_143),
.A2(n_102),
.B(n_133),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_206),
.B(n_207),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_134),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_161),
.B1(n_173),
.B2(n_168),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_158),
.A2(n_161),
.B1(n_149),
.B2(n_172),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_197),
.A2(n_148),
.B1(n_53),
.B2(n_47),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_149),
.A2(n_52),
.B1(n_55),
.B2(n_82),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_202),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_203),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_145),
.B(n_102),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_204),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_201),
.A2(n_132),
.B(n_146),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_142),
.B(n_101),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_146),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_132),
.B(n_1),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_159),
.A2(n_155),
.B(n_142),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_189),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_190),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_209),
.B(n_215),
.Y(n_271)
);

AOI22x1_ASAP7_75t_SL g212 ( 
.A1(n_199),
.A2(n_147),
.B1(n_154),
.B2(n_155),
.Y(n_212)
);

AO21x1_ASAP7_75t_L g270 ( 
.A1(n_212),
.A2(n_230),
.B(n_179),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_189),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_153),
.B(n_160),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_217),
.A2(n_220),
.B(n_229),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_156),
.C(n_153),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_218),
.B(n_178),
.C(n_194),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_206),
.B(n_197),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_151),
.B1(n_147),
.B2(n_141),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_221),
.A2(n_238),
.B1(n_215),
.B2(n_217),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_151),
.B1(n_160),
.B2(n_141),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_232),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_162),
.Y(n_232)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_195),
.B(n_98),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_234),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_186),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_237),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_132),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_175),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_187),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_0),
.B(n_2),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_198),
.Y(n_253)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_242),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_243),
.Y(n_281)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_223),
.B(n_176),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_245),
.B(n_247),
.Y(n_287)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_252),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_222),
.A2(n_174),
.B1(n_188),
.B2(n_191),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_216),
.B1(n_221),
.B2(n_210),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_254),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_200),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_255),
.A2(n_267),
.B1(n_268),
.B2(n_234),
.Y(n_279)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_257),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_211),
.B(n_205),
.Y(n_257)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_260),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_224),
.B(n_177),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_270),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_223),
.B(n_177),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_218),
.C(n_224),
.Y(n_273)
);

XOR2x1_ASAP7_75t_SL g263 ( 
.A(n_220),
.B(n_184),
.Y(n_263)
);

AOI21xp33_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_264),
.B(n_226),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_225),
.B(n_232),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_278),
.C(n_291),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_275),
.A2(n_276),
.B1(n_280),
.B2(n_285),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_250),
.A2(n_216),
.B1(n_210),
.B2(n_234),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_234),
.C(n_222),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_269),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_238),
.B1(n_230),
.B2(n_240),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_255),
.A2(n_229),
.B1(n_219),
.B2(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_258),
.A2(n_237),
.B1(n_219),
.B2(n_228),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_249),
.A2(n_233),
.B1(n_213),
.B2(n_239),
.Y(n_289)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_249),
.A2(n_271),
.B1(n_260),
.B2(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_148),
.C(n_236),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_269),
.A2(n_236),
.B1(n_101),
.B2(n_96),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_244),
.B1(n_265),
.B2(n_256),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_261),
.A2(n_101),
.B1(n_55),
.B2(n_52),
.Y(n_294)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_261),
.B(n_270),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_299),
.A2(n_308),
.B(n_0),
.Y(n_335)
);

BUFx12_ASAP7_75t_L g300 ( 
.A(n_291),
.Y(n_300)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_271),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_301),
.Y(n_321)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_303),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_273),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_314),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_306),
.B(n_309),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_276),
.A2(n_253),
.B(n_251),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_254),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_259),
.C(n_251),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_293),
.C(n_294),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_286),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_312),
.A2(n_318),
.B1(n_296),
.B2(n_277),
.Y(n_326)
);

A2O1A1O1Ixp25_ASAP7_75t_L g314 ( 
.A1(n_295),
.A2(n_287),
.B(n_284),
.C(n_286),
.D(n_293),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_295),
.A2(n_268),
.B(n_267),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_285),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_275),
.B(n_246),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_30),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_329),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_323),
.B(n_327),
.Y(n_344)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_326),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_317),
.A2(n_296),
.B1(n_266),
.B2(n_281),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_292),
.C(n_242),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_298),
.A2(n_243),
.B1(n_96),
.B2(n_60),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_330),
.B(n_333),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_332),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_304),
.B(n_7),
.Y(n_332)
);

XNOR2x1_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_7),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_298),
.A2(n_7),
.B1(n_16),
.B2(n_13),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_321),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_335),
.A2(n_315),
.B(n_303),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_322),
.A2(n_299),
.B(n_310),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_9),
.Y(n_361)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_339),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_320),
.A2(n_297),
.B1(n_308),
.B2(n_313),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_342),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_341),
.A2(n_334),
.B1(n_331),
.B2(n_324),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_300),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_306),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_348),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_323),
.A2(n_305),
.B(n_302),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_300),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_319),
.A2(n_307),
.B1(n_316),
.B2(n_314),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_347),
.A2(n_8),
.B1(n_13),
.B2(n_10),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_307),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_330),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_6),
.Y(n_360)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_352),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_337),
.A2(n_324),
.B1(n_333),
.B2(n_332),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_355),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_8),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_349),
.C(n_346),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_357),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_SL g359 ( 
.A(n_338),
.B(n_6),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_359),
.A2(n_349),
.B(n_9),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_360),
.B(n_361),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_344),
.B(n_9),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_362),
.B(n_10),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_340),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_367),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_351),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_368),
.B(n_371),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_358),
.A2(n_347),
.B(n_341),
.Y(n_369)
);

AO21x1_ASAP7_75t_L g377 ( 
.A1(n_369),
.A2(n_3),
.B(n_4),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_372),
.B(n_33),
.C(n_4),
.Y(n_379)
);

AOI322xp5_ASAP7_75t_L g374 ( 
.A1(n_368),
.A2(n_357),
.A3(n_361),
.B1(n_356),
.B2(n_346),
.C1(n_2),
.C2(n_5),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_374),
.A2(n_376),
.B1(n_365),
.B2(n_370),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_365),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_376)
);

AOI21x1_ASAP7_75t_L g381 ( 
.A1(n_377),
.A2(n_378),
.B(n_366),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_SL g378 ( 
.A(n_364),
.B(n_33),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_379),
.A2(n_4),
.B(n_5),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_381),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_375),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_382),
.A2(n_383),
.B(n_373),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_384),
.A2(n_374),
.B(n_5),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_385),
.Y(n_387)
);


endmodule