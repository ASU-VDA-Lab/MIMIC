module fake_jpeg_1413_n_52 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_31;
wire n_17;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_7),
.B(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_20),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_19),
.A2(n_30),
.B1(n_31),
.B2(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_23),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_6),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B(n_29),
.Y(n_32)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

AOI21xp33_ASAP7_75t_SL g29 ( 
.A1(n_10),
.A2(n_16),
.B(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_17),
.A2(n_15),
.B1(n_10),
.B2(n_9),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_21),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_30),
.B1(n_28),
.B2(n_23),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_43),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_37),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_43),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_39),
.B1(n_35),
.B2(n_41),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_44),
.B(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_50),
.A2(n_47),
.B(n_45),
.Y(n_51)
);

OAI21x1_ASAP7_75t_SL g52 ( 
.A1(n_51),
.A2(n_36),
.B(n_42),
.Y(n_52)
);


endmodule