module fake_jpeg_23182_n_138 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx10_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_30),
.B(n_32),
.Y(n_55)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_33),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_25),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_15),
.B1(n_29),
.B2(n_26),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_49),
.B1(n_51),
.B2(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_26),
.B1(n_17),
.B2(n_25),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_22),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_37),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_30),
.B1(n_36),
.B2(n_35),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_48),
.B1(n_32),
.B2(n_27),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_28),
.B1(n_19),
.B2(n_23),
.Y(n_49)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_20),
.B1(n_24),
.B2(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_45),
.Y(n_65)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_3),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_45),
.B(n_50),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_30),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_62),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_24),
.B1(n_21),
.B2(n_14),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_61),
.B1(n_68),
.B2(n_69),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_32),
.B1(n_38),
.B2(n_14),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_65),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_70),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_38),
.B1(n_5),
.B2(n_4),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_8),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_70),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_43),
.B(n_53),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_57),
.C(n_64),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_56),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_81),
.C(n_79),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_93),
.Y(n_108)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_43),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_80),
.B1(n_68),
.B2(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_99),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_65),
.C(n_74),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_91),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_77),
.B(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_77),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_102),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_78),
.B1(n_88),
.B2(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

OAI322xp33_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_112),
.A3(n_106),
.B1(n_107),
.B2(n_110),
.C1(n_109),
.C2(n_103),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_63),
.B(n_44),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_82),
.C(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_112),
.B(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_119),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_85),
.B(n_96),
.C(n_99),
.D(n_101),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_116),
.C(n_118),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_106),
.Y(n_121)
);

XOR2x2_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_53),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_111),
.B(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_120),
.A2(n_111),
.B1(n_104),
.B2(n_54),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_124),
.B1(n_116),
.B2(n_44),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_54),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_126),
.B(n_54),
.Y(n_129)
);

OAI21x1_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_117),
.B(n_115),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_130),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_125),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_131),
.B(n_133),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_121),
.Y(n_134)
);

OAI321xp33_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_44),
.A3(n_72),
.B1(n_73),
.B2(n_132),
.C(n_133),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_136),
.Y(n_138)
);


endmodule