module fake_ibex_470_n_665 (n_64, n_3, n_73, n_65, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_70, n_7, n_20, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_13, n_61, n_14, n_0, n_12, n_42, n_77, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_83, n_32, n_53, n_50, n_11, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_54, n_19, n_665);

input n_64;
input n_3;
input n_73;
input n_65;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_70;
input n_7;
input n_20;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_13;
input n_61;
input n_14;
input n_0;
input n_12;
input n_42;
input n_77;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_54;
input n_19;

output n_665;

wire n_151;
wire n_85;
wire n_599;
wire n_507;
wire n_540;
wire n_395;
wire n_84;
wire n_171;
wire n_103;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_108;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_452;
wire n_86;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_638;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_94;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_457;
wire n_88;
wire n_357;
wire n_412;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_90;
wire n_449;
wire n_547;
wire n_176;
wire n_216;
wire n_652;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_645;
wire n_500;
wire n_542;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_556;
wire n_189;
wire n_498;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_89;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_561;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_91;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_228;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_106;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_550;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_109;
wire n_127;
wire n_121;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_122;
wire n_523;
wire n_116;
wire n_614;
wire n_370;
wire n_431;
wire n_574;
wire n_289;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_136;
wire n_261;
wire n_521;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_654;
wire n_656;
wire n_437;
wire n_602;
wire n_355;
wire n_474;
wire n_594;
wire n_636;
wire n_407;
wire n_102;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_99;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_623;
wire n_585;
wire n_530;
wire n_356;
wire n_104;
wire n_420;
wire n_543;
wire n_483;
wire n_580;
wire n_141;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_576;
wire n_230;
wire n_96;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_618;
wire n_488;
wire n_139;
wire n_514;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_98;
wire n_129;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_87;
wire n_262;
wire n_439;
wire n_433;
wire n_643;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_554;
wire n_553;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_605;
wire n_539;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_624;
wire n_411;
wire n_135;
wire n_520;
wire n_658;
wire n_512;
wire n_615;
wire n_283;
wire n_366;
wire n_397;
wire n_111;
wire n_627;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_92;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_650;
wire n_409;
wire n_582;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_633;
wire n_532;
wire n_95;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_118;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_639;
wire n_303;
wire n_362;
wire n_93;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_97;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_631;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_160;
wire n_657;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVxp33_ASAP7_75t_SL g85 ( 
.A(n_1),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_15),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_43),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_5),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_5),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_24),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_0),
.Y(n_105)
);

INVxp67_ASAP7_75t_SL g106 ( 
.A(n_70),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_59),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_16),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_14),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_15),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_21),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_7),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_48),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_11),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_37),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_35),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_42),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_27),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_3),
.Y(n_132)
);

INVxp33_ASAP7_75t_SL g133 ( 
.A(n_50),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_7),
.Y(n_134)
);

NOR2xp67_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_61),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_0),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_38),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVxp33_ASAP7_75t_SL g139 ( 
.A(n_77),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_22),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_14),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_26),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_52),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_8),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_3),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_4),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g149 ( 
.A(n_8),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_80),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_6),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_51),
.Y(n_152)
);

INVx4_ASAP7_75t_R g153 ( 
.A(n_30),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_34),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_17),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_92),
.Y(n_157)
);

OAI21x1_ASAP7_75t_L g158 ( 
.A1(n_84),
.A2(n_31),
.B(n_71),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_2),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_94),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_9),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_104),
.B(n_9),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_98),
.B(n_10),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_118),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_118),
.B(n_10),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_112),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_136),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_86),
.B(n_11),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_91),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_85),
.B(n_12),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_98),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_127),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_R g196 ( 
.A(n_87),
.B(n_40),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_110),
.B(n_12),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_127),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_110),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_151),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_93),
.B(n_13),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_141),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_95),
.A2(n_44),
.B(n_64),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_151),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_87),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_90),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_90),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_117),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_147),
.B(n_13),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_107),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_128),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_128),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_133),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_96),
.A2(n_36),
.B(n_63),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_131),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_99),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_102),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_133),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_103),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_108),
.B(n_16),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_113),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_114),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_115),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_139),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_111),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_165),
.B(n_154),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_139),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_119),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_169),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_111),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_159),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_116),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_111),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_159),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_169),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_159),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_169),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_145),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_169),
.Y(n_253)
);

AO22x2_ASAP7_75t_L g254 ( 
.A1(n_161),
.A2(n_129),
.B1(n_152),
.B2(n_144),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_168),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_169),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_179),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_199),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_210),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_171),
.Y(n_260)
);

AND2x4_ASAP7_75t_L g261 ( 
.A(n_161),
.B(n_163),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_214),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_140),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_212),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_189),
.B(n_126),
.C(n_143),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_192),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_212),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_186),
.Y(n_269)
);

AO22x2_ASAP7_75t_L g270 ( 
.A1(n_163),
.A2(n_124),
.B1(n_138),
.B2(n_137),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_187),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_192),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_192),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_199),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_221),
.B(n_226),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_130),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_193),
.A2(n_85),
.B1(n_111),
.B2(n_97),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_208),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_164),
.B(n_111),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_229),
.B(n_225),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_164),
.B(n_125),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g283 ( 
.A(n_182),
.B(n_122),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_192),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_211),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_200),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_205),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_205),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_225),
.B(n_106),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_205),
.Y(n_290)
);

NAND2x1p5_ASAP7_75t_L g291 ( 
.A(n_197),
.B(n_121),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_205),
.Y(n_292)
);

AO22x2_ASAP7_75t_L g293 ( 
.A1(n_197),
.A2(n_101),
.B1(n_17),
.B2(n_153),
.Y(n_293)
);

AND2x6_ASAP7_75t_L g294 ( 
.A(n_231),
.B(n_135),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_226),
.B(n_18),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_231),
.B(n_20),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_188),
.B(n_23),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_205),
.Y(n_298)
);

AO22x2_ASAP7_75t_L g299 ( 
.A1(n_193),
.A2(n_25),
.B1(n_45),
.B2(n_55),
.Y(n_299)
);

OR2x2_ASAP7_75t_SL g300 ( 
.A(n_170),
.B(n_56),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_158),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_191),
.B(n_57),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_160),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_160),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_202),
.Y(n_305)
);

AO22x2_ASAP7_75t_L g306 ( 
.A1(n_177),
.A2(n_72),
.B1(n_203),
.B2(n_213),
.Y(n_306)
);

AND2x4_ASAP7_75t_L g307 ( 
.A(n_204),
.B(n_185),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_172),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_174),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_158),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_176),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_166),
.B(n_190),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_228),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_166),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_206),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_173),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_211),
.B(n_215),
.Y(n_317)
);

OAI221xp5_ASAP7_75t_L g318 ( 
.A1(n_201),
.A2(n_207),
.B1(n_223),
.B2(n_173),
.C(n_175),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_175),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_190),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_209),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_180),
.A2(n_181),
.B1(n_198),
.B2(n_195),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_209),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_223),
.B(n_220),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_178),
.B(n_183),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_215),
.B(n_220),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_303),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_280),
.Y(n_328)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_280),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_247),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_257),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_322),
.Y(n_332)
);

AND2x2_ASAP7_75t_SL g333 ( 
.A(n_261),
.B(n_206),
.Y(n_333)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_316),
.Y(n_334)
);

OR2x6_ASAP7_75t_SL g335 ( 
.A(n_286),
.B(n_198),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_240),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_269),
.B(n_219),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_257),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_306),
.A2(n_293),
.B1(n_299),
.B2(n_313),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_247),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_258),
.Y(n_341)
);

NAND2xp33_ASAP7_75t_SL g342 ( 
.A(n_324),
.B(n_326),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_269),
.B(n_219),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_289),
.B(n_178),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_274),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_289),
.B(n_183),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_235),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_261),
.B(n_207),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_243),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_250),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_262),
.B(n_232),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_279),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_241),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_240),
.Y(n_354)
);

AO22x1_ASAP7_75t_L g355 ( 
.A1(n_317),
.A2(n_195),
.B1(n_157),
.B2(n_162),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_239),
.B(n_184),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_241),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_281),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_239),
.B(n_157),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_291),
.B(n_162),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_276),
.B(n_232),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_285),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_291),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_263),
.B(n_184),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_244),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_237),
.B(n_282),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_244),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_282),
.B(n_196),
.Y(n_369)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_303),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_236),
.B(n_206),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_271),
.B(n_222),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_281),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_R g375 ( 
.A(n_259),
.B(n_222),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_314),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_314),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_222),
.Y(n_378)
);

OR2x6_ASAP7_75t_L g379 ( 
.A(n_299),
.B(n_293),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_248),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_301),
.Y(n_381)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_238),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_305),
.B(n_307),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_245),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_234),
.B(n_242),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_254),
.A2(n_270),
.B1(n_326),
.B2(n_318),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_266),
.B(n_234),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_322),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_275),
.A2(n_270),
.B1(n_254),
.B2(n_277),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_265),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_268),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_242),
.B(n_264),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_308),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_309),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_306),
.Y(n_396)
);

NOR3xp33_ASAP7_75t_SL g397 ( 
.A(n_277),
.B(n_266),
.C(n_325),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_320),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_251),
.Y(n_399)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_301),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_253),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_301),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_283),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_300),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_311),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_R g406 ( 
.A(n_295),
.B(n_310),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_272),
.Y(n_407)
);

CKINVDCx11_ASAP7_75t_R g408 ( 
.A(n_335),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_358),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_260),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_340),
.Y(n_414)
);

OAI21x1_ASAP7_75t_SL g415 ( 
.A1(n_339),
.A2(n_297),
.B(n_302),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_362),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_R g418 ( 
.A(n_332),
.B(n_249),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_379),
.A2(n_318),
.B1(n_255),
.B2(n_252),
.Y(n_419)
);

CKINVDCx8_ASAP7_75t_R g420 ( 
.A(n_379),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_264),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_405),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_252),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_341),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_378),
.A2(n_312),
.B(n_315),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_331),
.B(n_310),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_352),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_338),
.B(n_310),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_312),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_345),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_363),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_405),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_386),
.B(n_321),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_348),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_348),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_336),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_348),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_339),
.A2(n_302),
.B1(n_297),
.B2(n_296),
.Y(n_438)
);

BUFx4f_ASAP7_75t_L g439 ( 
.A(n_379),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_334),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_378),
.A2(n_342),
.B(n_373),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_396),
.A2(n_294),
.B1(n_319),
.B2(n_304),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_336),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_367),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_354),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_354),
.Y(n_446)
);

AOI21xp33_ASAP7_75t_L g447 ( 
.A1(n_371),
.A2(n_296),
.B(n_323),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_333),
.A2(n_315),
.B(n_287),
.Y(n_448)
);

OAI22xp33_ASAP7_75t_L g449 ( 
.A1(n_390),
.A2(n_315),
.B1(n_246),
.B2(n_256),
.Y(n_449)
);

BUFx12f_ASAP7_75t_L g450 ( 
.A(n_403),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_351),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_387),
.A2(n_298),
.B1(n_292),
.B2(n_290),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_372),
.B(n_294),
.Y(n_453)
);

OR2x6_ASAP7_75t_L g454 ( 
.A(n_355),
.B(n_238),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_365),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_351),
.A2(n_294),
.B1(n_273),
.B2(n_288),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_370),
.Y(n_457)
);

BUFx10_ASAP7_75t_L g458 ( 
.A(n_351),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_334),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_334),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_359),
.B(n_294),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_334),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_394),
.A2(n_238),
.B1(n_246),
.B2(n_256),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_370),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_360),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_372),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_334),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_365),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_333),
.A2(n_246),
.B(n_256),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_356),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_342),
.A2(n_267),
.B(n_278),
.C(n_284),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g472 ( 
.A(n_361),
.B(n_267),
.C(n_278),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_366),
.B(n_267),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_368),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_327),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_364),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_381),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_395),
.B(n_278),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_332),
.Y(n_479)
);

OAI21xp33_ASAP7_75t_SL g480 ( 
.A1(n_392),
.A2(n_284),
.B(n_380),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_347),
.B(n_284),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_361),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_426),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_419),
.A2(n_384),
.B1(n_397),
.B2(n_349),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_409),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_411),
.B(n_404),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_411),
.B(n_343),
.Y(n_488)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_457),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_L g490 ( 
.A1(n_439),
.A2(n_389),
.B1(n_403),
.B2(n_369),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_433),
.B(n_337),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_424),
.B(n_344),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_426),
.Y(n_493)
);

OAI22xp33_ASAP7_75t_L g494 ( 
.A1(n_439),
.A2(n_389),
.B1(n_368),
.B2(n_329),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_459),
.B(n_375),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_417),
.B(n_346),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_416),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_417),
.B(n_364),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_428),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_433),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_473),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_438),
.A2(n_423),
.B1(n_421),
.B2(n_429),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_438),
.A2(n_328),
.B1(n_329),
.B2(n_391),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_420),
.A2(n_328),
.B1(n_329),
.B2(n_391),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_428),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_421),
.A2(n_328),
.B1(n_364),
.B2(n_370),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_423),
.A2(n_353),
.B1(n_357),
.B2(n_385),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_476),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_475),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_451),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_481),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_412),
.B(n_353),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_408),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_429),
.A2(n_353),
.B1(n_385),
.B2(n_327),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_430),
.B(n_431),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_441),
.A2(n_425),
.B(n_448),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_436),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_415),
.A2(n_385),
.B1(n_376),
.B2(n_377),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_461),
.A2(n_398),
.B1(n_376),
.B2(n_377),
.Y(n_519)
);

INVx6_ASAP7_75t_L g520 ( 
.A(n_458),
.Y(n_520)
);

OAI22xp33_ASAP7_75t_L g521 ( 
.A1(n_459),
.A2(n_402),
.B1(n_400),
.B2(n_381),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_435),
.B(n_398),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_481),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_478),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_L g525 ( 
.A1(n_454),
.A2(n_400),
.B1(n_402),
.B2(n_381),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_479),
.A2(n_400),
.B1(n_402),
.B2(n_383),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_427),
.B(n_383),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_437),
.B(n_375),
.Y(n_528)
);

A2O1A1Ixp33_ASAP7_75t_L g529 ( 
.A1(n_447),
.A2(n_399),
.B(n_401),
.C(n_407),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_477),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_L g531 ( 
.A(n_477),
.B(n_406),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_448),
.A2(n_381),
.B(n_399),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_442),
.A2(n_406),
.B1(n_382),
.B2(n_401),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_449),
.A2(n_382),
.B1(n_407),
.B2(n_452),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_427),
.B(n_382),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_414),
.Y(n_536)
);

OAI22xp33_ASAP7_75t_L g537 ( 
.A1(n_454),
.A2(n_434),
.B1(n_456),
.B2(n_452),
.Y(n_537)
);

OA21x2_ASAP7_75t_L g538 ( 
.A1(n_469),
.A2(n_382),
.B(n_447),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_457),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_418),
.Y(n_540)
);

O2A1O1Ixp33_ASAP7_75t_L g541 ( 
.A1(n_465),
.A2(n_480),
.B(n_445),
.C(n_446),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_SL g542 ( 
.A(n_477),
.B(n_432),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_422),
.A2(n_454),
.B1(n_440),
.B2(n_467),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_458),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_450),
.Y(n_545)
);

AOI21x1_ASAP7_75t_L g546 ( 
.A1(n_469),
.A2(n_463),
.B(n_472),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_R g547 ( 
.A(n_444),
.B(n_464),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_466),
.B(n_453),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_482),
.A2(n_453),
.B1(n_443),
.B2(n_455),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g550 ( 
.A1(n_516),
.A2(n_471),
.B(n_478),
.Y(n_550)
);

CKINVDCx14_ASAP7_75t_R g551 ( 
.A(n_513),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_500),
.A2(n_468),
.B1(n_474),
.B2(n_464),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_488),
.B(n_413),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_532),
.A2(n_463),
.B(n_460),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_489),
.B(n_462),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_546),
.A2(n_538),
.B(n_518),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_502),
.A2(n_484),
.B1(n_491),
.B2(n_494),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_502),
.B(n_487),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_540),
.A2(n_494),
.B1(n_486),
.B2(n_498),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_503),
.A2(n_528),
.B1(n_490),
.B2(n_506),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_SL g561 ( 
.A(n_547),
.B(n_495),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_485),
.B(n_523),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_503),
.A2(n_490),
.B1(n_506),
.B2(n_527),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_530),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_547),
.A2(n_536),
.B1(n_513),
.B2(n_497),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_509),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_530),
.Y(n_567)
);

A2O1A1Ixp33_ASAP7_75t_L g568 ( 
.A1(n_541),
.A2(n_518),
.B(n_507),
.C(n_514),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_515),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_530),
.Y(n_570)
);

AOI21x1_ASAP7_75t_L g571 ( 
.A1(n_538),
.A2(n_495),
.B(n_534),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_527),
.A2(n_501),
.B1(n_510),
.B2(n_537),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_537),
.A2(n_492),
.B1(n_496),
.B2(n_515),
.Y(n_573)
);

OAI221xp5_ASAP7_75t_L g574 ( 
.A1(n_515),
.A2(n_507),
.B1(n_519),
.B2(n_514),
.C(n_517),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_512),
.A2(n_497),
.B1(n_504),
.B2(n_508),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_511),
.A2(n_524),
.B1(n_525),
.B2(n_543),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_529),
.A2(n_521),
.B(n_519),
.Y(n_577)
);

OAI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_520),
.A2(n_489),
.B1(n_535),
.B2(n_544),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_526),
.A2(n_548),
.B1(n_522),
.B2(n_493),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_483),
.Y(n_580)
);

OA21x2_ASAP7_75t_L g581 ( 
.A1(n_529),
.A2(n_499),
.B(n_505),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_539),
.B(n_489),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_545),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_520),
.A2(n_535),
.B1(n_489),
.B2(n_539),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_520),
.B(n_530),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_542),
.A2(n_538),
.B1(n_525),
.B2(n_533),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_542),
.A2(n_379),
.B1(n_339),
.B2(n_439),
.Y(n_587)
);

AOI221xp5_ASAP7_75t_L g588 ( 
.A1(n_559),
.A2(n_521),
.B1(n_531),
.B2(n_557),
.C(n_573),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_558),
.B(n_572),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_555),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_556),
.Y(n_591)
);

OAI21x1_ASAP7_75t_L g592 ( 
.A1(n_556),
.A2(n_571),
.B(n_554),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_564),
.Y(n_593)
);

OAI33xp33_ASAP7_75t_L g594 ( 
.A1(n_578),
.A2(n_576),
.A3(n_580),
.B1(n_566),
.B2(n_582),
.B3(n_583),
.Y(n_594)
);

AOI221xp5_ASAP7_75t_L g595 ( 
.A1(n_558),
.A2(n_574),
.B1(n_587),
.B2(n_560),
.C(n_563),
.Y(n_595)
);

NAND3xp33_ASAP7_75t_L g596 ( 
.A(n_586),
.B(n_576),
.C(n_577),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_562),
.B(n_566),
.Y(n_597)
);

AOI322xp5_ASAP7_75t_L g598 ( 
.A1(n_565),
.A2(n_551),
.A3(n_569),
.B1(n_561),
.B2(n_562),
.C1(n_579),
.C2(n_575),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_585),
.Y(n_599)
);

AOI221xp5_ASAP7_75t_SL g600 ( 
.A1(n_574),
.A2(n_568),
.B1(n_577),
.B2(n_578),
.C(n_549),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_580),
.B(n_553),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_565),
.A2(n_553),
.B1(n_552),
.B2(n_584),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g603 ( 
.A(n_550),
.B(n_552),
.C(n_584),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_564),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_581),
.A2(n_582),
.B1(n_555),
.B2(n_585),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_R g606 ( 
.A(n_555),
.B(n_564),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_567),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_555),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_567),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_598),
.A2(n_581),
.B(n_554),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_604),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_604),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_597),
.B(n_581),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_597),
.B(n_581),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_598),
.A2(n_602),
.B(n_588),
.Y(n_615)
);

NAND4xp25_ASAP7_75t_L g616 ( 
.A(n_600),
.B(n_567),
.C(n_570),
.D(n_550),
.Y(n_616)
);

AOI33xp33_ASAP7_75t_L g617 ( 
.A1(n_595),
.A2(n_550),
.A3(n_570),
.B1(n_605),
.B2(n_608),
.B3(n_591),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_601),
.B(n_589),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_589),
.B(n_570),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_601),
.B(n_550),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_606),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_600),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_599),
.Y(n_623)
);

OAI33xp33_ASAP7_75t_L g624 ( 
.A1(n_622),
.A2(n_618),
.A3(n_613),
.B1(n_616),
.B2(n_596),
.B3(n_615),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_619),
.B(n_596),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_611),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_623),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_620),
.B(n_591),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_621),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_614),
.B(n_591),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_614),
.B(n_605),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_627),
.B(n_621),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_626),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_624),
.A2(n_615),
.B1(n_594),
.B2(n_620),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_626),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_629),
.A2(n_599),
.B1(n_619),
.B2(n_625),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_631),
.B(n_617),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_629),
.A2(n_603),
.B(n_610),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_625),
.A2(n_603),
.B1(n_608),
.B2(n_616),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_633),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_638),
.A2(n_611),
.B(n_593),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_632),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_636),
.B(n_631),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_R g644 ( 
.A(n_637),
.B(n_628),
.Y(n_644)
);

NOR2xp67_ASAP7_75t_L g645 ( 
.A(n_639),
.B(n_628),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_643),
.B(n_634),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_644),
.A2(n_635),
.B1(n_590),
.B2(n_630),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_641),
.A2(n_628),
.B(n_630),
.Y(n_648)
);

AO22x2_ASAP7_75t_L g649 ( 
.A1(n_642),
.A2(n_628),
.B1(n_612),
.B2(n_590),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_642),
.Y(n_650)
);

XOR2xp5_ASAP7_75t_L g651 ( 
.A(n_640),
.B(n_590),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_649),
.B(n_645),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_646),
.B(n_612),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_650),
.A2(n_648),
.B(n_647),
.Y(n_654)
);

OA22x2_ASAP7_75t_SL g655 ( 
.A1(n_651),
.A2(n_644),
.B1(n_604),
.B2(n_607),
.Y(n_655)
);

NAND4xp25_ASAP7_75t_L g656 ( 
.A(n_654),
.B(n_590),
.C(n_609),
.D(n_593),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_652),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_653),
.B(n_592),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_657),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_659),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_660),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_661),
.Y(n_662)
);

INVxp67_ASAP7_75t_SL g663 ( 
.A(n_661),
.Y(n_663)
);

AOI322xp5_ASAP7_75t_L g664 ( 
.A1(n_663),
.A2(n_656),
.A3(n_658),
.B1(n_655),
.B2(n_607),
.C1(n_609),
.C2(n_592),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_664),
.A2(n_662),
.B(n_607),
.Y(n_665)
);


endmodule