module fake_jpeg_3832_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_38),
.Y(n_48)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_28),
.B1(n_31),
.B2(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_41),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_2),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_3),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_28),
.B1(n_19),
.B2(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_42),
.A2(n_60),
.B1(n_32),
.B2(n_24),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_17),
.B(n_30),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_49),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_47),
.B1(n_34),
.B2(n_38),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_30),
.C(n_17),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_55),
.Y(n_62)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_21),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_19),
.B1(n_22),
.B2(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_57),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_39),
.B(n_34),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_69),
.B(n_56),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_75),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_32),
.B1(n_33),
.B2(n_24),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_82),
.B1(n_48),
.B2(n_51),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_43),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_32),
.B1(n_36),
.B2(n_5),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_76),
.A2(n_60),
.B1(n_47),
.B2(n_45),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_49),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_27),
.B1(n_18),
.B2(n_25),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_61),
.Y(n_94)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_46),
.A2(n_27),
.B1(n_29),
.B2(n_23),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_85),
.B(n_88),
.Y(n_115)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_64),
.B(n_50),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_92),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_51),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_48),
.C(n_53),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_67),
.C(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_49),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_97),
.Y(n_121)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_101),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_3),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_107),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_97),
.C(n_12),
.Y(n_141)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_74),
.B1(n_73),
.B2(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_112),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_63),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_90),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_103),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_59),
.B1(n_36),
.B2(n_71),
.Y(n_112)
);

AOI22x1_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_36),
.B1(n_50),
.B2(n_43),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_120),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_84),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_77),
.B(n_4),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_70),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_134),
.C(n_135),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_SL g128 ( 
.A1(n_116),
.A2(n_88),
.A3(n_91),
.B1(n_96),
.B2(n_92),
.C1(n_83),
.C2(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_98),
.B(n_89),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_140),
.B(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_139),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_50),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_50),
.Y(n_135)
);

BUFx6f_ASAP7_75t_SL g136 ( 
.A(n_114),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_59),
.A3(n_43),
.B1(n_86),
.B2(n_75),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_75),
.Y(n_142)
);

OAI21x1_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_122),
.B(n_112),
.Y(n_143)
);

NOR2xp67_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_131),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_156),
.B(n_142),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_115),
.B1(n_119),
.B2(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_115),
.B1(n_124),
.B2(n_106),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_155),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_118),
.B1(n_114),
.B2(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_118),
.B(n_123),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_132),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_66),
.B1(n_104),
.B2(n_6),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_167),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_162),
.B(n_146),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_127),
.B(n_135),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_163),
.A2(n_170),
.B1(n_12),
.B2(n_14),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_134),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_165),
.B(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_148),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_166),
.A2(n_169),
.B(n_147),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_141),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_136),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_172),
.B(n_177),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_144),
.B(n_152),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_173),
.B(n_175),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_151),
.B1(n_157),
.B2(n_156),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_157),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_178),
.Y(n_186)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_165),
.B(n_164),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_13),
.B(n_14),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_158),
.B1(n_170),
.B2(n_167),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_188),
.B1(n_8),
.B2(n_9),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_7),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_180),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_176),
.A2(n_104),
.B1(n_66),
.B2(n_13),
.Y(n_188)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_174),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_193),
.B1(n_186),
.B2(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_194),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_183),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_104),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_8),
.B(n_11),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_194),
.C(n_181),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_195),
.B1(n_196),
.B2(n_8),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_184),
.C(n_9),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);


endmodule