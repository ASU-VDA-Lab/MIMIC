module fake_jpeg_16483_n_108 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_22),
.B(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_0),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_52),
.Y(n_61)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx5_ASAP7_75t_SL g57 ( 
.A(n_53),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_44),
.B1(n_39),
.B2(n_35),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_55),
.B1(n_38),
.B2(n_41),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_44),
.B1(n_39),
.B2(n_35),
.Y(n_55)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_41),
.B(n_42),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_76),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_78),
.C(n_4),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_16),
.B1(n_30),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_73),
.B1(n_59),
.B2(n_7),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_15),
.B1(n_28),
.B2(n_26),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_1),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_1),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_2),
.C(n_4),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_58),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_2),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_90),
.B1(n_6),
.B2(n_32),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_87),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_89),
.B1(n_6),
.B2(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_5),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_74),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_77),
.C(n_67),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_95),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_101),
.B(n_98),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_93),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_98),
.B(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_80),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_90),
.A3(n_89),
.B1(n_96),
.B2(n_81),
.C1(n_19),
.C2(n_21),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_10),
.Y(n_107)
);

AOI221xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.C(n_24),
.Y(n_108)
);


endmodule