module fake_jpeg_12268_n_27 (n_3, n_2, n_1, n_0, n_4, n_5, n_27);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_27;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_2),
.Y(n_6)
);

INVx5_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_4),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

MAJx2_ASAP7_75t_L g11 ( 
.A(n_6),
.B(n_5),
.C(n_1),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_14),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_8),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_13),
.A2(n_8),
.B(n_9),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_9),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_19),
.B(n_2),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_21),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_7),
.B(n_9),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_18),
.Y(n_24)
);

OAI21x1_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_16),
.B(n_21),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_26),
.C(n_23),
.Y(n_27)
);

AOI322xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_3),
.A3(n_4),
.B1(n_7),
.B2(n_9),
.C1(n_16),
.C2(n_22),
.Y(n_26)
);


endmodule