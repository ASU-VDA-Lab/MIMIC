module fake_jpeg_27283_n_83 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_51),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_1),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_55),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_44),
.B(n_46),
.C(n_39),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_10),
.B(n_11),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_45),
.B1(n_38),
.B2(n_8),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_62),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_12),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_13),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.C(n_64),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_72),
.Y(n_74)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_73),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_73),
.B1(n_63),
.B2(n_56),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_74),
.B(n_63),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_60),
.B1(n_59),
.B2(n_20),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_24),
.Y(n_80)
);

AOI322xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_26),
.A3(n_28),
.B1(n_29),
.B2(n_31),
.C1(n_32),
.C2(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_34),
.Y(n_82)
);

BUFx24_ASAP7_75t_SL g83 ( 
.A(n_82),
.Y(n_83)
);


endmodule