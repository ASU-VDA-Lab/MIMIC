module fake_jpeg_1743_n_110 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_35),
.B1(n_32),
.B2(n_38),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_47),
.B1(n_54),
.B2(n_36),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_38),
.B1(n_30),
.B2(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_39),
.B1(n_29),
.B2(n_37),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_36),
.B1(n_33),
.B2(n_3),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_36),
.B1(n_37),
.B2(n_33),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_58),
.B1(n_53),
.B2(n_6),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_63),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_54),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_62),
.Y(n_65)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_4),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_5),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_52),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_69),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_51),
.B(n_50),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_53),
.C(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_18),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_74),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_70),
.B1(n_68),
.B2(n_74),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_SL g96 ( 
.A1(n_76),
.A2(n_79),
.B(n_20),
.Y(n_96)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_86),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_55),
.B(n_60),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_19),
.C(n_26),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_84),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_5),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_81),
.C(n_70),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_14),
.C(n_21),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_7),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_7),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_16),
.B(n_23),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_8),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_96),
.C(n_22),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_96),
.B1(n_28),
.B2(n_87),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.Y(n_102)
);

AOI221xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_100),
.B1(n_88),
.B2(n_97),
.C(n_93),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_98),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_89),
.B(n_102),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_8),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_10),
.B(n_11),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_10),
.Y(n_110)
);


endmodule