module fake_jpeg_30423_n_140 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_11),
.B(n_6),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_62),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_58),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_53),
.B(n_47),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_48),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_76),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_2),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_49),
.B1(n_56),
.B2(n_54),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_62),
.B1(n_59),
.B2(n_51),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_1),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_3),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_73),
.B1(n_79),
.B2(n_80),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_95),
.B1(n_9),
.B2(n_10),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_2),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_27),
.B(n_42),
.C(n_41),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_3),
.B(n_4),
.Y(n_100)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_43),
.B1(n_25),
.B2(n_26),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_4),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_104),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_5),
.B(n_8),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_117)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_9),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_10),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_111),
.Y(n_121)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_40),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_95),
.C(n_92),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_115),
.C(n_96),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_14),
.C(n_16),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_119),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_29),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_30),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_127),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_100),
.B(n_105),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_129),
.B(n_31),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_104),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_121),
.B1(n_120),
.B2(n_123),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_97),
.B(n_32),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_130),
.B(n_132),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_124),
.B1(n_116),
.B2(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.C(n_133),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_33),
.B(n_35),
.Y(n_138)
);

AOI221xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.C(n_39),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_97),
.Y(n_140)
);


endmodule