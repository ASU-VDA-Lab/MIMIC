module fake_jpeg_16407_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_7),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_60),
.Y(n_93)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_16),
.B(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_63),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_66),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_68),
.Y(n_117)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_70),
.Y(n_120)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_73),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_26),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_35),
.Y(n_98)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_77),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_78),
.Y(n_89)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_30),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_41),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_40),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_81),
.Y(n_136)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_39),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_39),
.C(n_41),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_74),
.C(n_77),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_29),
.B1(n_33),
.B2(n_42),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_90),
.A2(n_91),
.B1(n_103),
.B2(n_128),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_35),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_95),
.B(n_104),
.Y(n_156)
);

CKINVDCx12_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_98),
.B(n_13),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_61),
.A2(n_42),
.B1(n_25),
.B2(n_34),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_70),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_52),
.Y(n_112)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_55),
.A2(n_32),
.B1(n_30),
.B2(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_130),
.B1(n_131),
.B2(n_12),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_54),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_63),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_26),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_134),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_68),
.A2(n_49),
.B1(n_57),
.B2(n_83),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_60),
.A2(n_34),
.B1(n_31),
.B2(n_27),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_64),
.A2(n_27),
.B1(n_25),
.B2(n_22),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_81),
.A2(n_22),
.B1(n_39),
.B2(n_3),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_13),
.B1(n_5),
.B2(n_6),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_82),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_69),
.B(n_0),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_72),
.B(n_1),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_110),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_152),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_47),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_141),
.B(n_149),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_145),
.B(n_185),
.Y(n_217)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_65),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_155),
.Y(n_197)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_157),
.B(n_158),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_136),
.B1(n_111),
.B2(n_94),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_1),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_167),
.Y(n_200)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_163),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_78),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_165),
.B(n_171),
.Y(n_192)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_169),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_1),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_172),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_11),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

BUFx12_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_1),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_179),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_96),
.B(n_102),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_176),
.B(n_177),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_99),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_116),
.A2(n_14),
.B1(n_15),
.B2(n_114),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_178),
.A2(n_181),
.B1(n_116),
.B2(n_121),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_125),
.B(n_14),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_131),
.B(n_15),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_182),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_129),
.A2(n_121),
.B1(n_94),
.B2(n_118),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_113),
.B(n_85),
.Y(n_182)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_183),
.B(n_184),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_88),
.B(n_126),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_143),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_207),
.C(n_164),
.Y(n_237)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_136),
.C(n_93),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_190),
.B(n_193),
.Y(n_243)
);

NOR2x1_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_122),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_195),
.A2(n_183),
.B1(n_150),
.B2(n_148),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_141),
.A2(n_84),
.B(n_117),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_196),
.A2(n_164),
.B(n_199),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_208),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_105),
.C(n_101),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_139),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_144),
.A2(n_132),
.B1(n_105),
.B2(n_89),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_209),
.A2(n_212),
.B1(n_214),
.B2(n_221),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_146),
.A2(n_157),
.B1(n_167),
.B2(n_161),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_175),
.A2(n_179),
.B1(n_185),
.B2(n_147),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_149),
.B(n_100),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_219),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_100),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_162),
.A2(n_132),
.B1(n_108),
.B2(n_89),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_147),
.B1(n_138),
.B2(n_154),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_222),
.A2(n_231),
.B1(n_245),
.B2(n_198),
.Y(n_268)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_151),
.B(n_173),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_223),
.A2(n_225),
.B(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_163),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_187),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_227),
.Y(n_252)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_217),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_142),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_235),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_142),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_237),
.C(n_248),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_160),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_238),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_240),
.Y(n_269)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_168),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_205),
.Y(n_267)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_244),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_194),
.A2(n_108),
.B1(n_169),
.B2(n_174),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_214),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_211),
.B(n_216),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_215),
.C(n_199),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_201),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_220),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_209),
.B1(n_197),
.B2(n_204),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_251),
.A2(n_272),
.B1(n_245),
.B2(n_231),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_253),
.B(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

OAI32xp33_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_195),
.A3(n_202),
.B1(n_221),
.B2(n_203),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_233),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_186),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_270),
.C(n_222),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_241),
.B(n_203),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_198),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_229),
.B(n_205),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_264),
.B(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_267),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_191),
.C(n_216),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_233),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_236),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_279),
.C(n_287),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_229),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_232),
.C(n_246),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_283),
.B1(n_268),
.B2(n_270),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_224),
.Y(n_282)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_269),
.Y(n_284)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_271),
.Y(n_292)
);

A2O1A1O1Ixp25_ASAP7_75t_L g286 ( 
.A1(n_250),
.A2(n_228),
.B(n_247),
.C(n_248),
.D(n_242),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_251),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_262),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_247),
.C(n_239),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_290),
.C(n_263),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_238),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_302),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_299),
.C(n_300),
.Y(n_314)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_265),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_290),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_250),
.B1(n_265),
.B2(n_255),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_303),
.B1(n_273),
.B2(n_277),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_256),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_263),
.B1(n_255),
.B2(n_259),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_288),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_315),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_304),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_299),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_301),
.B(n_261),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_312),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_293),
.B(n_276),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_282),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_313),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_273),
.Y(n_315)
);

AOI31xp67_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_286),
.A3(n_291),
.B(n_253),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_320),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_315),
.A2(n_285),
.B(n_302),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_321),
.C(n_314),
.Y(n_325)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_322),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_316),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_328),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_305),
.B(n_306),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_252),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_306),
.A3(n_300),
.B1(n_314),
.B2(n_295),
.C1(n_278),
.C2(n_275),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_316),
.B1(n_295),
.B2(n_323),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_331),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_258),
.B(n_272),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_258),
.B(n_328),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_330),
.B(n_329),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_335),
.A2(n_336),
.B1(n_227),
.B2(n_211),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_191),
.Y(n_338)
);


endmodule