module fake_jpeg_25421_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_7),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_18),
.B1(n_33),
.B2(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_18),
.B1(n_33),
.B2(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_33),
.B(n_25),
.C(n_32),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_28),
.B1(n_27),
.B2(n_32),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_19),
.Y(n_79)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_20),
.C(n_26),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_35),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_65),
.B(n_69),
.Y(n_92)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_42),
.B(n_27),
.C(n_30),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_79),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_18),
.B1(n_33),
.B2(n_32),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_0),
.B(n_1),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_16),
.B(n_31),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_18),
.B1(n_21),
.B2(n_31),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_29),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_87),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_21),
.B1(n_16),
.B2(n_31),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_19),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_21),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_52),
.B(n_19),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_61),
.Y(n_111)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_56),
.B(n_40),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_93),
.Y(n_144)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_91),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_112),
.B(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_65),
.A2(n_27),
.B(n_30),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_65),
.A2(n_30),
.B(n_29),
.Y(n_114)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_89),
.C(n_82),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_43),
.C(n_41),
.Y(n_146)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_86),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_124),
.B(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_79),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_69),
.C(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_127),
.B(n_135),
.Y(n_175)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_72),
.B1(n_47),
.B2(n_51),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_129),
.A2(n_138),
.B1(n_140),
.B2(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_90),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_134),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_66),
.B1(n_80),
.B2(n_88),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_69),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_64),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_136),
.A2(n_149),
.B(n_107),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_141),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_55),
.B1(n_51),
.B2(n_57),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_105),
.B(n_16),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_139),
.B(n_142),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_73),
.B1(n_84),
.B2(n_83),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_92),
.B(n_78),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_100),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_92),
.B(n_84),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_101),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_147),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_81),
.Y(n_147)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_119),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_104),
.A2(n_93),
.B1(n_112),
.B2(n_97),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_150),
.A2(n_174),
.B1(n_106),
.B2(n_24),
.Y(n_210)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_151),
.B(n_152),
.Y(n_206)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_93),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_158),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_156),
.Y(n_208)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_164),
.B1(n_179),
.B2(n_129),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_35),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_163),
.A2(n_172),
.B(n_178),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_99),
.B1(n_88),
.B2(n_80),
.Y(n_164)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_43),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_180),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_177),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_131),
.B(n_29),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_181),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_88),
.B1(n_80),
.B2(n_24),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_95),
.B(n_94),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_182),
.B(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_135),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_20),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_46),
.B1(n_50),
.B2(n_38),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_120),
.B(n_54),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_139),
.B(n_66),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_134),
.B(n_40),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_194),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_195),
.B1(n_197),
.B2(n_204),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_167),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_125),
.C(n_136),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_200),
.C(n_178),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_140),
.B(n_143),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_190),
.B(n_192),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_143),
.B(n_138),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_121),
.B(n_1),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_177),
.B1(n_164),
.B2(n_179),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_157),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_196),
.B(n_209),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_121),
.B1(n_123),
.B2(n_22),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_123),
.Y(n_199)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_43),
.C(n_116),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_211),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_0),
.B(n_2),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_202),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_180),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_203),
.B(n_116),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_0),
.B(n_2),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_210),
.B1(n_194),
.B2(n_154),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_106),
.B(n_43),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_159),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_215),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_211),
.B(n_212),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_222),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_200),
.C(n_198),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_216),
.C(n_235),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_150),
.B1(n_178),
.B2(n_167),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_225),
.B1(n_233),
.B2(n_210),
.Y(n_243)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_229),
.Y(n_258)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_182),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_188),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_166),
.Y(n_224)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_186),
.A2(n_152),
.B1(n_154),
.B2(n_165),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_204),
.B1(n_192),
.B2(n_187),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_208),
.B(n_166),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_234),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_26),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_201),
.A2(n_23),
.B1(n_22),
.B2(n_24),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_209),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_26),
.Y(n_237)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_197),
.B1(n_191),
.B2(n_190),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_238),
.A2(n_213),
.B1(n_230),
.B2(n_233),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_242),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_193),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_243),
.A2(n_17),
.B1(n_26),
.B2(n_3),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_244),
.A2(n_218),
.B1(n_238),
.B2(n_248),
.Y(n_265)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_252),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_183),
.Y(n_247)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_255),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_203),
.C(n_193),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_222),
.C(n_236),
.Y(n_264)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_220),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_254),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_202),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_218),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_219),
.Y(n_261)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_253),
.A2(n_227),
.B(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_249),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_266),
.B(n_242),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_213),
.B1(n_187),
.B2(n_183),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_273),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_205),
.B1(n_23),
.B2(n_22),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_23),
.B1(n_116),
.B2(n_26),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_258),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_259),
.C(n_266),
.Y(n_291)
);

NOR3xp33_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_256),
.C(n_251),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_284),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_12),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_240),
.Y(n_281)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

AO221x1_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_257),
.B1(n_17),
.B2(n_4),
.C(n_6),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_283),
.A2(n_12),
.B1(n_15),
.B2(n_4),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_256),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_264),
.C(n_259),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_287),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_17),
.C(n_40),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_268),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_292),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_291),
.B(n_293),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_272),
.C(n_270),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_273),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_269),
.B1(n_17),
.B2(n_4),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_297),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_0),
.B1(n_3),
.B2(n_6),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_286),
.B(n_12),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_301),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_17),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_279),
.B(n_280),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_304),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_277),
.A3(n_282),
.B1(n_287),
.B2(n_9),
.C1(n_11),
.C2(n_13),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_11),
.C(n_15),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_309),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_297),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_6),
.C(n_9),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_313),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_299),
.C(n_11),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_306),
.B(n_13),
.Y(n_314)
);

AOI21xp33_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_316),
.B(n_317),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_14),
.C(n_3),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_304),
.Y(n_317)
);

O2A1O1Ixp33_ASAP7_75t_SL g318 ( 
.A1(n_311),
.A2(n_14),
.B(n_40),
.C(n_315),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_319),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_320),
.C(n_14),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_40),
.Y(n_324)
);


endmodule