module fake_netlist_1_8313_n_685 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_166, n_162, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_685);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_685;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_424;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_406;
wire n_395;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_57), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_100), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_112), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_21), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_62), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_88), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_126), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_93), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_146), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_139), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_122), .Y(n_186) );
INVxp67_ASAP7_75t_L g187 ( .A(n_37), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_171), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_111), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_121), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_169), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_41), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_59), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_84), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_132), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_160), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_90), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_35), .B(n_65), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_66), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_149), .B(n_172), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_119), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_0), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_7), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_20), .Y(n_204) );
INVxp33_ASAP7_75t_L g205 ( .A(n_23), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_91), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_42), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_162), .Y(n_208) );
INVxp67_ASAP7_75t_SL g209 ( .A(n_48), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_71), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_136), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_7), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_67), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_148), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_156), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_140), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_80), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_107), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_28), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_125), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_19), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_143), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_174), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_166), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_52), .Y(n_225) );
BUFx3_ASAP7_75t_L g226 ( .A(n_69), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_18), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_163), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_141), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_131), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_158), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_65), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_50), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_118), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_99), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_159), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_3), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_110), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_134), .Y(n_239) );
INVxp67_ASAP7_75t_SL g240 ( .A(n_101), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_34), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_109), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_14), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_4), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_68), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_44), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_120), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_108), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_98), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_51), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_138), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_161), .Y(n_252) );
INVxp33_ASAP7_75t_SL g253 ( .A(n_113), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_63), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_102), .Y(n_255) );
CKINVDCx16_ASAP7_75t_R g256 ( .A(n_117), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_144), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_79), .Y(n_258) );
BUFx5_ASAP7_75t_L g259 ( .A(n_152), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_147), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_97), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_35), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_133), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_94), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_114), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_145), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_74), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_137), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_135), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_12), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_33), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_85), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_68), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_11), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_53), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_226), .B(n_0), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_259), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_259), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_202), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_202), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_259), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_178), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_259), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_203), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_259), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_205), .B(n_1), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_259), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_203), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_207), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_207), .Y(n_290) );
OAI22xp5_ASAP7_75t_SL g291 ( .A1(n_175), .A2(n_5), .B1(n_2), .B2(n_4), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_226), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_244), .Y(n_293) );
BUFx8_ASAP7_75t_L g294 ( .A(n_251), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_186), .Y(n_295) );
AND2x6_ASAP7_75t_L g296 ( .A(n_178), .B(n_72), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_205), .B(n_5), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_244), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_176), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_186), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_181), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_183), .Y(n_302) );
OAI22xp5_ASAP7_75t_SL g303 ( .A1(n_175), .A2(n_9), .B1(n_6), .B2(n_8), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_185), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_187), .B(n_8), .Y(n_305) );
NAND2xp33_ASAP7_75t_R g306 ( .A(n_253), .B(n_73), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_276), .B(n_179), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_282), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_276), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_294), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_276), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_282), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_294), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_297), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_286), .B(n_180), .Y(n_316) );
INVx8_ASAP7_75t_L g317 ( .A(n_296), .Y(n_317) );
INVx5_ASAP7_75t_L g318 ( .A(n_296), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_299), .B(n_253), .Y(n_319) );
OR2x6_ASAP7_75t_L g320 ( .A(n_291), .B(n_198), .Y(n_320) );
INVx8_ASAP7_75t_L g321 ( .A(n_296), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_301), .B(n_228), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_301), .B(n_256), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_282), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_292), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_286), .B(n_192), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_302), .B(n_206), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_296), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_302), .B(n_193), .Y(n_329) );
INVx4_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_304), .B(n_199), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_292), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_305), .A2(n_182), .B1(n_214), .B2(n_195), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_295), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_294), .Y(n_335) );
BUFx10_ASAP7_75t_L g336 ( .A(n_296), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_279), .B(n_199), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_279), .B(n_212), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_280), .B(n_213), .Y(n_339) );
NOR2xp33_ASAP7_75t_R g340 ( .A(n_311), .B(n_306), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_315), .B(n_177), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_314), .B(n_238), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_328), .B(n_190), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_319), .B(n_277), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_337), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_323), .B(n_196), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_320), .A2(n_257), .B1(n_238), .B2(n_303), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_337), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_334), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_322), .B(n_196), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_334), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_335), .B(n_280), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_308), .B(n_277), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_316), .B(n_222), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_338), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_338), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_316), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_339), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_326), .B(n_284), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_333), .B(n_219), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_308), .B(n_277), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_325), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_317), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_326), .A2(n_227), .B1(n_246), .B2(n_245), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_326), .B(n_258), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_331), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_332), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_329), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_313), .Y(n_370) );
OR2x6_ASAP7_75t_L g371 ( .A(n_320), .B(n_221), .Y(n_371) );
AOI21x1_ASAP7_75t_L g372 ( .A1(n_310), .A2(n_281), .B(n_278), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_312), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_330), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_327), .Y(n_375) );
INVx8_ASAP7_75t_L g376 ( .A(n_317), .Y(n_376) );
INVx4_ASAP7_75t_L g377 ( .A(n_321), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_321), .A2(n_270), .B1(n_275), .B2(n_271), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_318), .B(n_268), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_313), .Y(n_380) );
INVx5_ASAP7_75t_L g381 ( .A(n_321), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_318), .B(n_278), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_318), .B(n_278), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_318), .B(n_281), .Y(n_384) );
OR2x6_ASAP7_75t_L g385 ( .A(n_307), .B(n_225), .Y(n_385) );
OAI22xp5_ASAP7_75t_SL g386 ( .A1(n_318), .A2(n_237), .B1(n_241), .B2(n_204), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_336), .B(n_281), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_336), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_307), .B(n_283), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_309), .B(n_283), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_309), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_367), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_355), .B(n_356), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_352), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_342), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_344), .A2(n_287), .B(n_285), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
OA22x2_ASAP7_75t_L g398 ( .A1(n_360), .A2(n_209), .B1(n_233), .B2(n_232), .Y(n_398) );
INVx5_ASAP7_75t_L g399 ( .A(n_385), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_369), .Y(n_400) );
NAND2x1p5_ASAP7_75t_L g401 ( .A(n_381), .B(n_293), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_381), .B(n_184), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_387), .A2(n_287), .B(n_240), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_345), .B(n_300), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_348), .A2(n_243), .B1(n_254), .B2(n_250), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_373), .B(n_262), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_358), .Y(n_407) );
A2O1A1Ixp33_ASAP7_75t_L g408 ( .A1(n_363), .A2(n_274), .B(n_273), .C(n_284), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_349), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_351), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_385), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_387), .A2(n_189), .B(n_188), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_359), .A2(n_289), .B1(n_298), .B2(n_290), .C(n_288), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_353), .A2(n_194), .B(n_191), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_341), .B(n_296), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_347), .B(n_293), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_353), .B(n_197), .Y(n_418) );
INVx5_ASAP7_75t_L g419 ( .A(n_385), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_368), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_365), .B(n_10), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_361), .B(n_201), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_389), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_386), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_340), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_375), .B(n_208), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_377), .B(n_211), .Y(n_427) );
OA22x2_ASAP7_75t_L g428 ( .A1(n_347), .A2(n_217), .B1(n_218), .B2(n_216), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_354), .B(n_220), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_390), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_L g431 ( .A1(n_350), .A2(n_230), .B(n_231), .C(n_224), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_366), .B(n_234), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_346), .B(n_242), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_364), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_378), .B(n_252), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_390), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_380), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_382), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_374), .B(n_255), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g440 ( .A(n_343), .B(n_215), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_382), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_370), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_383), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_383), .A2(n_261), .B(n_260), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_379), .A2(n_282), .B1(n_266), .B2(n_267), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_384), .B(n_264), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_391), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_388), .B(n_269), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_352), .Y(n_449) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_376), .Y(n_450) );
BUFx8_ASAP7_75t_SL g451 ( .A(n_371), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_357), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_372), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_367), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_372), .Y(n_455) );
OR2x6_ASAP7_75t_L g456 ( .A(n_371), .B(n_210), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_372), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_367), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_357), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_393), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_399), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_393), .Y(n_462) );
OAI21x1_ASAP7_75t_L g463 ( .A1(n_453), .A2(n_235), .B(n_229), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_392), .B(n_235), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_396), .A2(n_247), .B(n_239), .Y(n_465) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_455), .A2(n_248), .B(n_247), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_396), .A2(n_249), .B(n_248), .Y(n_467) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_457), .A2(n_265), .B(n_263), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_404), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_399), .Y(n_470) );
AO31x2_ASAP7_75t_L g471 ( .A1(n_415), .A2(n_265), .A3(n_272), .B(n_200), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_428), .A2(n_236), .B1(n_223), .B2(n_272), .Y(n_472) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_403), .A2(n_236), .B(n_223), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_454), .B(n_13), .Y(n_474) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_434), .Y(n_475) );
AO31x2_ASAP7_75t_L g476 ( .A1(n_415), .A2(n_324), .A3(n_14), .B(n_13), .Y(n_476) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_444), .A2(n_413), .B(n_416), .Y(n_477) );
OAI21x1_ASAP7_75t_L g478 ( .A1(n_444), .A2(n_324), .B(n_75), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_420), .Y(n_479) );
AO32x2_ASAP7_75t_L g480 ( .A1(n_405), .A2(n_15), .A3(n_16), .B1(n_17), .B2(n_18), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_428), .A2(n_16), .B1(n_19), .B2(n_20), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_398), .A2(n_22), .B1(n_23), .B2(n_24), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_431), .B(n_22), .C(n_25), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_423), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_458), .Y(n_485) );
OAI21x1_ASAP7_75t_L g486 ( .A1(n_447), .A2(n_77), .B(n_76), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_399), .Y(n_487) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_394), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_430), .Y(n_489) );
OAI21x1_ASAP7_75t_L g490 ( .A1(n_440), .A2(n_81), .B(n_78), .Y(n_490) );
OAI21x1_ASAP7_75t_SL g491 ( .A1(n_426), .A2(n_26), .B(n_27), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_436), .Y(n_492) );
BUFx2_ASAP7_75t_R g493 ( .A(n_451), .Y(n_493) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_426), .A2(n_83), .B(n_82), .Y(n_494) );
OAI21x1_ASAP7_75t_L g495 ( .A1(n_440), .A2(n_87), .B(n_86), .Y(n_495) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_429), .A2(n_92), .B(n_89), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_400), .B(n_29), .Y(n_497) );
INVx5_ASAP7_75t_L g498 ( .A(n_450), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_397), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_407), .B(n_29), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_443), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_406), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_419), .B(n_30), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_406), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_437), .Y(n_505) );
NAND2x1p5_ASAP7_75t_L g506 ( .A(n_419), .B(n_30), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_398), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_507) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_446), .A2(n_96), .B(n_95), .Y(n_508) );
AOI222xp33_ASAP7_75t_L g509 ( .A1(n_424), .A2(n_36), .B1(n_37), .B2(n_38), .C1(n_39), .C2(n_40), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_438), .Y(n_510) );
BUFx2_ASAP7_75t_SL g511 ( .A(n_419), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_409), .Y(n_512) );
OAI22xp33_ASAP7_75t_L g513 ( .A1(n_456), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_410), .Y(n_514) );
INVx6_ASAP7_75t_L g515 ( .A(n_419), .Y(n_515) );
OAI21x1_ASAP7_75t_L g516 ( .A1(n_401), .A2(n_123), .B(n_173), .Y(n_516) );
OAI21x1_ASAP7_75t_L g517 ( .A1(n_442), .A2(n_124), .B(n_170), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_418), .A2(n_43), .B1(n_45), .B2(n_46), .Y(n_518) );
OAI211xp5_ASAP7_75t_L g519 ( .A1(n_414), .A2(n_45), .B(n_47), .C(n_49), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_452), .Y(n_520) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_429), .A2(n_127), .B(n_168), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_433), .A2(n_53), .B(n_54), .C(n_55), .Y(n_522) );
INVxp67_ASAP7_75t_L g523 ( .A(n_449), .Y(n_523) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_434), .Y(n_524) );
OAI22xp33_ASAP7_75t_L g525 ( .A1(n_417), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_525) );
OAI21x1_ASAP7_75t_L g526 ( .A1(n_402), .A2(n_128), .B(n_167), .Y(n_526) );
OAI21x1_ASAP7_75t_L g527 ( .A1(n_445), .A2(n_129), .B(n_165), .Y(n_527) );
INVx4_ASAP7_75t_SL g528 ( .A(n_434), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_421), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_529) );
AO31x2_ASAP7_75t_L g530 ( .A1(n_408), .A2(n_60), .A3(n_61), .B(n_62), .Y(n_530) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_432), .A2(n_130), .B(n_164), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_459), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_441), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g534 ( .A(n_412), .B(n_64), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_422), .B(n_66), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_435), .A2(n_67), .B(n_70), .Y(n_536) );
BUFx2_ASAP7_75t_L g537 ( .A(n_395), .Y(n_537) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_439), .A2(n_103), .B(n_104), .Y(n_538) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_448), .A2(n_105), .B(n_106), .Y(n_539) );
AND2x6_ASAP7_75t_SL g540 ( .A(n_493), .B(n_427), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_485), .B(n_425), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_498), .B(n_411), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_479), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_533), .Y(n_544) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_498), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_483), .B(n_115), .C(n_116), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_465), .A2(n_467), .B(n_535), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_497), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_497), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_498), .B(n_142), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_500), .Y(n_551) );
AOI222xp33_ASAP7_75t_L g552 ( .A1(n_525), .A2(n_150), .B1(n_153), .B2(n_154), .C1(n_155), .C2(n_157), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_500), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_465), .A2(n_467), .B(n_477), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_510), .B(n_484), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_488), .A2(n_506), .B1(n_472), .B2(n_534), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_506), .A2(n_472), .B1(n_507), .B2(n_482), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_474), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_489), .B(n_492), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_499), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_482), .A2(n_507), .B1(n_481), .B2(n_529), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_481), .A2(n_529), .B1(n_513), .B2(n_518), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_501), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_477), .A2(n_473), .B(n_463), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_505), .B(n_512), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_520), .Y(n_566) );
OAI211xp5_ASAP7_75t_L g567 ( .A1(n_509), .A2(n_519), .B(n_522), .C(n_536), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_532), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_464), .A2(n_523), .B1(n_537), .B2(n_461), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_470), .B(n_487), .Y(n_570) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_503), .A2(n_511), .B1(n_491), .B2(n_515), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_514), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_508), .A2(n_494), .B(n_468), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_530), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_480), .B(n_530), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_471), .B(n_530), .Y(n_576) );
OAI211xp5_ASAP7_75t_L g577 ( .A1(n_521), .A2(n_494), .B(n_508), .C(n_468), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_466), .A2(n_524), .B1(n_475), .B2(n_480), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_530), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_476), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_476), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_480), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_478), .A2(n_496), .B(n_531), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_539), .A2(n_538), .B1(n_475), .B2(n_524), .C(n_471), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_528), .B(n_524), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_476), .B(n_471), .Y(n_586) );
AOI22xp5_ASAP7_75t_SL g587 ( .A1(n_528), .A2(n_476), .B1(n_495), .B2(n_490), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_528), .B(n_527), .Y(n_588) );
BUFx3_ASAP7_75t_L g589 ( .A(n_516), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_526), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g591 ( .A1(n_486), .A2(n_504), .B(n_502), .C(n_469), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_517), .B(n_392), .Y(n_592) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_498), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g594 ( .A1(n_465), .A2(n_467), .B(n_396), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_460), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_460), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_460), .B(n_462), .Y(n_597) );
OA21x2_ASAP7_75t_L g598 ( .A1(n_573), .A2(n_584), .B(n_583), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_595), .B(n_596), .Y(n_599) );
NOR2x1_ASAP7_75t_SL g600 ( .A(n_545), .B(n_593), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_566), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_568), .Y(n_602) );
OR2x2_ASAP7_75t_SL g603 ( .A(n_576), .B(n_580), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_570), .B(n_544), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_563), .B(n_597), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_555), .B(n_559), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_543), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_560), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_555), .B(n_559), .Y(n_609) );
INVx3_ASAP7_75t_L g610 ( .A(n_545), .Y(n_610) );
INVx3_ASAP7_75t_L g611 ( .A(n_593), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_565), .B(n_572), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_585), .B(n_593), .Y(n_613) );
OA21x2_ASAP7_75t_L g614 ( .A1(n_564), .A2(n_577), .B(n_554), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_548), .B(n_549), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_551), .B(n_553), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_581), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_558), .B(n_574), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_586), .B(n_575), .Y(n_619) );
BUFx3_ASAP7_75t_L g620 ( .A(n_542), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_579), .B(n_562), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_582), .B(n_561), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_569), .B(n_557), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_541), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_550), .B(n_591), .Y(n_625) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_542), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_547), .B(n_552), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_550), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_557), .B(n_556), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g630 ( .A(n_589), .B(n_587), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_556), .B(n_567), .Y(n_631) );
INVx3_ASAP7_75t_L g632 ( .A(n_592), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_594), .B(n_571), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_594), .B(n_588), .Y(n_634) );
OR2x2_ASAP7_75t_SL g635 ( .A(n_540), .B(n_546), .Y(n_635) );
BUFx2_ASAP7_75t_L g636 ( .A(n_590), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_578), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_628), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_619), .B(n_622), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_622), .B(n_606), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_606), .B(n_609), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_618), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_612), .B(n_633), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_621), .B(n_629), .Y(n_644) );
BUFx3_ASAP7_75t_L g645 ( .A(n_620), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_599), .B(n_605), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_604), .B(n_603), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_617), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_615), .B(n_616), .Y(n_649) );
OR2x6_ASAP7_75t_L g650 ( .A(n_630), .B(n_625), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_631), .B(n_627), .Y(n_651) );
BUFx3_ASAP7_75t_L g652 ( .A(n_620), .Y(n_652) );
AND2x2_ASAP7_75t_SL g653 ( .A(n_623), .B(n_625), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_632), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_632), .Y(n_655) );
AND2x4_ASAP7_75t_L g656 ( .A(n_625), .B(n_634), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_601), .B(n_602), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_607), .B(n_608), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_639), .B(n_637), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_649), .B(n_624), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_640), .B(n_636), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_646), .B(n_626), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_644), .B(n_614), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_647), .B(n_598), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_643), .B(n_598), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_648), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_641), .B(n_613), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_659), .B(n_651), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_661), .B(n_642), .Y(n_669) );
XNOR2xp5_ASAP7_75t_L g670 ( .A(n_660), .B(n_653), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_665), .B(n_656), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_670), .A2(n_650), .B1(n_662), .B2(n_667), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_668), .B(n_663), .Y(n_673) );
XNOR2xp5_ASAP7_75t_L g674 ( .A(n_672), .B(n_635), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_673), .B(n_669), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_674), .A2(n_658), .B1(n_657), .B2(n_671), .C(n_664), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_676), .B(n_675), .Y(n_677) );
NOR3x1_ASAP7_75t_L g678 ( .A(n_677), .B(n_655), .C(n_654), .Y(n_678) );
XNOR2xp5_ASAP7_75t_L g679 ( .A(n_678), .B(n_652), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_679), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_680), .Y(n_681) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_681), .B(n_610), .C(n_611), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_682), .Y(n_683) );
AOI22xp5_ASAP7_75t_SL g684 ( .A1(n_683), .A2(n_645), .B1(n_610), .B2(n_638), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_684), .A2(n_600), .B(n_666), .Y(n_685) );
endmodule