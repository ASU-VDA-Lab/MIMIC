module fake_netlist_1_3242_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
NOR2xp33_ASAP7_75t_L g3 ( .A(n_1), .B(n_2), .Y(n_3) );
CKINVDCx5p33_ASAP7_75t_R g4 ( .A(n_1), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_3), .Y(n_5) );
AOI21xp5_ASAP7_75t_SL g6 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_5), .B(n_4), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
AOI222xp33_ASAP7_75t_SL g9 ( .A1(n_8), .A2(n_5), .B1(n_1), .B2(n_0), .C1(n_2), .C2(n_6), .Y(n_9) );
NOR2x1_ASAP7_75t_L g10 ( .A(n_9), .B(n_7), .Y(n_10) );
OAI21xp5_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_5), .B(n_0), .Y(n_11) );
AO21x2_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_2), .B(n_0), .Y(n_12) );
endmodule