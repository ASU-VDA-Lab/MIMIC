module fake_jpeg_22781_n_348 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_52),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_31),
.B1(n_32),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_53),
.A2(n_80),
.B1(n_81),
.B2(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_66),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_26),
.Y(n_59)
);

OR2x4_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_65),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_22),
.B1(n_32),
.B2(n_31),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_69),
.B(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_33),
.C(n_28),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_31),
.B1(n_32),
.B2(n_22),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_29),
.B1(n_35),
.B2(n_18),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_41),
.A2(n_33),
.B1(n_18),
.B2(n_30),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_79),
.Y(n_90)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_34),
.B1(n_17),
.B2(n_33),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_24),
.B1(n_34),
.B2(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_59),
.B(n_39),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_39),
.C(n_58),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_88),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_83),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_40),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_106),
.B1(n_62),
.B2(n_56),
.Y(n_124)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_94),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_37),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_112),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_42),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_61),
.B(n_30),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_102),
.B(n_103),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_16),
.B(n_37),
.C(n_29),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_24),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_104),
.B(n_119),
.Y(n_148)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_35),
.B1(n_29),
.B2(n_25),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_63),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_107),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_43),
.B1(n_51),
.B2(n_35),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_55),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_111),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_25),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

BUFx24_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_114),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_25),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_113),
.Y(n_142)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_118),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_39),
.Y(n_120)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_35),
.B1(n_29),
.B2(n_16),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_62),
.B1(n_56),
.B2(n_66),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_124),
.B1(n_130),
.B2(n_133),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_85),
.C(n_100),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_84),
.A2(n_86),
.B1(n_88),
.B2(n_103),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_83),
.A2(n_19),
.B(n_16),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_140),
.B(n_119),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_95),
.A2(n_19),
.B1(n_16),
.B2(n_2),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_94),
.B1(n_92),
.B2(n_116),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_111),
.Y(n_163)
);

AOI31xp33_ASAP7_75t_L g143 ( 
.A1(n_95),
.A2(n_19),
.A3(n_16),
.B(n_14),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_143),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_146),
.A2(n_117),
.B1(n_101),
.B2(n_91),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_0),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_148),
.Y(n_159)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_154),
.Y(n_198)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_176),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_93),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_156),
.B(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

O2A1O1Ixp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_130),
.B(n_125),
.C(n_143),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_139),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_163),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_121),
.B1(n_112),
.B2(n_115),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_160),
.A2(n_171),
.B1(n_175),
.B2(n_184),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_161),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_140),
.B(n_131),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_164),
.A2(n_186),
.B(n_126),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_172),
.C(n_180),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_141),
.B(n_139),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_137),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_148),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_173),
.B1(n_183),
.B2(n_134),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_137),
.B(n_93),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_170),
.B(n_177),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_110),
.B1(n_117),
.B2(n_91),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_90),
.C(n_107),
.Y(n_172)
);

AO21x2_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_114),
.B(n_98),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_174),
.A2(n_134),
.B1(n_144),
.B2(n_126),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_123),
.A2(n_114),
.B1(n_101),
.B2(n_118),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_118),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_118),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_178),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_105),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_114),
.C(n_109),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_14),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_182),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_11),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_124),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_3),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_141),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_12),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_189),
.A2(n_138),
.B1(n_4),
.B2(n_5),
.Y(n_245)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_122),
.Y(n_196)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_203),
.Y(n_241)
);

FAx1_ASAP7_75t_SL g232 ( 
.A(n_202),
.B(n_172),
.CI(n_159),
.CON(n_232),
.SN(n_232)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_210),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_219),
.B1(n_168),
.B2(n_180),
.Y(n_225)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_213),
.A2(n_217),
.B(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_156),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_158),
.A2(n_150),
.B1(n_144),
.B2(n_152),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_167),
.B(n_3),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_185),
.B(n_164),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_161),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_221),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_165),
.C(n_166),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_242),
.C(n_202),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_225),
.B(n_232),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_190),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_194),
.A2(n_197),
.B(n_213),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_229),
.A2(n_234),
.B1(n_235),
.B2(n_245),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_162),
.B1(n_183),
.B2(n_170),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_239),
.Y(n_265)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_219),
.A2(n_162),
.B1(n_175),
.B2(n_184),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_205),
.A2(n_175),
.B1(n_186),
.B2(n_176),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_236),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_198),
.B(n_186),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_237),
.B(n_217),
.Y(n_261)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_175),
.C(n_155),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_210),
.A2(n_215),
.B1(n_218),
.B2(n_206),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_216),
.B1(n_206),
.B2(n_204),
.Y(n_260)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_249),
.Y(n_252)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_240),
.B(n_200),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_253),
.B(n_232),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_266),
.C(n_270),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_257),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_195),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_263),
.B1(n_234),
.B2(n_246),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_269),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_188),
.B1(n_189),
.B2(n_201),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_220),
.C(n_192),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_236),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_267),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_192),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_220),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_250),
.A2(n_243),
.B1(n_244),
.B2(n_241),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_273),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_258),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_268),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_235),
.B1(n_247),
.B2(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_277),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_223),
.B1(n_239),
.B2(n_224),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_260),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_251),
.A2(n_245),
.B1(n_248),
.B2(n_227),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_226),
.B1(n_224),
.B2(n_248),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_229),
.B1(n_232),
.B2(n_231),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_253),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_265),
.A2(n_207),
.B1(n_199),
.B2(n_228),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_289),
.B(n_273),
.Y(n_302)
);

XNOR2x2_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_212),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_269),
.B(n_255),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_293),
.B(n_277),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_294),
.A2(n_303),
.B(n_279),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_271),
.B(n_262),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_295),
.A2(n_287),
.B(n_288),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_304),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_191),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_297),
.B(n_300),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_254),
.C(n_266),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_301),
.C(n_306),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_272),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_270),
.C(n_257),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_280),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_191),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_3),
.C(n_4),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_315),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_309),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_279),
.B1(n_291),
.B2(n_287),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_310),
.A2(n_319),
.B1(n_306),
.B2(n_296),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_303),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_274),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_320),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_281),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_286),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_318),
.C(n_3),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_275),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_292),
.B(n_278),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_308),
.A2(n_298),
.B1(n_307),
.B2(n_295),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_317),
.B1(n_313),
.B2(n_315),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_323),
.A2(n_330),
.B(n_4),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_292),
.Y(n_324)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_324),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_321),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_316),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_314),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_313),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_4),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_336),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_334),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_335),
.A2(n_337),
.B(n_330),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_329),
.Y(n_337)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_339),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_325),
.C(n_7),
.Y(n_340)
);

AOI221xp5_ASAP7_75t_L g342 ( 
.A1(n_340),
.A2(n_333),
.B1(n_332),
.B2(n_8),
.C(n_9),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_342),
.A2(n_343),
.B(n_338),
.Y(n_344)
);

AOI322xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C1(n_341),
.C2(n_330),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_10),
.C(n_6),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_7),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_10),
.Y(n_348)
);


endmodule