module fake_netlist_6_206_n_1955 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1955);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1955;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_141),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_22),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_23),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_52),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_125),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_119),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_20),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_135),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_65),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_105),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_146),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_112),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_157),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_63),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_38),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_56),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_2),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_126),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_111),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_9),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_92),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_33),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_151),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_17),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_16),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_72),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_16),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_90),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_117),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_2),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_29),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_54),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_139),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_99),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_38),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_162),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_89),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_19),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_22),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_42),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_175),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_57),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_81),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_21),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_174),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_62),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_71),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_158),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_170),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_56),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_39),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_91),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_115),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_40),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_8),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_53),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_164),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_86),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_66),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_144),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_77),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_177),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_124),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_118),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_94),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_167),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_93),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_21),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_123),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_166),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_101),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_176),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_110),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_107),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_13),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_31),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_19),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_148),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_44),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_88),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_62),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_14),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_73),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_127),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_4),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_13),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_50),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_100),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_44),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_52),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_114),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_78),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_26),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_37),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_17),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_15),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_79),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_11),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_54),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_109),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_149),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_64),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_75),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_43),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_26),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_10),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_76),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_132),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_153),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_63),
.Y(n_300)
);

BUFx2_ASAP7_75t_SL g301 ( 
.A(n_165),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_59),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_102),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_85),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_42),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_57),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_122),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_18),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_4),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_87),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_59),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_121),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_67),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_25),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_6),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_50),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_83),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_49),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_6),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_108),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_154),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_106),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_65),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_104),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_97),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_25),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_46),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_35),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_30),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_129),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_28),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_96),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_43),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_169),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_36),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_37),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_48),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_51),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_30),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_33),
.Y(n_340)
);

INVxp33_ASAP7_75t_R g341 ( 
.A(n_12),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_32),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_69),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_53),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_67),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_178),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_32),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_168),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_24),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_64),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_12),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_46),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_58),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_68),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_41),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_55),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_211),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_265),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_185),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_187),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_188),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_255),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_190),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_211),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_270),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_192),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_211),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_318),
.B(n_0),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_211),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_265),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_211),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_195),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_336),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_211),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_196),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_336),
.B(n_1),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_274),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_222),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_277),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_183),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_222),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_197),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_222),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_222),
.Y(n_384)
);

INVxp33_ASAP7_75t_SL g385 ( 
.A(n_184),
.Y(n_385)
);

INVxp33_ASAP7_75t_SL g386 ( 
.A(n_189),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_222),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_277),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_240),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_222),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_318),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_349),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_198),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_204),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_231),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_205),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_295),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_349),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_349),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_240),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_215),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_240),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_216),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_220),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_343),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_181),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_182),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_221),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_231),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_224),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_181),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_226),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_348),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_233),
.Y(n_418)
);

INVxp33_ASAP7_75t_SL g419 ( 
.A(n_191),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_235),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_343),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_238),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_239),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_251),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_183),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_207),
.B(n_1),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_295),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_266),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_247),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_266),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_248),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_186),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_186),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_250),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_252),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_200),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_200),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_203),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_251),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_203),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_253),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_206),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_256),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_207),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_206),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_208),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_444),
.B(n_209),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_426),
.B(n_332),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_388),
.B(n_332),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_357),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_357),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_444),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_416),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_364),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_388),
.B(n_207),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_444),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_364),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_367),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_367),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_369),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_369),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_371),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_371),
.B(n_209),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_374),
.Y(n_464)
);

OA21x2_ASAP7_75t_L g465 ( 
.A1(n_374),
.A2(n_381),
.B(n_378),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_378),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_381),
.Y(n_467)
);

NOR2x1_ASAP7_75t_L g468 ( 
.A(n_426),
.B(n_243),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_388),
.B(n_390),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_383),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_390),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_389),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_383),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_387),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_392),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_398),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_392),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_393),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_393),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

OR2x6_ASAP7_75t_L g484 ( 
.A(n_368),
.B(n_301),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_394),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_268),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_428),
.B(n_317),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_401),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_401),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_417),
.B(n_243),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_417),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_425),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_425),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_410),
.B(n_268),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_432),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_368),
.B(n_243),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_432),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_436),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_446),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_436),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_437),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_437),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_438),
.A2(n_356),
.B(n_218),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_440),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_440),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_403),
.B(n_259),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_442),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_442),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_415),
.B(n_291),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_400),
.B(n_266),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_445),
.Y(n_517)
);

OA21x2_ASAP7_75t_L g518 ( 
.A1(n_445),
.A2(n_218),
.B(n_208),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_403),
.B(n_259),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_413),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_446),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_405),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_405),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_408),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_515),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_465),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_457),
.Y(n_527)
);

OAI21xp33_ASAP7_75t_SL g528 ( 
.A1(n_499),
.A2(n_439),
.B(n_424),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_448),
.B(n_385),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_471),
.B(n_360),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_448),
.B(n_361),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_448),
.A2(n_434),
.B1(n_435),
.B2(n_429),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_471),
.B(n_363),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_469),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_465),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_501),
.A2(n_373),
.B1(n_370),
.B2(n_358),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_465),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_465),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_483),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_465),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_516),
.B(n_366),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_469),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_469),
.B(n_408),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_469),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_471),
.B(n_372),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_457),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_501),
.A2(n_370),
.B1(n_358),
.B2(n_427),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_453),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_516),
.A2(n_400),
.B1(n_379),
.B2(n_428),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_457),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_453),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_471),
.B(n_409),
.Y(n_554)
);

INVx5_ASAP7_75t_L g555 ( 
.A(n_456),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_494),
.B(n_375),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_501),
.A2(n_391),
.B1(n_227),
.B2(n_230),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_456),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_455),
.B(n_259),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_457),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_483),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_494),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_516),
.B(n_382),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_472),
.B(n_379),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_522),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_456),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_494),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_499),
.B(n_396),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_494),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_456),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_L g571 ( 
.A(n_468),
.B(n_254),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_488),
.A2(n_443),
.B1(n_419),
.B2(n_386),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_522),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_515),
.B(n_397),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_456),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_522),
.Y(n_576)
);

CKINVDCx6p67_ASAP7_75t_R g577 ( 
.A(n_488),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_449),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_461),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_461),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_501),
.A2(n_391),
.B1(n_227),
.B2(n_230),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_449),
.B(n_399),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_461),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_501),
.A2(n_246),
.B1(n_258),
.B2(n_219),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_464),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_456),
.Y(n_586)
);

BUFx4f_ASAP7_75t_L g587 ( 
.A(n_509),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_472),
.B(n_430),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_449),
.B(n_430),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_449),
.A2(n_406),
.B1(n_407),
.B2(n_404),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_455),
.B(n_297),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_464),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_484),
.A2(n_412),
.B1(n_418),
.B2(n_414),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_464),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_464),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_466),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_483),
.B(n_420),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_523),
.Y(n_598)
);

INVxp67_ASAP7_75t_SL g599 ( 
.A(n_487),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_523),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_523),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_466),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_524),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_524),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_487),
.B(n_409),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_484),
.A2(n_441),
.B1(n_431),
.B2(n_423),
.Y(n_606)
);

BUFx8_ASAP7_75t_SL g607 ( 
.A(n_479),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_456),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_484),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_483),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_466),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_524),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_509),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_483),
.B(n_422),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_483),
.B(n_411),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_466),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_455),
.B(n_193),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_455),
.B(n_320),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_484),
.A2(n_217),
.B1(n_237),
.B2(n_223),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_501),
.B(n_317),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_468),
.B(n_254),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_497),
.B(n_421),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_493),
.B(n_321),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_501),
.B(n_317),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_509),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_509),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_493),
.B(n_421),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_493),
.B(n_257),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_476),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_456),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_509),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_479),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_476),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_468),
.B(n_254),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_484),
.A2(n_210),
.B1(n_212),
.B2(n_199),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_497),
.B(n_359),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_509),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_493),
.B(n_317),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_497),
.B(n_362),
.Y(n_639)
);

BUFx4f_ASAP7_75t_L g640 ( 
.A(n_509),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_498),
.B(n_365),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_498),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_456),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_484),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_476),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_456),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_476),
.Y(n_647)
);

AND2x6_ASAP7_75t_L g648 ( 
.A(n_512),
.B(n_297),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_450),
.B(n_261),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_478),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_498),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_484),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_500),
.B(n_502),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_484),
.A2(n_306),
.B1(n_245),
.B2(n_244),
.Y(n_654)
);

NAND3xp33_ASAP7_75t_L g655 ( 
.A(n_512),
.B(n_376),
.C(n_380),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_478),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_518),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_512),
.A2(n_377),
.B1(n_376),
.B2(n_273),
.Y(n_658)
);

BUFx6f_ASAP7_75t_SL g659 ( 
.A(n_519),
.Y(n_659)
);

INVx5_ASAP7_75t_L g660 ( 
.A(n_459),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_500),
.B(n_380),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_500),
.B(n_433),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_512),
.B(n_433),
.C(n_229),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_479),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_519),
.A2(n_258),
.B1(n_355),
.B2(n_354),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_478),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_519),
.A2(n_518),
.B1(n_504),
.B2(n_505),
.Y(n_667)
);

AND3x2_ASAP7_75t_L g668 ( 
.A(n_520),
.B(n_297),
.C(n_194),
.Y(n_668)
);

AND2x6_ASAP7_75t_L g669 ( 
.A(n_519),
.B(n_254),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_502),
.B(n_228),
.Y(n_670)
);

NOR2x1p5_ASAP7_75t_L g671 ( 
.A(n_502),
.B(n_232),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_518),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_518),
.B(n_505),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_450),
.B(n_263),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_519),
.B(n_281),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_518),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_574),
.B(n_520),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_599),
.B(n_504),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_554),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_538),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_L g681 ( 
.A(n_529),
.B(n_520),
.C(n_180),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_534),
.B(n_504),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_543),
.B(n_518),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_538),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_589),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_578),
.A2(n_290),
.B1(n_293),
.B2(n_282),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_543),
.B(n_518),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_534),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_544),
.B(n_504),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_587),
.B(n_254),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_672),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_538),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_568),
.B(n_341),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_544),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_587),
.B(n_254),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_525),
.B(n_341),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_648),
.A2(n_519),
.B1(n_504),
.B2(n_225),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_672),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_542),
.B(n_504),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_SL g700 ( 
.A1(n_531),
.A2(n_214),
.B1(n_264),
.B2(n_262),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_578),
.B(n_519),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_676),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_605),
.B(n_505),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_605),
.B(n_508),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_525),
.B(n_234),
.Y(n_705)
);

BUFx12f_ASAP7_75t_L g706 ( 
.A(n_664),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_587),
.B(n_506),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_554),
.B(n_506),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_525),
.B(n_249),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_673),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_554),
.B(n_506),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_617),
.B(n_506),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_673),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_618),
.B(n_506),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_623),
.B(n_506),
.Y(n_715)
);

AND2x4_ASAP7_75t_SL g716 ( 
.A(n_577),
.B(n_266),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_676),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_640),
.B(n_506),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_538),
.B(n_506),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_661),
.B(n_508),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_565),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_565),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_538),
.B(n_506),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_L g724 ( 
.A(n_541),
.B(n_269),
.C(n_267),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_548),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_640),
.B(n_506),
.Y(n_726)
);

NOR3xp33_ASAP7_75t_L g727 ( 
.A(n_563),
.B(n_272),
.C(n_271),
.Y(n_727)
);

NAND3xp33_ASAP7_75t_L g728 ( 
.A(n_528),
.B(n_655),
.C(n_663),
.Y(n_728)
);

BUFx8_ASAP7_75t_L g729 ( 
.A(n_564),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_598),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_588),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_640),
.B(n_299),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_613),
.A2(n_463),
.B(n_447),
.C(n_514),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_548),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_667),
.B(n_303),
.Y(n_735)
);

AND2x4_ASAP7_75t_SL g736 ( 
.A(n_577),
.B(n_201),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_598),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_600),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_600),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_548),
.B(n_463),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_588),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_548),
.B(n_463),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_548),
.B(n_450),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_567),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_627),
.B(n_451),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_653),
.B(n_451),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_590),
.B(n_275),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_553),
.Y(n_748)
);

NOR2x1p5_ASAP7_75t_L g749 ( 
.A(n_589),
.B(n_283),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_562),
.B(n_451),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_636),
.A2(n_641),
.B1(n_639),
.B2(n_624),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_601),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_601),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_603),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_603),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_604),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_L g757 ( 
.A(n_559),
.B(n_179),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_562),
.B(n_454),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_569),
.B(n_454),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_648),
.A2(n_194),
.B1(n_179),
.B2(n_202),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_569),
.B(n_454),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_604),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_567),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_609),
.B(n_304),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_609),
.B(n_307),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_612),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_582),
.B(n_284),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_612),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_593),
.B(n_286),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_613),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_573),
.B(n_458),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_576),
.B(n_458),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_642),
.B(n_458),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_651),
.B(n_470),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_625),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_648),
.A2(n_591),
.B1(n_559),
.B2(n_625),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_626),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_626),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_628),
.B(n_470),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_644),
.B(n_310),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_644),
.B(n_312),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_671),
.B(n_202),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_631),
.Y(n_783)
);

BUFx12f_ASAP7_75t_L g784 ( 
.A(n_664),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_559),
.B(n_214),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_620),
.A2(n_322),
.B1(n_325),
.B2(n_330),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_606),
.B(n_288),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_631),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_648),
.A2(n_287),
.B1(n_225),
.B2(n_242),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_652),
.B(n_447),
.Y(n_790)
);

AND2x6_ASAP7_75t_SL g791 ( 
.A(n_662),
.B(n_219),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_637),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_526),
.B(n_470),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_526),
.B(n_473),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_530),
.B(n_242),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_637),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_535),
.B(n_537),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_657),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_535),
.B(n_473),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_537),
.B(n_473),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_657),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_540),
.B(n_549),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_540),
.Y(n_803)
);

NOR2xp67_ASAP7_75t_SL g804 ( 
.A(n_652),
.B(n_301),
.Y(n_804)
);

AO221x1_ASAP7_75t_L g805 ( 
.A1(n_619),
.A2(n_654),
.B1(n_635),
.B2(n_549),
.C(n_350),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_658),
.B(n_289),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_622),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_527),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_572),
.A2(n_287),
.B1(n_324),
.B2(n_346),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_559),
.B(n_474),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_527),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_559),
.B(n_260),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_559),
.B(n_474),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_546),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_591),
.B(n_649),
.Y(n_815)
);

O2A1O1Ixp5_ASAP7_75t_L g816 ( 
.A1(n_675),
.A2(n_447),
.B(n_477),
.C(n_474),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_SL g817 ( 
.A(n_553),
.B(n_213),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_591),
.B(n_477),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_546),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_591),
.A2(n_648),
.B1(n_638),
.B2(n_614),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_591),
.B(n_674),
.Y(n_821)
);

NAND2xp33_ASAP7_75t_L g822 ( 
.A(n_591),
.B(n_260),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_552),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_652),
.B(n_597),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_SL g825 ( 
.A(n_550),
.B(n_236),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_560),
.Y(n_826)
);

AO22x2_ASAP7_75t_L g827 ( 
.A1(n_564),
.A2(n_262),
.B1(n_278),
.B2(n_264),
.Y(n_827)
);

AO22x2_ASAP7_75t_L g828 ( 
.A1(n_551),
.A2(n_278),
.B1(n_298),
.B2(n_324),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_560),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_539),
.B(n_298),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_648),
.B(n_477),
.Y(n_831)
);

INVxp67_ASAP7_75t_SL g832 ( 
.A(n_558),
.Y(n_832)
);

INVx8_ASAP7_75t_L g833 ( 
.A(n_659),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_669),
.Y(n_834)
);

OAI22xp33_ASAP7_75t_L g835 ( 
.A1(n_532),
.A2(n_334),
.B1(n_346),
.B2(n_313),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_533),
.B(n_480),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_545),
.B(n_556),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_539),
.B(n_334),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_659),
.A2(n_521),
.B1(n_517),
.B2(n_514),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_547),
.B(n_508),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_670),
.B(n_480),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_539),
.B(n_480),
.Y(n_842)
);

BUFx4_ASAP7_75t_L g843 ( 
.A(n_607),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_659),
.A2(n_557),
.B1(n_581),
.B2(n_584),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_536),
.B(n_246),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_571),
.A2(n_521),
.B(n_517),
.C(n_514),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_710),
.A2(n_665),
.B1(n_329),
.B2(n_347),
.Y(n_847)
);

O2A1O1Ixp5_ASAP7_75t_L g848 ( 
.A1(n_830),
.A2(n_615),
.B(n_561),
.C(n_610),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_740),
.A2(n_610),
.B(n_561),
.Y(n_849)
);

BUFx8_ASAP7_75t_SL g850 ( 
.A(n_843),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_SL g851 ( 
.A(n_748),
.B(n_607),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_728),
.A2(n_837),
.B1(n_751),
.B2(n_795),
.Y(n_852)
);

NAND2x1p5_ASAP7_75t_L g853 ( 
.A(n_680),
.B(n_561),
.Y(n_853)
);

AOI33xp33_ASAP7_75t_L g854 ( 
.A1(n_835),
.A2(n_340),
.A3(n_326),
.B1(n_323),
.B2(n_309),
.B3(n_347),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_680),
.B(n_610),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_680),
.B(n_558),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_742),
.A2(n_621),
.B(n_571),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_807),
.B(n_558),
.Y(n_858)
);

CKINVDCx11_ASAP7_75t_R g859 ( 
.A(n_706),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_677),
.B(n_668),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_713),
.A2(n_241),
.B1(n_302),
.B2(n_632),
.Y(n_861)
);

BUFx8_ASAP7_75t_L g862 ( 
.A(n_706),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_690),
.A2(n_580),
.B(n_579),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_720),
.B(n_688),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_720),
.B(n_566),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_790),
.A2(n_634),
.B(n_621),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_790),
.A2(n_634),
.B(n_570),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_694),
.B(n_566),
.Y(n_868)
);

OAI21xp33_ASAP7_75t_L g869 ( 
.A1(n_806),
.A2(n_294),
.B(n_292),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_809),
.A2(n_513),
.B(n_521),
.C(n_517),
.Y(n_870)
);

AO21x1_ASAP7_75t_L g871 ( 
.A1(n_690),
.A2(n_279),
.B(n_276),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_703),
.B(n_566),
.Y(n_872)
);

OAI21xp33_ASAP7_75t_L g873 ( 
.A1(n_747),
.A2(n_300),
.B(n_296),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_721),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_703),
.B(n_704),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_704),
.B(n_570),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_735),
.A2(n_510),
.B(n_513),
.C(n_656),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_701),
.B(n_570),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_769),
.A2(n_329),
.B(n_326),
.C(n_323),
.Y(n_879)
);

NAND2x1p5_ASAP7_75t_L g880 ( 
.A(n_680),
.B(n_575),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_701),
.B(n_575),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_680),
.A2(n_586),
.B(n_575),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_795),
.B(n_586),
.Y(n_883)
);

O2A1O1Ixp5_ASAP7_75t_L g884 ( 
.A1(n_830),
.A2(n_586),
.B(n_608),
.C(n_630),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_705),
.B(n_632),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_721),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_722),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_795),
.B(n_841),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_685),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_725),
.A2(n_630),
.B(n_608),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_691),
.B(n_608),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_748),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_725),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_683),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_725),
.A2(n_734),
.B(n_723),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_722),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_784),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_691),
.B(n_630),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_695),
.A2(n_580),
.B(n_579),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_731),
.B(n_305),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_698),
.B(n_643),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_725),
.A2(n_646),
.B(n_643),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_725),
.A2(n_646),
.B(n_643),
.Y(n_903)
);

CKINVDCx16_ASAP7_75t_R g904 ( 
.A(n_817),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_744),
.B(n_510),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_734),
.B(n_646),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_784),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_739),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_698),
.B(n_702),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_734),
.A2(n_555),
.B(n_452),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_695),
.A2(n_743),
.B(n_797),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_702),
.B(n_717),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_787),
.A2(n_309),
.B(n_285),
.C(n_280),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_L g914 ( 
.A(n_693),
.B(n_311),
.C(n_308),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_739),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_734),
.A2(n_555),
.B(n_452),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_717),
.B(n_583),
.Y(n_917)
);

BUFx12f_ASAP7_75t_L g918 ( 
.A(n_729),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_734),
.A2(n_555),
.B(n_452),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_836),
.B(n_583),
.Y(n_920)
);

OR2x6_ASAP7_75t_L g921 ( 
.A(n_833),
.B(n_285),
.Y(n_921)
);

INVx5_ASAP7_75t_L g922 ( 
.A(n_834),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_770),
.B(n_585),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_770),
.A2(n_340),
.B(n_350),
.C(n_353),
.Y(n_924)
);

AO21x1_ASAP7_75t_L g925 ( 
.A1(n_732),
.A2(n_353),
.B(n_356),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_764),
.A2(n_669),
.B1(n_666),
.B2(n_611),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_729),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_755),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_719),
.A2(n_555),
.B(n_452),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_833),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_792),
.B(n_585),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_709),
.B(n_510),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_792),
.B(n_592),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_755),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_776),
.A2(n_629),
.B1(n_666),
.B2(n_594),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_802),
.A2(n_555),
.B(n_660),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_741),
.B(n_314),
.Y(n_937)
);

AND2x4_ASAP7_75t_SL g938 ( 
.A(n_834),
.B(n_354),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_798),
.B(n_592),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_756),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_798),
.B(n_594),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_730),
.B(n_595),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_737),
.B(n_595),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_744),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_738),
.B(n_596),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_840),
.B(n_315),
.Y(n_946)
);

AND2x2_ASAP7_75t_SL g947 ( 
.A(n_757),
.B(n_355),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_756),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_684),
.B(n_596),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_815),
.A2(n_660),
.B(n_629),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_782),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_735),
.A2(n_513),
.B(n_656),
.C(n_650),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_821),
.A2(n_660),
.B(n_611),
.Y(n_953)
);

OAI21xp33_ASAP7_75t_L g954 ( 
.A1(n_767),
.A2(n_845),
.B(n_840),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_752),
.B(n_602),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_824),
.A2(n_660),
.B(n_616),
.Y(n_956)
);

NOR2xp67_ASAP7_75t_L g957 ( 
.A(n_786),
.B(n_686),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_824),
.A2(n_660),
.B(n_616),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_683),
.A2(n_650),
.B(n_647),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_753),
.B(n_602),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_844),
.A2(n_647),
.B1(n_645),
.B2(n_633),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_754),
.B(n_633),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_712),
.A2(n_645),
.B(n_503),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_833),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_762),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_687),
.A2(n_669),
.B1(n_495),
.B2(n_507),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_833),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_687),
.A2(n_669),
.B(n_460),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_714),
.A2(n_511),
.B(n_507),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_L g970 ( 
.A1(n_838),
.A2(n_511),
.B(n_507),
.C(n_503),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_820),
.A2(n_495),
.B1(n_319),
.B2(n_327),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_763),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_779),
.B(n_503),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_766),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_845),
.A2(n_511),
.B(n_507),
.C(n_503),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_764),
.A2(n_669),
.B1(n_511),
.B2(n_489),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_696),
.B(n_316),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_684),
.B(n_495),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_766),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_678),
.B(n_669),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_803),
.B(n_481),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_825),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_715),
.A2(n_478),
.B(n_496),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_763),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_707),
.A2(n_496),
.B(n_482),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_716),
.B(n_328),
.Y(n_986)
);

NAND2xp33_ASAP7_75t_L g987 ( 
.A(n_834),
.B(n_331),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_765),
.A2(n_489),
.B1(n_481),
.B2(n_491),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_765),
.A2(n_486),
.B(n_481),
.C(n_491),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_775),
.B(n_485),
.Y(n_990)
);

NOR2x1_ASAP7_75t_L g991 ( 
.A(n_749),
.B(n_460),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_780),
.A2(n_489),
.B(n_485),
.C(n_491),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_780),
.A2(n_490),
.B(n_486),
.C(n_485),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_684),
.B(n_495),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_777),
.B(n_486),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_707),
.A2(n_496),
.B(n_482),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_718),
.A2(n_496),
.B(n_482),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_SL g998 ( 
.A(n_729),
.B(n_333),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_716),
.B(n_335),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_778),
.B(n_490),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_783),
.B(n_490),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_781),
.A2(n_460),
.B(n_495),
.C(n_482),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_768),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_718),
.A2(n_726),
.B(n_842),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_768),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_692),
.B(n_495),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_726),
.A2(n_460),
.B(n_475),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_788),
.B(n_460),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_679),
.Y(n_1009)
);

OAI21xp33_ASAP7_75t_L g1010 ( 
.A1(n_681),
.A2(n_351),
.B(n_338),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_828),
.A2(n_352),
.B(n_339),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_692),
.B(n_492),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_796),
.A2(n_337),
.B(n_342),
.C(n_344),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_733),
.A2(n_460),
.B(n_345),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_808),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_801),
.B(n_459),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_736),
.B(n_3),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_781),
.A2(n_492),
.B1(n_475),
.B2(n_467),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_679),
.A2(n_805),
.B1(n_732),
.B2(n_838),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_692),
.B(n_459),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_810),
.B(n_492),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_813),
.B(n_492),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_808),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_708),
.A2(n_475),
.B(n_467),
.Y(n_1024)
);

INVx5_ASAP7_75t_L g1025 ( 
.A(n_834),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_736),
.B(n_3),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_782),
.B(n_5),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_682),
.B(n_5),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_689),
.A2(n_475),
.B(n_467),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_746),
.B(n_459),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_819),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_711),
.A2(n_475),
.B(n_467),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_745),
.B(n_459),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_819),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_846),
.A2(n_492),
.B(n_475),
.C(n_467),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_699),
.B(n_459),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_826),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_832),
.B(n_459),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_782),
.A2(n_492),
.B1(n_475),
.B2(n_467),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_964),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_849),
.A2(n_812),
.B(n_785),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_965),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_875),
.B(n_888),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_951),
.B(n_724),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_954),
.B(n_861),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1004),
.A2(n_793),
.B(n_794),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_852),
.A2(n_816),
.B(n_727),
.C(n_839),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_853),
.A2(n_857),
.B(n_911),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_984),
.B(n_944),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_977),
.B(n_889),
.Y(n_1050)
);

AND2x6_ASAP7_75t_L g1051 ( 
.A(n_964),
.B(n_834),
.Y(n_1051)
);

CKINVDCx8_ASAP7_75t_R g1052 ( 
.A(n_904),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_974),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_879),
.A2(n_700),
.B(n_773),
.C(n_772),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_864),
.B(n_932),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_865),
.B(n_799),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_965),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_974),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_964),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_892),
.Y(n_1060)
);

AOI22x1_ASAP7_75t_L g1061 ( 
.A1(n_866),
.A2(n_828),
.B1(n_827),
.B2(n_811),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_889),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_893),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_879),
.A2(n_774),
.B(n_771),
.C(n_812),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_944),
.Y(n_1065)
);

AOI21xp33_ASAP7_75t_L g1066 ( 
.A1(n_946),
.A2(n_828),
.B(n_827),
.Y(n_1066)
);

OAI21xp33_ASAP7_75t_L g1067 ( 
.A1(n_946),
.A2(n_828),
.B(n_827),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_984),
.B(n_818),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1028),
.B(n_827),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1003),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1003),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1028),
.B(n_750),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_964),
.Y(n_1073)
);

INVxp67_ASAP7_75t_L g1074 ( 
.A(n_1017),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_957),
.B(n_697),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1005),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_972),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_977),
.B(n_791),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_913),
.A2(n_757),
.B(n_785),
.C(n_822),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_853),
.A2(n_822),
.B(n_800),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_982),
.B(n_831),
.Y(n_1081)
);

O2A1O1Ixp5_ASAP7_75t_L g1082 ( 
.A1(n_925),
.A2(n_804),
.B(n_759),
.C(n_761),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_895),
.A2(n_758),
.B(n_789),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1005),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_930),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_905),
.B(n_760),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_905),
.B(n_914),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_893),
.A2(n_826),
.B(n_829),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_855),
.A2(n_829),
.B(n_823),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_874),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_872),
.B(n_814),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_SL g1092 ( 
.A1(n_975),
.A2(n_173),
.B(n_172),
.C(n_171),
.Y(n_1092)
);

AOI33xp33_ASAP7_75t_L g1093 ( 
.A1(n_885),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.B3(n_11),
.Y(n_1093)
);

AO21x2_ASAP7_75t_L g1094 ( 
.A1(n_1019),
.A2(n_136),
.B(n_80),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_855),
.A2(n_475),
.B(n_467),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_876),
.B(n_492),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1021),
.A2(n_475),
.B(n_467),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_909),
.A2(n_475),
.B(n_467),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_940),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_973),
.B(n_492),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_947),
.A2(n_492),
.B1(n_467),
.B2(n_462),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_860),
.B(n_7),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1015),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_860),
.B(n_14),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1013),
.A2(n_15),
.B(n_18),
.C(n_20),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_920),
.B(n_492),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_972),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1015),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_979),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_912),
.A2(n_883),
.B(n_881),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_886),
.B(n_462),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_SL g1112 ( 
.A(n_907),
.B(n_462),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_878),
.A2(n_462),
.B(n_459),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_SL g1114 ( 
.A(n_862),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1009),
.B(n_462),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_894),
.A2(n_462),
.B1(n_459),
.B2(n_27),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_967),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_947),
.A2(n_462),
.B1(n_459),
.B2(n_27),
.Y(n_1118)
);

NOR3xp33_ASAP7_75t_SL g1119 ( 
.A(n_873),
.B(n_23),
.C(n_24),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_869),
.B(n_900),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1011),
.A2(n_462),
.B(n_31),
.C(n_34),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_SL g1122 ( 
.A1(n_1014),
.A2(n_161),
.B(n_160),
.C(n_159),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1013),
.A2(n_462),
.B(n_34),
.C(n_35),
.Y(n_1123)
);

AOI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_971),
.A2(n_28),
.B(n_36),
.Y(n_1124)
);

NAND2xp33_ASAP7_75t_SL g1125 ( 
.A(n_967),
.B(n_39),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_887),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_867),
.A2(n_147),
.B(n_145),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_959),
.A2(n_142),
.B(n_140),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1023),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_894),
.A2(n_40),
.B1(n_41),
.B2(n_45),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1026),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_922),
.B(n_1025),
.Y(n_1132)
);

AOI22x1_ASAP7_75t_L g1133 ( 
.A1(n_896),
.A2(n_138),
.B1(n_134),
.B2(n_133),
.Y(n_1133)
);

BUFx12f_ASAP7_75t_L g1134 ( 
.A(n_859),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_922),
.B(n_131),
.Y(n_1135)
);

AO21x1_ASAP7_75t_L g1136 ( 
.A1(n_877),
.A2(n_45),
.B(n_47),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_966),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_908),
.B(n_128),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_915),
.B(n_51),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_928),
.B(n_120),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_897),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1027),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_922),
.Y(n_1143)
);

OR2x6_ASAP7_75t_SL g1144 ( 
.A(n_850),
.B(n_55),
.Y(n_1144)
);

AND2x6_ASAP7_75t_L g1145 ( 
.A(n_991),
.B(n_116),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_921),
.B(n_922),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1023),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_966),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_862),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_918),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_934),
.B(n_103),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_856),
.A2(n_98),
.B(n_95),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_948),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_900),
.A2(n_937),
.B(n_999),
.C(n_952),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_924),
.A2(n_60),
.B(n_61),
.C(n_66),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_1025),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1025),
.Y(n_1157)
);

OR2x6_ASAP7_75t_L g1158 ( 
.A(n_927),
.B(n_74),
.Y(n_1158)
);

INVx6_ASAP7_75t_L g1159 ( 
.A(n_1025),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_856),
.A2(n_82),
.B(n_69),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_924),
.A2(n_68),
.B(n_70),
.C(n_71),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_937),
.B(n_70),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_986),
.B(n_72),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_999),
.B(n_1010),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_998),
.B(n_847),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_975),
.A2(n_870),
.B(n_858),
.C(n_1035),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_938),
.B(n_1034),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_851),
.B(n_921),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_921),
.B(n_868),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_906),
.A2(n_848),
.B(n_980),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_906),
.A2(n_1033),
.B(n_882),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_938),
.B(n_847),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_978),
.B(n_994),
.Y(n_1173)
);

BUFx8_ASAP7_75t_L g1174 ( 
.A(n_1031),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_854),
.B(n_981),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1037),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1030),
.B(n_990),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_978),
.B(n_994),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_923),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_995),
.B(n_1000),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1001),
.B(n_942),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_854),
.B(n_1039),
.Y(n_1182)
);

BUFx12f_ASAP7_75t_L g1183 ( 
.A(n_880),
.Y(n_1183)
);

NOR2xp67_ASAP7_75t_SL g1184 ( 
.A(n_968),
.B(n_903),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_880),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_890),
.A2(n_902),
.B(n_891),
.Y(n_1186)
);

AO21x1_ASAP7_75t_L g1187 ( 
.A1(n_989),
.A2(n_992),
.B(n_993),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_961),
.Y(n_1188)
);

NOR2x1_ASAP7_75t_L g1189 ( 
.A(n_987),
.B(n_1006),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_943),
.B(n_962),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_945),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_898),
.A2(n_901),
.B(n_1038),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1006),
.B(n_949),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1035),
.A2(n_960),
.B(n_955),
.C(n_871),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_SL g1195 ( 
.A(n_1002),
.B(n_935),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_R g1196 ( 
.A(n_1008),
.B(n_1016),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_931),
.A2(n_939),
.B1(n_933),
.B2(n_941),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_988),
.B(n_976),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_926),
.B(n_917),
.Y(n_1199)
);

CKINVDCx6p67_ASAP7_75t_R g1200 ( 
.A(n_1134),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1050),
.B(n_949),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1176),
.Y(n_1202)
);

INVxp67_ASAP7_75t_SL g1203 ( 
.A(n_1077),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1062),
.B(n_1022),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1078),
.B(n_1120),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1186),
.A2(n_1171),
.B(n_1048),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1046),
.A2(n_963),
.B(n_1022),
.Y(n_1207)
);

OAI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1055),
.A2(n_1018),
.B1(n_1036),
.B2(n_1020),
.Y(n_1208)
);

AOI221x1_ASAP7_75t_L g1209 ( 
.A1(n_1066),
.A2(n_1067),
.B1(n_1124),
.B2(n_1154),
.C(n_1121),
.Y(n_1209)
);

OA21x2_ASAP7_75t_L g1210 ( 
.A1(n_1170),
.A2(n_863),
.B(n_899),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1065),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_1174),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1090),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1099),
.Y(n_1214)
);

AO21x1_ASAP7_75t_L g1215 ( 
.A1(n_1066),
.A2(n_969),
.B(n_953),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1046),
.A2(n_1021),
.B(n_950),
.Y(n_1216)
);

BUFx8_ASAP7_75t_L g1217 ( 
.A(n_1149),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1045),
.A2(n_1012),
.B1(n_996),
.B2(n_997),
.Y(n_1218)
);

NOR2xp67_ASAP7_75t_L g1219 ( 
.A(n_1074),
.B(n_1007),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1164),
.A2(n_1012),
.B1(n_985),
.B2(n_958),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_1107),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1102),
.A2(n_956),
.B(n_1029),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1097),
.A2(n_929),
.B(n_983),
.Y(n_1223)
);

AOI221x1_ASAP7_75t_L g1224 ( 
.A1(n_1124),
.A2(n_1032),
.B1(n_1024),
.B2(n_936),
.C(n_919),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1109),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1041),
.A2(n_884),
.B(n_910),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1089),
.A2(n_970),
.B(n_916),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1192),
.A2(n_1110),
.B(n_1113),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1053),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1177),
.A2(n_1080),
.B(n_1180),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1058),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1180),
.A2(n_1056),
.B(n_1181),
.Y(n_1232)
);

AOI221xp5_ASAP7_75t_L g1233 ( 
.A1(n_1104),
.A2(n_1130),
.B1(n_1148),
.B2(n_1137),
.C(n_1162),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_SL g1234 ( 
.A1(n_1122),
.A2(n_1047),
.B(n_1075),
.C(n_1123),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1174),
.Y(n_1235)
);

AOI31xp67_ASAP7_75t_L g1236 ( 
.A1(n_1199),
.A2(n_1198),
.A3(n_1069),
.B(n_1072),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1095),
.A2(n_1098),
.B(n_1088),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1166),
.A2(n_1083),
.B(n_1194),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1096),
.A2(n_1111),
.B(n_1100),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1056),
.A2(n_1181),
.B(n_1190),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1190),
.A2(n_1043),
.B(n_1197),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1043),
.A2(n_1197),
.B(n_1195),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1055),
.A2(n_1143),
.B(n_1106),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1049),
.B(n_1146),
.Y(n_1244)
);

OAI21xp33_ASAP7_75t_L g1245 ( 
.A1(n_1119),
.A2(n_1118),
.B(n_1165),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1187),
.A2(n_1136),
.A3(n_1128),
.B(n_1193),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1064),
.A2(n_1188),
.B(n_1082),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1131),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1191),
.B(n_1179),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1111),
.A2(n_1100),
.B(n_1138),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_1060),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1087),
.A2(n_1044),
.B1(n_1169),
.B2(n_1168),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1138),
.A2(n_1140),
.B(n_1151),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1142),
.B(n_1163),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_SL g1255 ( 
.A1(n_1130),
.A2(n_1148),
.B(n_1137),
.Y(n_1255)
);

AOI221x1_ASAP7_75t_L g1256 ( 
.A1(n_1127),
.A2(n_1125),
.B1(n_1160),
.B2(n_1116),
.C(n_1182),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1061),
.A2(n_1091),
.B(n_1140),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1079),
.A2(n_1091),
.B(n_1086),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1071),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1052),
.B(n_1141),
.Y(n_1260)
);

AO21x1_ASAP7_75t_L g1261 ( 
.A1(n_1105),
.A2(n_1175),
.B(n_1054),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1059),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1151),
.A2(n_1115),
.B(n_1139),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1143),
.A2(n_1132),
.B(n_1189),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1167),
.A2(n_1081),
.B(n_1068),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1076),
.B(n_1070),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1044),
.B(n_1049),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1172),
.A2(n_1116),
.B1(n_1159),
.B2(n_1146),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1114),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1084),
.Y(n_1270)
);

BUFx10_ASAP7_75t_L g1271 ( 
.A(n_1158),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1112),
.B(n_1068),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1103),
.A2(n_1108),
.B(n_1147),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1129),
.A2(n_1152),
.B(n_1133),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1042),
.B(n_1057),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1126),
.B(n_1153),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1092),
.A2(n_1094),
.B(n_1173),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1178),
.A2(n_1184),
.A3(n_1094),
.B(n_1040),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1155),
.A2(n_1161),
.B(n_1093),
.C(n_1135),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1159),
.A2(n_1158),
.B1(n_1063),
.B2(n_1156),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1185),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1196),
.B(n_1063),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1156),
.A2(n_1157),
.B(n_1185),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1159),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1156),
.A2(n_1157),
.B(n_1101),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1157),
.A2(n_1185),
.B(n_1117),
.Y(n_1286)
);

OAI22x1_ASAP7_75t_L g1287 ( 
.A1(n_1040),
.A2(n_1144),
.B1(n_1158),
.B2(n_1145),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1085),
.A2(n_1117),
.B(n_1059),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1085),
.A2(n_1117),
.B(n_1059),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1051),
.A2(n_1145),
.B(n_1183),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1073),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1051),
.B(n_1145),
.Y(n_1292)
);

AOI211x1_ASAP7_75t_L g1293 ( 
.A1(n_1145),
.A2(n_1051),
.B(n_1073),
.C(n_1085),
.Y(n_1293)
);

OAI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1150),
.A2(n_1073),
.B1(n_1145),
.B2(n_1051),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1051),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1176),
.Y(n_1296)
);

BUFx10_ASAP7_75t_L g1297 ( 
.A(n_1060),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1186),
.A2(n_1171),
.B(n_1048),
.Y(n_1298)
);

CKINVDCx11_ASAP7_75t_R g1299 ( 
.A(n_1134),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1050),
.B(n_885),
.Y(n_1300)
);

BUFx12f_ASAP7_75t_L g1301 ( 
.A(n_1134),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1154),
.A2(n_677),
.B(n_1078),
.C(n_529),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1048),
.A2(n_1046),
.B(n_725),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1043),
.B(n_1055),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1170),
.A2(n_1048),
.B(n_1046),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1043),
.B(n_1055),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1176),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1187),
.A2(n_1170),
.A3(n_1035),
.B(n_1048),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1048),
.A2(n_725),
.B(n_680),
.Y(n_1309)
);

O2A1O1Ixp33_ASAP7_75t_SL g1310 ( 
.A1(n_1154),
.A2(n_1121),
.B(n_1066),
.C(n_1122),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1187),
.A2(n_1170),
.A3(n_1035),
.B(n_1048),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1048),
.A2(n_1046),
.B(n_725),
.Y(n_1312)
);

AO32x2_ASAP7_75t_L g1313 ( 
.A1(n_1130),
.A2(n_1148),
.A3(n_1137),
.B1(n_1116),
.B2(n_1197),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1055),
.A2(n_875),
.B1(n_852),
.B2(n_1118),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1050),
.B(n_885),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1070),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1176),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_SL g1318 ( 
.A(n_1078),
.B(n_751),
.C(n_677),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1048),
.A2(n_1046),
.B(n_725),
.Y(n_1319)
);

NOR2x1_ASAP7_75t_SL g1320 ( 
.A(n_1156),
.B(n_1157),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1154),
.A2(n_677),
.B(n_1078),
.C(n_529),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1048),
.A2(n_725),
.B(n_680),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1176),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1176),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1043),
.B(n_1055),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1050),
.B(n_904),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1050),
.B(n_885),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1176),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1176),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1159),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1176),
.Y(n_1331)
);

AO32x2_ASAP7_75t_L g1332 ( 
.A1(n_1130),
.A2(n_1148),
.A3(n_1137),
.B1(n_1116),
.B2(n_1197),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1187),
.A2(n_1170),
.A3(n_1035),
.B(n_1048),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1159),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1048),
.A2(n_725),
.B(n_680),
.Y(n_1335)
);

AO31x2_ASAP7_75t_L g1336 ( 
.A1(n_1187),
.A2(n_1170),
.A3(n_1035),
.B(n_1048),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1062),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1120),
.A2(n_1045),
.B(n_1154),
.C(n_1164),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_SL g1339 ( 
.A1(n_1154),
.A2(n_1121),
.B(n_1066),
.C(n_1122),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1176),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1048),
.A2(n_725),
.B(n_680),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1048),
.A2(n_725),
.B(n_680),
.Y(n_1342)
);

NOR2xp67_ASAP7_75t_L g1343 ( 
.A(n_1074),
.B(n_706),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1055),
.A2(n_875),
.B1(n_852),
.B2(n_1118),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1048),
.A2(n_725),
.B(n_680),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1186),
.A2(n_1171),
.B(n_1048),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1176),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1048),
.A2(n_1046),
.B(n_725),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1176),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1174),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1048),
.A2(n_1046),
.B(n_725),
.Y(n_1351)
);

AOI31xp67_ASAP7_75t_L g1352 ( 
.A1(n_1199),
.A2(n_1019),
.A3(n_852),
.B(n_824),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1055),
.A2(n_875),
.B1(n_852),
.B2(n_1118),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1048),
.A2(n_1046),
.B(n_725),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1060),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1062),
.Y(n_1356)
);

AO21x1_ASAP7_75t_L g1357 ( 
.A1(n_1120),
.A2(n_1066),
.B(n_1072),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1176),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1048),
.A2(n_1046),
.B(n_725),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1318),
.A2(n_1233),
.B1(n_1205),
.B2(n_1245),
.Y(n_1360)
);

OAI21xp33_ASAP7_75t_L g1361 ( 
.A1(n_1338),
.A2(n_1321),
.B(n_1302),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1300),
.A2(n_1327),
.B1(n_1315),
.B2(n_1353),
.Y(n_1362)
);

CKINVDCx6p67_ASAP7_75t_R g1363 ( 
.A(n_1301),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1255),
.A2(n_1233),
.B1(n_1252),
.B2(n_1306),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1261),
.A2(n_1353),
.B1(n_1314),
.B2(n_1344),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1299),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1314),
.A2(n_1344),
.B1(n_1242),
.B2(n_1357),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1337),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_1240),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1304),
.A2(n_1306),
.B1(n_1325),
.B2(n_1238),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1304),
.A2(n_1325),
.B1(n_1326),
.B2(n_1282),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1271),
.A2(n_1267),
.B1(n_1280),
.B2(n_1201),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1282),
.A2(n_1232),
.B1(n_1249),
.B2(n_1221),
.Y(n_1373)
);

BUFx8_ASAP7_75t_SL g1374 ( 
.A(n_1251),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1238),
.A2(n_1258),
.B1(n_1247),
.B2(n_1287),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1262),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1276),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1254),
.B(n_1244),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1202),
.Y(n_1379)
);

CKINVDCx11_ASAP7_75t_R g1380 ( 
.A(n_1355),
.Y(n_1380)
);

BUFx4f_ASAP7_75t_SL g1381 ( 
.A(n_1200),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1356),
.Y(n_1382)
);

INVx8_ASAP7_75t_L g1383 ( 
.A(n_1262),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1262),
.Y(n_1384)
);

BUFx8_ASAP7_75t_L g1385 ( 
.A(n_1235),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1211),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1213),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1297),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1284),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1214),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1249),
.A2(n_1343),
.B1(n_1272),
.B2(n_1203),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1217),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1297),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_1217),
.Y(n_1394)
);

CKINVDCx11_ASAP7_75t_R g1395 ( 
.A(n_1271),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1244),
.B(n_1248),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1316),
.Y(n_1397)
);

BUFx12f_ASAP7_75t_L g1398 ( 
.A(n_1212),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1269),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1241),
.B(n_1204),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1260),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1284),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1280),
.A2(n_1279),
.B1(n_1268),
.B2(n_1347),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1258),
.A2(n_1247),
.B1(n_1268),
.B2(n_1296),
.Y(n_1404)
);

INVx6_ASAP7_75t_L g1405 ( 
.A(n_1320),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1330),
.Y(n_1406)
);

INVx2_ASAP7_75t_R g1407 ( 
.A(n_1295),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1225),
.B(n_1307),
.Y(n_1408)
);

OAI21xp33_ASAP7_75t_L g1409 ( 
.A1(n_1222),
.A2(n_1331),
.B(n_1329),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1350),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1317),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1323),
.A2(n_1324),
.B1(n_1358),
.B2(n_1340),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1313),
.A2(n_1332),
.B1(n_1277),
.B2(n_1292),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1330),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1328),
.B(n_1349),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1270),
.Y(n_1416)
);

BUFx12f_ASAP7_75t_L g1417 ( 
.A(n_1334),
.Y(n_1417)
);

INVx6_ASAP7_75t_L g1418 ( 
.A(n_1334),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1219),
.A2(n_1229),
.B1(n_1231),
.B2(n_1259),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1290),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1277),
.A2(n_1230),
.B1(n_1332),
.B2(n_1313),
.Y(n_1421)
);

OAI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1209),
.A2(n_1256),
.B1(n_1332),
.B2(n_1313),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1275),
.A2(n_1215),
.B1(n_1265),
.B2(n_1305),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1266),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1281),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1266),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1291),
.Y(n_1427)
);

CKINVDCx11_ASAP7_75t_R g1428 ( 
.A(n_1294),
.Y(n_1428)
);

BUFx8_ASAP7_75t_L g1429 ( 
.A(n_1288),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1292),
.A2(n_1243),
.B1(n_1264),
.B2(n_1285),
.Y(n_1430)
);

BUFx12f_ASAP7_75t_L g1431 ( 
.A(n_1288),
.Y(n_1431)
);

OAI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1303),
.A2(n_1354),
.B1(n_1351),
.B2(n_1348),
.Y(n_1432)
);

BUFx12f_ASAP7_75t_L g1433 ( 
.A(n_1289),
.Y(n_1433)
);

BUFx4f_ASAP7_75t_L g1434 ( 
.A(n_1263),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1234),
.A2(n_1339),
.B1(n_1310),
.B2(n_1208),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1236),
.Y(n_1436)
);

BUFx12f_ASAP7_75t_L g1437 ( 
.A(n_1289),
.Y(n_1437)
);

BUFx8_ASAP7_75t_L g1438 ( 
.A(n_1286),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1263),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1305),
.A2(n_1285),
.B1(n_1253),
.B2(n_1257),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1293),
.A2(n_1359),
.B1(n_1319),
.B2(n_1312),
.Y(n_1441)
);

CKINVDCx11_ASAP7_75t_R g1442 ( 
.A(n_1283),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1257),
.A2(n_1303),
.B1(n_1354),
.B2(n_1351),
.Y(n_1443)
);

CKINVDCx6p67_ASAP7_75t_R g1444 ( 
.A(n_1278),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1274),
.B(n_1359),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1207),
.A2(n_1216),
.B1(n_1312),
.B2(n_1348),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1319),
.A2(n_1220),
.B1(n_1218),
.B2(n_1345),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1207),
.A2(n_1216),
.B1(n_1239),
.B2(n_1210),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1226),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1210),
.A2(n_1250),
.B1(n_1226),
.B2(n_1228),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1309),
.A2(n_1322),
.B1(n_1335),
.B2(n_1342),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1308),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1308),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1341),
.A2(n_1206),
.B1(n_1346),
.B2(n_1298),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1352),
.A2(n_1246),
.B1(n_1237),
.B2(n_1227),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1246),
.A2(n_1223),
.B1(n_1311),
.B2(n_1333),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1246),
.Y(n_1457)
);

BUFx8_ASAP7_75t_SL g1458 ( 
.A(n_1224),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1336),
.B(n_1311),
.Y(n_1459)
);

BUFx10_ASAP7_75t_L g1460 ( 
.A(n_1333),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1333),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1336),
.A2(n_1338),
.B(n_1321),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1336),
.A2(n_751),
.B1(n_1338),
.B2(n_677),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1276),
.Y(n_1464)
);

INVx6_ASAP7_75t_L g1465 ( 
.A(n_1297),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_SL g1466 ( 
.A(n_1297),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1318),
.A2(n_1233),
.B1(n_1045),
.B2(n_1205),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1300),
.A2(n_1078),
.B1(n_817),
.B2(n_516),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1297),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1300),
.A2(n_1078),
.B1(n_817),
.B2(n_516),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1262),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1318),
.A2(n_1078),
.B1(n_885),
.B2(n_453),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1300),
.A2(n_1078),
.B1(n_817),
.B2(n_516),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1297),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1276),
.Y(n_1475)
);

CKINVDCx8_ASAP7_75t_R g1476 ( 
.A(n_1235),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_1251),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1273),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1318),
.A2(n_1233),
.B1(n_1045),
.B2(n_1205),
.Y(n_1479)
);

INVx8_ASAP7_75t_L g1480 ( 
.A(n_1262),
.Y(n_1480)
);

BUFx12f_ASAP7_75t_L g1481 ( 
.A(n_1299),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1276),
.Y(n_1482)
);

BUFx8_ASAP7_75t_SL g1483 ( 
.A(n_1301),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1276),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1338),
.A2(n_751),
.B1(n_677),
.B2(n_1233),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1273),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1300),
.B(n_1315),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1337),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1300),
.B(n_1315),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1300),
.A2(n_1078),
.B1(n_817),
.B2(n_516),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1337),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1276),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1276),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1337),
.Y(n_1494)
);

BUFx12f_ASAP7_75t_L g1495 ( 
.A(n_1299),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1300),
.A2(n_1078),
.B1(n_817),
.B2(n_516),
.Y(n_1496)
);

CKINVDCx16_ASAP7_75t_R g1497 ( 
.A(n_1251),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1273),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1338),
.A2(n_751),
.B1(n_677),
.B2(n_1233),
.Y(n_1499)
);

BUFx4f_ASAP7_75t_L g1500 ( 
.A(n_1301),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1300),
.A2(n_1078),
.B1(n_817),
.B2(n_516),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1452),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1368),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1452),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1413),
.B(n_1462),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1453),
.Y(n_1506)
);

BUFx12f_ASAP7_75t_SL g1507 ( 
.A(n_1420),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1459),
.B(n_1367),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1386),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1453),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1449),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1485),
.A2(n_1499),
.B1(n_1479),
.B2(n_1467),
.Y(n_1512)
);

BUFx10_ASAP7_75t_L g1513 ( 
.A(n_1466),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1369),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1369),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1367),
.B(n_1365),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1439),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1370),
.B(n_1364),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1445),
.A2(n_1454),
.B(n_1451),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1436),
.A2(n_1421),
.B(n_1450),
.Y(n_1520)
);

NAND4xp25_ASAP7_75t_SL g1521 ( 
.A(n_1468),
.B(n_1501),
.C(n_1496),
.D(n_1490),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1451),
.A2(n_1450),
.B(n_1447),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1488),
.Y(n_1523)
);

OAI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1467),
.A2(n_1479),
.B1(n_1470),
.B2(n_1473),
.C(n_1472),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1370),
.B(n_1364),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1446),
.A2(n_1448),
.B(n_1441),
.Y(n_1526)
);

NOR2x1_ASAP7_75t_R g1527 ( 
.A(n_1366),
.B(n_1481),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1494),
.Y(n_1528)
);

NOR2x1_ASAP7_75t_SL g1529 ( 
.A(n_1403),
.B(n_1431),
.Y(n_1529)
);

CKINVDCx11_ASAP7_75t_R g1530 ( 
.A(n_1495),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1400),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1438),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1457),
.Y(n_1533)
);

OAI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1463),
.A2(n_1361),
.B(n_1365),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1461),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1458),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1487),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1439),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1478),
.A2(n_1498),
.B(n_1486),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1434),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1421),
.A2(n_1456),
.B(n_1375),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1423),
.A2(n_1404),
.B(n_1435),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1360),
.A2(n_1362),
.B1(n_1428),
.B2(n_1372),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1461),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1432),
.A2(n_1375),
.B(n_1422),
.Y(n_1545)
);

AO21x2_ASAP7_75t_L g1546 ( 
.A1(n_1432),
.A2(n_1422),
.B(n_1409),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1434),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1371),
.B(n_1373),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1444),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1460),
.Y(n_1550)
);

AOI222xp33_ASAP7_75t_L g1551 ( 
.A1(n_1360),
.A2(n_1428),
.B1(n_1489),
.B2(n_1404),
.C1(n_1377),
.C2(n_1484),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1460),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1426),
.B(n_1379),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1426),
.Y(n_1554)
);

INVx3_ASAP7_75t_SL g1555 ( 
.A(n_1405),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1387),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1390),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1411),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1438),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1416),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1424),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1464),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1382),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1475),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1423),
.A2(n_1419),
.B(n_1412),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1482),
.B(n_1492),
.Y(n_1566)
);

INVxp33_ASAP7_75t_SL g1567 ( 
.A(n_1380),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1493),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1419),
.B(n_1412),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1429),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1397),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1429),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1391),
.A2(n_1430),
.B(n_1455),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1491),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1374),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1433),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1443),
.A2(n_1440),
.B(n_1408),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1415),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1437),
.Y(n_1579)
);

NAND2xp33_ASAP7_75t_L g1580 ( 
.A(n_1393),
.B(n_1474),
.Y(n_1580)
);

AOI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1427),
.A2(n_1396),
.B(n_1378),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1407),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1442),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1407),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1442),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1389),
.A2(n_1405),
.B(n_1395),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1405),
.Y(n_1587)
);

INVx8_ASAP7_75t_L g1588 ( 
.A(n_1383),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1376),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1469),
.A2(n_1402),
.B(n_1406),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1414),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1476),
.A2(n_1465),
.B1(n_1401),
.B2(n_1425),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1465),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1414),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1536),
.A2(n_1465),
.B1(n_1466),
.B2(n_1500),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1531),
.B(n_1497),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1505),
.B(n_1471),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1557),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_SL g1599 ( 
.A1(n_1524),
.A2(n_1394),
.B(n_1392),
.C(n_1395),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1537),
.B(n_1399),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1511),
.B(n_1477),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1512),
.A2(n_1500),
.B(n_1406),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1505),
.B(n_1471),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1508),
.B(n_1384),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1536),
.A2(n_1381),
.B1(n_1418),
.B2(n_1402),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1556),
.Y(n_1606)
);

OAI211xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1534),
.A2(n_1388),
.B(n_1385),
.C(n_1381),
.Y(n_1607)
);

BUFx4f_ASAP7_75t_SL g1608 ( 
.A(n_1513),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1578),
.B(n_1418),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1556),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1508),
.B(n_1418),
.Y(n_1611)
);

A2O1A1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1534),
.A2(n_1545),
.B(n_1548),
.C(n_1542),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1578),
.B(n_1385),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1547),
.B(n_1383),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1518),
.A2(n_1417),
.B(n_1363),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1547),
.B(n_1480),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1556),
.B(n_1398),
.Y(n_1617)
);

A2O1A1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1548),
.A2(n_1480),
.B(n_1410),
.C(n_1483),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1541),
.B(n_1546),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1518),
.A2(n_1480),
.B(n_1525),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_SL g1621 ( 
.A1(n_1529),
.A2(n_1590),
.B(n_1525),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1521),
.A2(n_1573),
.B(n_1543),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_SL g1623 ( 
.A1(n_1529),
.A2(n_1590),
.B(n_1569),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1521),
.A2(n_1573),
.B(n_1551),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1541),
.B(n_1546),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1562),
.B(n_1564),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1541),
.B(n_1546),
.Y(n_1627)
);

A2O1A1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1542),
.A2(n_1516),
.B(n_1577),
.C(n_1565),
.Y(n_1628)
);

AOI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1516),
.A2(n_1569),
.B1(n_1577),
.B2(n_1563),
.C(n_1568),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1558),
.B(n_1560),
.Y(n_1630)
);

O2A1O1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1551),
.A2(n_1580),
.B(n_1585),
.C(n_1583),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1511),
.B(n_1566),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1565),
.A2(n_1526),
.B(n_1522),
.C(n_1515),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1566),
.B(n_1558),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1567),
.B(n_1592),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1560),
.B(n_1582),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1582),
.B(n_1584),
.Y(n_1637)
);

OR2x6_ASAP7_75t_L g1638 ( 
.A(n_1526),
.B(n_1522),
.Y(n_1638)
);

OR2x6_ASAP7_75t_L g1639 ( 
.A(n_1540),
.B(n_1519),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1584),
.B(n_1553),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1586),
.A2(n_1585),
.B(n_1583),
.Y(n_1641)
);

CKINVDCx8_ASAP7_75t_R g1642 ( 
.A(n_1575),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1553),
.B(n_1514),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1503),
.B(n_1509),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1544),
.B(n_1535),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1586),
.A2(n_1583),
.B(n_1585),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1576),
.A2(n_1579),
.B1(n_1570),
.B2(n_1592),
.Y(n_1647)
);

A2O1A1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1532),
.A2(n_1559),
.B(n_1572),
.C(n_1570),
.Y(n_1648)
);

AO21x2_ASAP7_75t_L g1649 ( 
.A1(n_1539),
.A2(n_1552),
.B(n_1533),
.Y(n_1649)
);

AO21x2_ASAP7_75t_L g1650 ( 
.A1(n_1552),
.A2(n_1533),
.B(n_1549),
.Y(n_1650)
);

AND2x2_ASAP7_75t_SL g1651 ( 
.A(n_1559),
.B(n_1572),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1523),
.B(n_1528),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1506),
.A2(n_1510),
.B(n_1504),
.Y(n_1653)
);

AO22x2_ASAP7_75t_L g1654 ( 
.A1(n_1550),
.A2(n_1549),
.B1(n_1510),
.B2(n_1506),
.Y(n_1654)
);

INVx4_ASAP7_75t_L g1655 ( 
.A(n_1559),
.Y(n_1655)
);

O2A1O1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1574),
.A2(n_1563),
.B(n_1594),
.C(n_1576),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1653),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1643),
.B(n_1561),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1619),
.B(n_1520),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1639),
.B(n_1517),
.Y(n_1660)
);

BUFx2_ASAP7_75t_L g1661 ( 
.A(n_1654),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1632),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1606),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1643),
.B(n_1554),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1619),
.B(n_1625),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1625),
.B(n_1520),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1606),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1610),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_SL g1669 ( 
.A(n_1624),
.B(n_1507),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1629),
.B(n_1581),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1636),
.B(n_1538),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1627),
.B(n_1502),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_1651),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1650),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1610),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1627),
.B(n_1517),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1640),
.B(n_1637),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1637),
.B(n_1538),
.Y(n_1678)
);

NOR3xp33_ASAP7_75t_L g1679 ( 
.A(n_1622),
.B(n_1572),
.C(n_1559),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1607),
.A2(n_1579),
.B1(n_1576),
.B2(n_1532),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1638),
.B(n_1633),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1598),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1650),
.Y(n_1683)
);

BUFx5_ASAP7_75t_L g1684 ( 
.A(n_1651),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1650),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1612),
.B(n_1579),
.C(n_1591),
.Y(n_1686)
);

INVx4_ASAP7_75t_L g1687 ( 
.A(n_1655),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1630),
.B(n_1571),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1596),
.A2(n_1532),
.B1(n_1572),
.B2(n_1530),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1662),
.B(n_1626),
.Y(n_1690)
);

INVxp67_ASAP7_75t_SL g1691 ( 
.A(n_1674),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1662),
.B(n_1644),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_L g1693 ( 
.A(n_1686),
.B(n_1612),
.C(n_1628),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1667),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1658),
.B(n_1652),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1678),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1667),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1671),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1658),
.B(n_1628),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1677),
.B(n_1638),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1678),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1665),
.B(n_1604),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1670),
.A2(n_1599),
.B1(n_1656),
.B2(n_1631),
.C(n_1633),
.Y(n_1703)
);

NOR3xp33_ASAP7_75t_L g1704 ( 
.A(n_1686),
.B(n_1599),
.C(n_1615),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1667),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1664),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1657),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1668),
.Y(n_1708)
);

OAI321xp33_ASAP7_75t_L g1709 ( 
.A1(n_1670),
.A2(n_1638),
.A3(n_1620),
.B1(n_1646),
.B2(n_1641),
.C(n_1581),
.Y(n_1709)
);

INVx4_ASAP7_75t_L g1710 ( 
.A(n_1687),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1678),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1660),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1665),
.B(n_1671),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1668),
.Y(n_1714)
);

OAI221xp5_ASAP7_75t_L g1715 ( 
.A1(n_1669),
.A2(n_1647),
.B1(n_1618),
.B2(n_1602),
.C(n_1648),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1675),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1675),
.Y(n_1717)
);

NAND3xp33_ASAP7_75t_L g1718 ( 
.A(n_1679),
.B(n_1638),
.C(n_1648),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1657),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1675),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1663),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1657),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1677),
.B(n_1654),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1677),
.B(n_1654),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1665),
.B(n_1634),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1673),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1661),
.B(n_1649),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1680),
.A2(n_1618),
.B1(n_1613),
.B2(n_1605),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1661),
.B(n_1649),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1676),
.B(n_1645),
.Y(n_1730)
);

INVx3_ASAP7_75t_L g1731 ( 
.A(n_1660),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1664),
.B(n_1682),
.Y(n_1732)
);

AOI33xp33_ASAP7_75t_L g1733 ( 
.A1(n_1681),
.A2(n_1597),
.A3(n_1603),
.B1(n_1604),
.B2(n_1617),
.B3(n_1611),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1663),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1707),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1721),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1723),
.B(n_1661),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1721),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1699),
.B(n_1672),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1723),
.B(n_1681),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1727),
.B(n_1672),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1724),
.B(n_1681),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1693),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1707),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1719),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1734),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1724),
.B(n_1659),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1712),
.B(n_1659),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1727),
.B(n_1672),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1734),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1694),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1706),
.B(n_1659),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1719),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1726),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1694),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1710),
.B(n_1660),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1698),
.B(n_1732),
.Y(n_1757)
);

NAND2x1_ASAP7_75t_L g1758 ( 
.A(n_1726),
.B(n_1660),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1697),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1697),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1705),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1700),
.B(n_1673),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1705),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1710),
.B(n_1660),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1729),
.B(n_1688),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1710),
.B(n_1660),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1708),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1729),
.B(n_1688),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1700),
.B(n_1673),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1713),
.B(n_1666),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1708),
.B(n_1666),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1714),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1714),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1712),
.B(n_1666),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1756),
.Y(n_1775)
);

INVxp67_ASAP7_75t_SL g1776 ( 
.A(n_1743),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1755),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1756),
.Y(n_1778)
);

O2A1O1Ixp5_ASAP7_75t_L g1779 ( 
.A1(n_1758),
.A2(n_1718),
.B(n_1728),
.C(n_1712),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1743),
.B(n_1733),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1755),
.Y(n_1781)
);

NOR2xp67_ASAP7_75t_SL g1782 ( 
.A(n_1762),
.B(n_1715),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1772),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1772),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1739),
.B(n_1725),
.Y(n_1785)
);

NAND2x1_ASAP7_75t_L g1786 ( 
.A(n_1756),
.B(n_1731),
.Y(n_1786)
);

OR2x2_ASAP7_75t_SL g1787 ( 
.A(n_1739),
.B(n_1692),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1735),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1736),
.Y(n_1789)
);

AO21x1_ASAP7_75t_L g1790 ( 
.A1(n_1758),
.A2(n_1704),
.B(n_1669),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1765),
.B(n_1725),
.Y(n_1791)
);

INVxp67_ASAP7_75t_L g1792 ( 
.A(n_1754),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1740),
.B(n_1731),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1754),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1765),
.B(n_1702),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1736),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1740),
.B(n_1731),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1756),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1757),
.B(n_1703),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1768),
.B(n_1692),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1735),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1737),
.A2(n_1679),
.B1(n_1680),
.B2(n_1635),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1757),
.B(n_1695),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1738),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1752),
.B(n_1690),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_1764),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1742),
.B(n_1730),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1738),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1752),
.B(n_1690),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1742),
.B(n_1737),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1764),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1737),
.B(n_1730),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1764),
.B(n_1696),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1746),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1764),
.B(n_1696),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1766),
.B(n_1701),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1766),
.A2(n_1709),
.B(n_1527),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1787),
.B(n_1768),
.Y(n_1818)
);

OR2x6_ASAP7_75t_L g1819 ( 
.A(n_1817),
.B(n_1595),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1787),
.B(n_1741),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1776),
.B(n_1747),
.Y(n_1821)
);

NOR2x1_ASAP7_75t_L g1822 ( 
.A(n_1799),
.B(n_1601),
.Y(n_1822)
);

NOR2x1_ASAP7_75t_R g1823 ( 
.A(n_1780),
.B(n_1527),
.Y(n_1823)
);

NOR2x1_ASAP7_75t_L g1824 ( 
.A(n_1777),
.B(n_1781),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1782),
.B(n_1747),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1810),
.B(n_1811),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1782),
.B(n_1747),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1810),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1785),
.B(n_1741),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1792),
.B(n_1762),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1811),
.B(n_1766),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1779),
.A2(n_1689),
.B(n_1685),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1785),
.B(n_1749),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1775),
.B(n_1766),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1811),
.B(n_1769),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1803),
.B(n_1769),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1790),
.B(n_1684),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1811),
.B(n_1748),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1790),
.B(n_1684),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1802),
.B(n_1642),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1807),
.B(n_1748),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1800),
.B(n_1749),
.Y(n_1842)
);

INVxp67_ASAP7_75t_L g1843 ( 
.A(n_1794),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1789),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1789),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1807),
.B(n_1748),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1788),
.Y(n_1847)
);

NAND4xp25_ASAP7_75t_L g1848 ( 
.A(n_1802),
.B(n_1689),
.C(n_1600),
.D(n_1617),
.Y(n_1848)
);

OAI31xp33_ASAP7_75t_L g1849 ( 
.A1(n_1798),
.A2(n_1673),
.A3(n_1674),
.B(n_1774),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1812),
.B(n_1774),
.Y(n_1850)
);

AOI221xp5_ASAP7_75t_SL g1851 ( 
.A1(n_1806),
.A2(n_1683),
.B1(n_1685),
.B2(n_1771),
.C(n_1774),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1796),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1800),
.B(n_1771),
.Y(n_1853)
);

INVx1_ASAP7_75t_SL g1854 ( 
.A(n_1822),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1824),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1844),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_SL g1857 ( 
.A(n_1823),
.B(n_1840),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1844),
.Y(n_1858)
);

NAND3xp33_ASAP7_75t_L g1859 ( 
.A(n_1843),
.B(n_1781),
.C(n_1777),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1837),
.A2(n_1775),
.B1(n_1778),
.B2(n_1812),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1839),
.A2(n_1778),
.B1(n_1805),
.B2(n_1809),
.Y(n_1861)
);

AOI211xp5_ASAP7_75t_SL g1862 ( 
.A1(n_1825),
.A2(n_1608),
.B(n_1783),
.C(n_1784),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1821),
.B(n_1791),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1835),
.B(n_1813),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1830),
.B(n_1795),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1845),
.Y(n_1866)
);

AOI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1832),
.A2(n_1784),
.B1(n_1783),
.B2(n_1814),
.C(n_1808),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1836),
.B(n_1795),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1845),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1835),
.B(n_1813),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_SL g1871 ( 
.A1(n_1848),
.A2(n_1816),
.B(n_1815),
.Y(n_1871)
);

OAI21xp33_ASAP7_75t_SL g1872 ( 
.A1(n_1827),
.A2(n_1797),
.B(n_1793),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1826),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1828),
.B(n_1818),
.Y(n_1874)
);

AOI31xp33_ASAP7_75t_L g1875 ( 
.A1(n_1818),
.A2(n_1791),
.A3(n_1815),
.B(n_1816),
.Y(n_1875)
);

INVx1_ASAP7_75t_SL g1876 ( 
.A(n_1820),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1852),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1852),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1820),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1867),
.A2(n_1854),
.B1(n_1859),
.B2(n_1876),
.C(n_1879),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1873),
.B(n_1828),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1855),
.Y(n_1882)
);

OAI31xp33_ASAP7_75t_L g1883 ( 
.A1(n_1862),
.A2(n_1849),
.A3(n_1834),
.B(n_1826),
.Y(n_1883)
);

OAI221xp5_ASAP7_75t_SL g1884 ( 
.A1(n_1871),
.A2(n_1819),
.B1(n_1851),
.B2(n_1842),
.C(n_1829),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1873),
.B(n_1841),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1875),
.A2(n_1819),
.B1(n_1863),
.B2(n_1874),
.Y(n_1886)
);

AOI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1857),
.A2(n_1819),
.B(n_1834),
.Y(n_1887)
);

O2A1O1Ixp33_ASAP7_75t_L g1888 ( 
.A1(n_1860),
.A2(n_1819),
.B(n_1847),
.C(n_1834),
.Y(n_1888)
);

OAI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1861),
.A2(n_1831),
.B(n_1842),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1874),
.Y(n_1890)
);

NAND4xp25_ASAP7_75t_SL g1891 ( 
.A(n_1872),
.B(n_1829),
.C(n_1833),
.D(n_1853),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1856),
.Y(n_1892)
);

AOI211xp5_ASAP7_75t_L g1893 ( 
.A1(n_1863),
.A2(n_1831),
.B(n_1853),
.C(n_1833),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1864),
.B(n_1841),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1865),
.B(n_1642),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1864),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1868),
.B(n_1846),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1870),
.B(n_1846),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1856),
.A2(n_1786),
.B(n_1796),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1890),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1896),
.B(n_1870),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1885),
.Y(n_1902)
);

NAND4xp25_ASAP7_75t_L g1903 ( 
.A(n_1880),
.B(n_1878),
.C(n_1877),
.D(n_1869),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1895),
.B(n_1513),
.Y(n_1904)
);

AOI211xp5_ASAP7_75t_L g1905 ( 
.A1(n_1884),
.A2(n_1866),
.B(n_1858),
.C(n_1869),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1894),
.B(n_1858),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1886),
.A2(n_1866),
.B(n_1847),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1882),
.B(n_1850),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1898),
.Y(n_1909)
);

INVxp67_ASAP7_75t_SL g1910 ( 
.A(n_1882),
.Y(n_1910)
);

AOI322xp5_ASAP7_75t_L g1911 ( 
.A1(n_1895),
.A2(n_1850),
.A3(n_1838),
.B1(n_1786),
.B2(n_1793),
.C1(n_1797),
.C2(n_1691),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1881),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1910),
.A2(n_1888),
.B(n_1891),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1901),
.B(n_1893),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1910),
.Y(n_1915)
);

NOR3xp33_ASAP7_75t_L g1916 ( 
.A(n_1904),
.B(n_1887),
.C(n_1889),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1900),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1911),
.B(n_1883),
.Y(n_1918)
);

NAND3xp33_ASAP7_75t_SL g1919 ( 
.A(n_1905),
.B(n_1897),
.C(n_1899),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1908),
.Y(n_1920)
);

OAI211xp5_ASAP7_75t_SL g1921 ( 
.A1(n_1902),
.A2(n_1892),
.B(n_1801),
.C(n_1788),
.Y(n_1921)
);

NOR3xp33_ASAP7_75t_L g1922 ( 
.A(n_1903),
.B(n_1838),
.C(n_1801),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1909),
.B(n_1804),
.Y(n_1923)
);

AND4x1_ASAP7_75t_L g1924 ( 
.A(n_1913),
.B(n_1907),
.C(n_1912),
.D(n_1513),
.Y(n_1924)
);

AOI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1918),
.A2(n_1907),
.B1(n_1906),
.B2(n_1804),
.Y(n_1925)
);

AOI222xp33_ASAP7_75t_L g1926 ( 
.A1(n_1919),
.A2(n_1814),
.B1(n_1808),
.B2(n_1683),
.C1(n_1801),
.C2(n_1788),
.Y(n_1926)
);

NAND4xp75_ASAP7_75t_L g1927 ( 
.A(n_1915),
.B(n_1513),
.C(n_1597),
.D(n_1603),
.Y(n_1927)
);

OAI21xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1917),
.A2(n_1614),
.B(n_1616),
.Y(n_1928)
);

AOI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1925),
.A2(n_1916),
.B1(n_1914),
.B2(n_1922),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1928),
.A2(n_1922),
.B1(n_1920),
.B2(n_1923),
.Y(n_1930)
);

AOI221xp5_ASAP7_75t_L g1931 ( 
.A1(n_1924),
.A2(n_1921),
.B1(n_1746),
.B2(n_1750),
.C(n_1751),
.Y(n_1931)
);

AOI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1926),
.A2(n_1750),
.B1(n_1760),
.B2(n_1759),
.C(n_1773),
.Y(n_1932)
);

AOI221xp5_ASAP7_75t_SL g1933 ( 
.A1(n_1927),
.A2(n_1773),
.B1(n_1751),
.B2(n_1767),
.C(n_1763),
.Y(n_1933)
);

OAI221xp5_ASAP7_75t_SL g1934 ( 
.A1(n_1925),
.A2(n_1593),
.B1(n_1770),
.B2(n_1587),
.C(n_1753),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1930),
.Y(n_1935)
);

NOR3xp33_ASAP7_75t_L g1936 ( 
.A(n_1929),
.B(n_1593),
.C(n_1655),
.Y(n_1936)
);

OAI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1934),
.A2(n_1735),
.B1(n_1744),
.B2(n_1745),
.Y(n_1937)
);

NAND4xp75_ASAP7_75t_L g1938 ( 
.A(n_1933),
.B(n_1761),
.C(n_1759),
.D(n_1760),
.Y(n_1938)
);

NAND2x1p5_ASAP7_75t_L g1939 ( 
.A(n_1931),
.B(n_1593),
.Y(n_1939)
);

XNOR2xp5_ASAP7_75t_L g1940 ( 
.A(n_1935),
.B(n_1932),
.Y(n_1940)
);

OAI321xp33_ASAP7_75t_L g1941 ( 
.A1(n_1939),
.A2(n_1587),
.A3(n_1609),
.B1(n_1770),
.B2(n_1589),
.C(n_1763),
.Y(n_1941)
);

OAI221xp5_ASAP7_75t_L g1942 ( 
.A1(n_1936),
.A2(n_1555),
.B1(n_1744),
.B2(n_1753),
.C(n_1745),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1940),
.Y(n_1943)
);

OAI22x1_ASAP7_75t_L g1944 ( 
.A1(n_1943),
.A2(n_1942),
.B1(n_1941),
.B2(n_1938),
.Y(n_1944)
);

XNOR2xp5_ASAP7_75t_L g1945 ( 
.A(n_1944),
.B(n_1937),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1944),
.B(n_1744),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1946),
.A2(n_1753),
.B1(n_1745),
.B2(n_1767),
.Y(n_1947)
);

NOR2x1_ASAP7_75t_L g1948 ( 
.A(n_1945),
.B(n_1761),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1948),
.A2(n_1588),
.B(n_1621),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1947),
.A2(n_1588),
.B(n_1623),
.Y(n_1950)
);

AOI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1949),
.A2(n_1701),
.B1(n_1711),
.B2(n_1555),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1951),
.B(n_1950),
.Y(n_1952)
);

NAND2xp33_ASAP7_75t_L g1953 ( 
.A(n_1952),
.B(n_1588),
.Y(n_1953)
);

AOI221xp5_ASAP7_75t_L g1954 ( 
.A1(n_1953),
.A2(n_1722),
.B1(n_1720),
.B2(n_1717),
.C(n_1716),
.Y(n_1954)
);

AOI211xp5_ASAP7_75t_L g1955 ( 
.A1(n_1954),
.A2(n_1555),
.B(n_1614),
.C(n_1616),
.Y(n_1955)
);


endmodule