module fake_jpeg_14602_n_138 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_30),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_5),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_5),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_10),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_24),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_55),
.Y(n_78)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_18),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_11),
.Y(n_63)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_68)
);

A2O1A1O1Ixp25_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_69),
.B(n_64),
.C(n_52),
.D(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_31),
.B(n_11),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_73),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_37),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_26),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_81),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_26),
.B1(n_67),
.B2(n_47),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_61),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_66),
.B1(n_57),
.B2(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_88),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_69),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_50),
.C(n_54),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_50),
.C(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_48),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_58),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_100),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_73),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_101),
.C(n_106),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_79),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_82),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_86),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_72),
.C(n_80),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_75),
.C(n_74),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_74),
.C(n_87),
.Y(n_112)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_97),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_121),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_124),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_112),
.B1(n_116),
.B2(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_117),
.B(n_108),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_129),
.B(n_128),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_109),
.B(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_131),
.B(n_134),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_135),
.Y(n_138)
);


endmodule