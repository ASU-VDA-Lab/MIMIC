module real_jpeg_32330_n_25 (n_17, n_8, n_0, n_21, n_2, n_185, n_180, n_10, n_175, n_9, n_178, n_186, n_12, n_24, n_176, n_6, n_183, n_177, n_179, n_23, n_11, n_14, n_7, n_22, n_18, n_3, n_174, n_5, n_4, n_173, n_181, n_1, n_182, n_20, n_19, n_184, n_16, n_15, n_13, n_25);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_185;
input n_180;
input n_10;
input n_175;
input n_9;
input n_178;
input n_186;
input n_12;
input n_24;
input n_176;
input n_6;
input n_183;
input n_177;
input n_179;
input n_23;
input n_11;
input n_14;
input n_7;
input n_22;
input n_18;
input n_3;
input n_174;
input n_5;
input n_4;
input n_173;
input n_181;
input n_1;
input n_182;
input n_20;
input n_19;
input n_184;
input n_16;
input n_15;
input n_13;

output n_25;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_0),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_1),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_1),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_2),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_2),
.B(n_41),
.Y(n_171)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_4),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_5),
.B(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_5),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_6),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_6),
.B(n_104),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_7),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_8),
.B(n_63),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_9),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_SL g70 ( 
.A1(n_11),
.A2(n_58),
.B(n_62),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_11),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_12),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_12),
.B(n_109),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_13),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_13),
.B(n_155),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_15),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_15),
.A2(n_95),
.A3(n_97),
.B1(n_102),
.B2(n_127),
.C1(n_129),
.C2(n_184),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_16),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_58),
.C(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_17),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_17),
.B(n_116),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_19),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_19),
.B(n_135),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_20),
.B(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_22),
.B(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_24),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_24),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_36),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_48),
.B(n_171),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_47),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_137),
.B(n_157),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_132),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI31xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_88),
.A3(n_114),
.B(n_122),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_81),
.C(n_82),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_73),
.B(n_80),
.Y(n_54)
);

OAI322xp33_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_64),
.A3(n_69),
.B1(n_70),
.B2(n_71),
.C1(n_72),
.C2(n_173),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_175),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_79),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_101),
.C(n_108),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_123),
.B(n_126),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_108),
.C(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_180),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OA21x2_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_145),
.C(n_149),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_166),
.C(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp67_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

OAI322xp33_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_151),
.A3(n_165),
.B1(n_168),
.B2(n_169),
.C1(n_170),
.C2(n_186),
.Y(n_164)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI321xp33_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_159),
.A3(n_160),
.B1(n_161),
.B2(n_164),
.C(n_185),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_174),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_176),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_177),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_178),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_179),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_181),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_182),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_183),
.Y(n_117)
);


endmodule