module fake_ibex_613_n_943 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_943);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_943;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_732;
wire n_673;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_857;
wire n_849;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_560;
wire n_429;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_566;
wire n_484;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_444;
wire n_200;
wire n_562;
wire n_506;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_905;
wire n_410;
wire n_762;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_927;
wire n_684;
wire n_775;
wire n_934;
wire n_784;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_10),
.Y(n_172)
);

BUFx2_ASAP7_75t_SL g173 ( 
.A(n_8),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_60),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_139),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_14),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_83),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_5),
.Y(n_180)
);

NOR2xp67_ASAP7_75t_L g181 ( 
.A(n_50),
.B(n_102),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_46),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_86),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_147),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_85),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_75),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_137),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_27),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_92),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_71),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_37),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_31),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_78),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_91),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_67),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_132),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_55),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_155),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_66),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_40),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_65),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_97),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_70),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_136),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_36),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_30),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_62),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_53),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_38),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_90),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_73),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_74),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_120),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_54),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_115),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_166),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_162),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_98),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_109),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_34),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_106),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_129),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_64),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_43),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_142),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_68),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_88),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_42),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_151),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_148),
.B(n_28),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_131),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_57),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_49),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_79),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_42),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_87),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_37),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_118),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_35),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_14),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_41),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_2),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_108),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_52),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_128),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_58),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_161),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_156),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_105),
.B(n_12),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_51),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_63),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_122),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_80),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_158),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_39),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_123),
.B(n_145),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_157),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_61),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_76),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_121),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_96),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_150),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_23),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_140),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_59),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_29),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_27),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_100),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_198),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_231),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_196),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_0),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_195),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

AND2x4_ASAP7_75t_L g288 ( 
.A(n_239),
.B(n_1),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_195),
.A2(n_94),
.B(n_169),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_190),
.Y(n_290)
);

BUFx8_ASAP7_75t_L g291 ( 
.A(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_248),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_259),
.Y(n_293)
);

AND2x4_ASAP7_75t_L g294 ( 
.A(n_215),
.B(n_3),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_172),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_250),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_201),
.A2(n_93),
.B(n_168),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_179),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_172),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_179),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_178),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_201),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_224),
.Y(n_304)
);

BUFx8_ASAP7_75t_SL g305 ( 
.A(n_204),
.Y(n_305)
);

OA21x2_ASAP7_75t_L g306 ( 
.A1(n_224),
.A2(n_95),
.B(n_167),
.Y(n_306)
);

AND2x4_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_4),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_179),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_179),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_232),
.B(n_6),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_229),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_6),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_223),
.B(n_7),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_232),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_229),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_238),
.B(n_9),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_238),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_178),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_318)
);

CKINVDCx6p67_ASAP7_75t_R g319 ( 
.A(n_198),
.Y(n_319)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_205),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_240),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_205),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_205),
.Y(n_323)
);

BUFx8_ASAP7_75t_SL g324 ( 
.A(n_204),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_240),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_205),
.Y(n_326)
);

BUFx12f_ASAP7_75t_L g327 ( 
.A(n_183),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g328 ( 
.A(n_247),
.B(n_47),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_247),
.B(n_276),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_225),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_180),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_170),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_225),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_171),
.Y(n_334)
);

OA21x2_ASAP7_75t_L g335 ( 
.A1(n_174),
.A2(n_101),
.B(n_165),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_266),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_277),
.B(n_11),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_225),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_177),
.Y(n_339)
);

BUFx12f_ASAP7_75t_L g340 ( 
.A(n_183),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_180),
.B(n_15),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_182),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_184),
.B(n_15),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_225),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_256),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_175),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_185),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g348 ( 
.A(n_199),
.B(n_48),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_256),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_182),
.B(n_16),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_173),
.B(n_16),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_207),
.B(n_17),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_271),
.B(n_18),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_208),
.Y(n_355)
);

NOR2x1_ASAP7_75t_L g356 ( 
.A(n_209),
.B(n_56),
.Y(n_356)
);

BUFx8_ASAP7_75t_L g357 ( 
.A(n_260),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_256),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_210),
.B(n_18),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_344),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_344),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_344),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_345),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_345),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_316),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_286),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_345),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_345),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_288),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_298),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_298),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_288),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_298),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_282),
.B(n_249),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_342),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_288),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_303),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_295),
.B(n_194),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_298),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_304),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_298),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_304),
.Y(n_386)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_294),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_308),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_327),
.Y(n_389)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_328),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

INVxp33_ASAP7_75t_SL g393 ( 
.A(n_293),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_294),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_314),
.B(n_273),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_291),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_294),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_291),
.Y(n_398)
);

AND2x6_ASAP7_75t_L g399 ( 
.A(n_313),
.B(n_211),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_307),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_307),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_307),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_337),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_319),
.B(n_212),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_308),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_346),
.B(n_186),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_343),
.A2(n_352),
.B1(n_353),
.B2(n_310),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_329),
.B(n_193),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_308),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_309),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_348),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_327),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_340),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_284),
.B(n_213),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_280),
.B(n_218),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_309),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_287),
.B(n_217),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_309),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_319),
.B(n_235),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_299),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_309),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_309),
.Y(n_423)
);

AOI21x1_ASAP7_75t_L g424 ( 
.A1(n_297),
.A2(n_222),
.B(n_221),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_352),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_322),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_322),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_322),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_281),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_322),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_322),
.Y(n_432)
);

NOR2x1p5_ASAP7_75t_L g433 ( 
.A(n_293),
.B(n_246),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_329),
.B(n_187),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_281),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_315),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_323),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_313),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_L g439 ( 
.A(n_348),
.B(n_328),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_323),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_329),
.B(n_189),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_315),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_317),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_341),
.Y(n_444)
);

AND2x2_ASAP7_75t_SL g445 ( 
.A(n_285),
.B(n_193),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_323),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_347),
.B(n_192),
.Y(n_447)
);

AND3x2_ASAP7_75t_L g448 ( 
.A(n_305),
.B(n_234),
.C(n_241),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_317),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_340),
.Y(n_450)
);

OAI22xp33_ASAP7_75t_L g451 ( 
.A1(n_351),
.A2(n_214),
.B1(n_278),
.B2(n_176),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_L g452 ( 
.A(n_348),
.B(n_197),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_290),
.B(n_251),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_323),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_321),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_355),
.B(n_253),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_L g457 ( 
.A(n_348),
.B(n_200),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_321),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_SL g459 ( 
.A(n_351),
.B(n_176),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_305),
.Y(n_460)
);

NAND3xp33_ASAP7_75t_L g461 ( 
.A(n_312),
.B(n_230),
.C(n_233),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_325),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_326),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_325),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_L g465 ( 
.A(n_348),
.B(n_202),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_332),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_332),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_326),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_292),
.B(n_203),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_296),
.B(n_206),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_301),
.A2(n_242),
.B1(n_258),
.B2(n_262),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_L g472 ( 
.A(n_328),
.B(n_216),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_334),
.B(n_219),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_328),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_334),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_330),
.Y(n_476)
);

INVxp33_ASAP7_75t_L g477 ( 
.A(n_324),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_336),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_330),
.Y(n_479)
);

NOR2x1p5_ASAP7_75t_L g480 ( 
.A(n_324),
.B(n_214),
.Y(n_480)
);

INVxp33_ASAP7_75t_L g481 ( 
.A(n_350),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_339),
.B(n_236),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_339),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_360),
.A2(n_328),
.B1(n_359),
.B2(n_356),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_478),
.B(n_357),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_478),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_478),
.B(n_357),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_444),
.B(n_357),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_462),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_226),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_227),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_462),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_396),
.B(n_228),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_462),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_378),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_360),
.A2(n_362),
.B1(n_368),
.B2(n_375),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_426),
.B(n_278),
.Y(n_497)
);

NOR3xp33_ASAP7_75t_L g498 ( 
.A(n_451),
.B(n_283),
.C(n_318),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_362),
.A2(n_328),
.B1(n_289),
.B2(n_306),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_453),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_456),
.B(n_254),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_453),
.B(n_263),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_445),
.A2(n_279),
.B1(n_188),
.B2(n_191),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_445),
.A2(n_279),
.B1(n_191),
.B2(n_264),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_398),
.B(n_265),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_416),
.B(n_268),
.Y(n_506)
);

A2O1A1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_400),
.A2(n_275),
.B(n_237),
.C(n_243),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_430),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_377),
.B(n_220),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_407),
.B(n_245),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_404),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_403),
.B(n_255),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_368),
.A2(n_289),
.B1(n_306),
.B2(n_270),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_372),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_473),
.B(n_257),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_434),
.B(n_272),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_433),
.B(n_264),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g518 ( 
.A(n_389),
.B(n_302),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_412),
.B(n_289),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_375),
.A2(n_306),
.B1(n_335),
.B2(n_320),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_420),
.B(n_421),
.Y(n_521)
);

NOR3xp33_ASAP7_75t_L g522 ( 
.A(n_459),
.B(n_181),
.C(n_267),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_425),
.B(n_300),
.Y(n_523)
);

O2A1O1Ixp5_ASAP7_75t_L g524 ( 
.A1(n_424),
.A2(n_300),
.B(n_320),
.C(n_349),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_382),
.B(n_19),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_435),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_435),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_441),
.B(n_300),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_408),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_408),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_399),
.A2(n_401),
.B1(n_402),
.B2(n_387),
.Y(n_531)
);

AO22x2_ASAP7_75t_L g532 ( 
.A1(n_375),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_532)
);

NOR3xp33_ASAP7_75t_L g533 ( 
.A(n_382),
.B(n_20),
.C(n_21),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_420),
.Y(n_534)
);

INVx8_ASAP7_75t_L g535 ( 
.A(n_387),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_411),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_387),
.B(n_300),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_379),
.A2(n_358),
.B1(n_354),
.B2(n_349),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_395),
.B(n_69),
.Y(n_539)
);

NAND2x1p5_ASAP7_75t_L g540 ( 
.A(n_450),
.B(n_358),
.Y(n_540)
);

NOR2xp67_ASAP7_75t_L g541 ( 
.A(n_389),
.B(n_413),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_482),
.B(n_330),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_482),
.B(n_333),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_450),
.B(n_22),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_399),
.A2(n_358),
.B1(n_354),
.B2(n_349),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_408),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_464),
.B(n_338),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_393),
.B(n_349),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_379),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_466),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_379),
.A2(n_349),
.B1(n_338),
.B2(n_333),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_415),
.B(n_418),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_L g553 ( 
.A(n_399),
.B(n_338),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_406),
.B(n_113),
.Y(n_554)
);

NOR3xp33_ASAP7_75t_L g555 ( 
.A(n_461),
.B(n_24),
.C(n_25),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_394),
.B(n_333),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_474),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_413),
.B(n_24),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_470),
.B(n_114),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_480),
.B(n_438),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_466),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_438),
.B(n_333),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_439),
.A2(n_112),
.B(n_164),
.Y(n_563)
);

NAND3xp33_ASAP7_75t_SL g564 ( 
.A(n_471),
.B(n_26),
.C(n_28),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_369),
.Y(n_565)
);

NAND2x1p5_ASAP7_75t_L g566 ( 
.A(n_397),
.B(n_30),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_414),
.B(n_31),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_467),
.B(n_32),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_390),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_447),
.B(n_117),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_475),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_475),
.Y(n_572)
);

BUFx6f_ASAP7_75t_SL g573 ( 
.A(n_477),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_483),
.Y(n_574)
);

INVx8_ASAP7_75t_L g575 ( 
.A(n_390),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_549),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_535),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_519),
.A2(n_465),
.B(n_452),
.Y(n_578)
);

A2O1A1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_514),
.A2(n_452),
.B(n_457),
.C(n_465),
.Y(n_579)
);

BUFx8_ASAP7_75t_SL g580 ( 
.A(n_573),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_499),
.A2(n_556),
.B(n_513),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_514),
.B(n_380),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_534),
.B(n_448),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_535),
.B(n_474),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_495),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_521),
.B(n_460),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_552),
.B(n_380),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_497),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_496),
.A2(n_504),
.B1(n_503),
.B2(n_531),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_513),
.A2(n_472),
.B(n_384),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_566),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_500),
.B(n_381),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_523),
.A2(n_381),
.B(n_384),
.Y(n_593)
);

AO21x1_ASAP7_75t_L g594 ( 
.A1(n_563),
.A2(n_566),
.B(n_522),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_544),
.Y(n_595)
);

AND2x6_ASAP7_75t_L g596 ( 
.A(n_544),
.B(n_386),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_488),
.B(n_392),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_565),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_510),
.B(n_436),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_511),
.B(n_436),
.Y(n_600)
);

BUFx12f_ASAP7_75t_L g601 ( 
.A(n_560),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_520),
.A2(n_442),
.B(n_443),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_520),
.A2(n_442),
.B(n_443),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_562),
.A2(n_449),
.B(n_455),
.Y(n_604)
);

NOR3xp33_ASAP7_75t_L g605 ( 
.A(n_498),
.B(n_460),
.C(n_449),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_573),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_512),
.A2(n_455),
.B(n_458),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_529),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_530),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_485),
.B(n_36),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_548),
.B(n_536),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_491),
.B(n_502),
.Y(n_612)
);

AND2x6_ASAP7_75t_SL g613 ( 
.A(n_560),
.B(n_38),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_515),
.A2(n_479),
.B(n_476),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_487),
.B(n_41),
.Y(n_615)
);

NOR2xp67_ASAP7_75t_L g616 ( 
.A(n_541),
.B(n_43),
.Y(n_616)
);

O2A1O1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_507),
.A2(n_361),
.B(n_371),
.C(n_370),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_533),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_575),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_546),
.Y(n_620)
);

NOR2x1_ASAP7_75t_R g621 ( 
.A(n_517),
.B(n_44),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_490),
.B(n_44),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_568),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_574),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_516),
.B(n_45),
.Y(n_625)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_522),
.B(n_363),
.C(n_364),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_524),
.A2(n_468),
.B(n_463),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_525),
.A2(n_365),
.B1(n_367),
.B2(n_366),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_501),
.B(n_72),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_550),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_575),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_561),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_518),
.A2(n_454),
.B1(n_446),
.B2(n_440),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_484),
.A2(n_572),
.B(n_526),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_533),
.B(n_437),
.C(n_432),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_506),
.B(n_77),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_493),
.B(n_81),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_560),
.B(n_431),
.Y(n_638)
);

O2A1O1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_564),
.A2(n_429),
.B(n_428),
.C(n_427),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_564),
.A2(n_428),
.B1(n_427),
.B2(n_423),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_509),
.B(n_99),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_558),
.B(n_104),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_489),
.A2(n_492),
.B(n_494),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_553),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_567),
.B(n_107),
.Y(n_645)
);

BUFx4f_ASAP7_75t_L g646 ( 
.A(n_540),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_508),
.A2(n_422),
.B(n_373),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_540),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_527),
.A2(n_388),
.B(n_417),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_571),
.A2(n_385),
.B1(n_410),
.B2(n_409),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_575),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_505),
.B(n_111),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_542),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_570),
.A2(n_405),
.B(n_391),
.C(n_383),
.Y(n_654)
);

INVx3_ASAP7_75t_SL g655 ( 
.A(n_532),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_557),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_537),
.A2(n_376),
.B(n_374),
.Y(n_657)
);

O2A1O1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_555),
.A2(n_373),
.B(n_124),
.C(n_127),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_543),
.A2(n_419),
.B(n_130),
.Y(n_659)
);

OAI21xp33_ASAP7_75t_SL g660 ( 
.A1(n_587),
.A2(n_571),
.B(n_563),
.Y(n_660)
);

O2A1O1Ixp5_ASAP7_75t_L g661 ( 
.A1(n_594),
.A2(n_581),
.B(n_611),
.C(n_629),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_585),
.Y(n_662)
);

AO31x2_ASAP7_75t_L g663 ( 
.A1(n_590),
.A2(n_547),
.A3(n_539),
.B(n_554),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_627),
.A2(n_603),
.B(n_602),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_624),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_577),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_579),
.A2(n_597),
.B(n_643),
.Y(n_667)
);

AO31x2_ASAP7_75t_L g668 ( 
.A1(n_654),
.A2(n_559),
.A3(n_528),
.B(n_532),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_634),
.A2(n_545),
.B(n_551),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_607),
.A2(n_551),
.B(n_538),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_619),
.Y(n_671)
);

AOI21xp33_ASAP7_75t_L g672 ( 
.A1(n_658),
.A2(n_569),
.B(n_419),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_596),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_593),
.A2(n_419),
.B(n_135),
.Y(n_674)
);

AO21x2_ASAP7_75t_L g675 ( 
.A1(n_635),
.A2(n_133),
.B(n_138),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_655),
.A2(n_143),
.B1(n_144),
.B2(n_149),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_612),
.A2(n_153),
.B(n_154),
.C(n_159),
.Y(n_677)
);

INVx5_ASAP7_75t_L g678 ( 
.A(n_619),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_601),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_622),
.A2(n_636),
.B(n_618),
.C(n_617),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_630),
.Y(n_681)
);

OA22x2_ASAP7_75t_L g682 ( 
.A1(n_615),
.A2(n_595),
.B1(n_589),
.B2(n_586),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_592),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_632),
.A2(n_618),
.B(n_639),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_588),
.B(n_583),
.Y(n_685)
);

AOI211x1_ASAP7_75t_L g686 ( 
.A1(n_626),
.A2(n_625),
.B(n_599),
.C(n_610),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_596),
.B(n_600),
.Y(n_687)
);

NOR2x1p5_ASAP7_75t_L g688 ( 
.A(n_606),
.B(n_591),
.Y(n_688)
);

OAI21x1_ASAP7_75t_SL g689 ( 
.A1(n_652),
.A2(n_641),
.B(n_598),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_591),
.B(n_638),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_645),
.A2(n_642),
.B1(n_615),
.B2(n_637),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_596),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_600),
.B(n_620),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_638),
.B(n_631),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_608),
.Y(n_695)
);

AO31x2_ASAP7_75t_L g696 ( 
.A1(n_650),
.A2(n_659),
.A3(n_628),
.B(n_614),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_580),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_638),
.B(n_609),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_640),
.A2(n_653),
.B(n_604),
.Y(n_699)
);

AO31x2_ASAP7_75t_L g700 ( 
.A1(n_647),
.A2(n_649),
.A3(n_657),
.B(n_576),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_637),
.A2(n_646),
.B1(n_616),
.B2(n_648),
.Y(n_701)
);

AO21x2_ASAP7_75t_L g702 ( 
.A1(n_633),
.A2(n_644),
.B(n_584),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_656),
.A2(n_651),
.B(n_621),
.C(n_613),
.Y(n_703)
);

OAI21x1_ASAP7_75t_SL g704 ( 
.A1(n_594),
.A2(n_597),
.B(n_563),
.Y(n_704)
);

AO31x2_ASAP7_75t_L g705 ( 
.A1(n_594),
.A2(n_581),
.A3(n_590),
.B(n_578),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_581),
.A2(n_590),
.B(n_578),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_577),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_655),
.A2(n_587),
.B1(n_582),
.B2(n_623),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_577),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_585),
.Y(n_710)
);

AO31x2_ASAP7_75t_L g711 ( 
.A1(n_594),
.A2(n_581),
.A3(n_590),
.B(n_578),
.Y(n_711)
);

AO31x2_ASAP7_75t_L g712 ( 
.A1(n_594),
.A2(n_581),
.A3(n_590),
.B(n_578),
.Y(n_712)
);

AO31x2_ASAP7_75t_L g713 ( 
.A1(n_594),
.A2(n_581),
.A3(n_590),
.B(n_578),
.Y(n_713)
);

AO31x2_ASAP7_75t_L g714 ( 
.A1(n_594),
.A2(n_581),
.A3(n_590),
.B(n_578),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_577),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_624),
.Y(n_716)
);

BUFx4f_ASAP7_75t_L g717 ( 
.A(n_577),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_655),
.A2(n_587),
.B1(n_582),
.B2(n_623),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_577),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_587),
.B(n_495),
.Y(n_720)
);

AOI221x1_ASAP7_75t_L g721 ( 
.A1(n_581),
.A2(n_522),
.B1(n_532),
.B2(n_533),
.C(n_605),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_624),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_624),
.Y(n_723)
);

OAI22x1_ASAP7_75t_L g724 ( 
.A1(n_655),
.A2(n_585),
.B1(n_495),
.B2(n_480),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_587),
.B(n_495),
.Y(n_725)
);

OAI21xp5_ASAP7_75t_L g726 ( 
.A1(n_581),
.A2(n_590),
.B(n_578),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_587),
.B(n_495),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_SL g728 ( 
.A1(n_579),
.A2(n_486),
.B(n_645),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_585),
.B(n_534),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_577),
.Y(n_730)
);

AO31x2_ASAP7_75t_L g731 ( 
.A1(n_594),
.A2(n_581),
.A3(n_590),
.B(n_578),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_577),
.Y(n_732)
);

BUFx4f_ASAP7_75t_SL g733 ( 
.A(n_601),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_585),
.B(n_495),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_587),
.B(n_495),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_585),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_624),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_581),
.A2(n_590),
.B(n_578),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_580),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_587),
.B(n_495),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_665),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_688),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_706),
.A2(n_738),
.B(n_726),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_720),
.B(n_725),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_708),
.A2(n_718),
.B1(n_691),
.B2(n_682),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_727),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_660),
.A2(n_684),
.B(n_667),
.Y(n_747)
);

AO21x2_ASAP7_75t_L g748 ( 
.A1(n_726),
.A2(n_738),
.B(n_704),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_739),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_735),
.B(n_740),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_691),
.A2(n_729),
.B1(n_734),
.B2(n_718),
.Y(n_751)
);

INVxp67_ASAP7_75t_SL g752 ( 
.A(n_710),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_684),
.A2(n_664),
.B(n_661),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_662),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_736),
.B(n_681),
.Y(n_755)
);

CKINVDCx6p67_ASAP7_75t_R g756 ( 
.A(n_697),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_717),
.Y(n_757)
);

BUFx2_ASAP7_75t_SL g758 ( 
.A(n_678),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_666),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_716),
.B(n_722),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_685),
.A2(n_701),
.B1(n_687),
.B2(n_698),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_717),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_686),
.B(n_674),
.C(n_672),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_693),
.B(n_723),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_694),
.B(n_692),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_SL g766 ( 
.A(n_703),
.B(n_676),
.C(n_701),
.Y(n_766)
);

OAI21xp5_ASAP7_75t_L g767 ( 
.A1(n_699),
.A2(n_669),
.B(n_728),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_669),
.A2(n_674),
.B(n_670),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_678),
.Y(n_769)
);

CKINVDCx11_ASAP7_75t_R g770 ( 
.A(n_732),
.Y(n_770)
);

AO22x2_ASAP7_75t_L g771 ( 
.A1(n_686),
.A2(n_673),
.B1(n_689),
.B2(n_690),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_690),
.B(n_678),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_724),
.A2(n_737),
.B1(n_695),
.B2(n_679),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_694),
.B(n_709),
.Y(n_774)
);

AO31x2_ASAP7_75t_L g775 ( 
.A1(n_677),
.A2(n_712),
.A3(n_705),
.B(n_714),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_733),
.Y(n_776)
);

BUFx2_ASAP7_75t_R g777 ( 
.A(n_707),
.Y(n_777)
);

OA21x2_ASAP7_75t_L g778 ( 
.A1(n_705),
.A2(n_711),
.B(n_714),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_L g779 ( 
.A(n_732),
.B(n_671),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_719),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_668),
.B(n_712),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_715),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_700),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_730),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_671),
.B(n_668),
.Y(n_785)
);

OR2x6_ASAP7_75t_L g786 ( 
.A(n_702),
.B(n_675),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_713),
.A2(n_731),
.B1(n_663),
.B2(n_696),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_713),
.A2(n_731),
.B(n_663),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_696),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_665),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_739),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_688),
.B(n_683),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_729),
.B(n_534),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_L g794 ( 
.A(n_686),
.B(n_721),
.C(n_680),
.Y(n_794)
);

INVxp67_ASAP7_75t_SL g795 ( 
.A(n_708),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_678),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_665),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_720),
.B(n_725),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_665),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_688),
.B(n_683),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_681),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_SL g802 ( 
.A1(n_745),
.A2(n_795),
.B1(n_744),
.B2(n_798),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_750),
.B(n_745),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_783),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_750),
.B(n_746),
.Y(n_805)
);

AOI21x1_ASAP7_75t_L g806 ( 
.A1(n_788),
.A2(n_743),
.B(n_786),
.Y(n_806)
);

BUFx12f_ASAP7_75t_L g807 ( 
.A(n_770),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_759),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_785),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_748),
.B(n_767),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_772),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_743),
.B(n_741),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_778),
.B(n_747),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_746),
.B(n_793),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_781),
.B(n_751),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_753),
.B(n_789),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_781),
.B(n_794),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_774),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_787),
.B(n_775),
.Y(n_819)
);

AOI21xp33_ASAP7_75t_L g820 ( 
.A1(n_794),
.A2(n_763),
.B(n_771),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_775),
.B(n_771),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_774),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_SL g823 ( 
.A1(n_792),
.A2(n_800),
.B1(n_752),
.B2(n_758),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_775),
.B(n_801),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_761),
.B(n_764),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_760),
.Y(n_826)
);

CKINVDCx14_ASAP7_75t_R g827 ( 
.A(n_776),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_805),
.Y(n_828)
);

NAND3xp33_ASAP7_75t_L g829 ( 
.A(n_802),
.B(n_773),
.C(n_788),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_812),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_812),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_824),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_SL g833 ( 
.A1(n_823),
.A2(n_766),
.B(n_792),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_814),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_806),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_809),
.B(n_797),
.Y(n_836)
);

NAND2x1p5_ASAP7_75t_L g837 ( 
.A(n_818),
.B(n_796),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_825),
.B(n_826),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_825),
.B(n_790),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_808),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_815),
.B(n_803),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_819),
.B(n_799),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_815),
.B(n_803),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_819),
.B(n_768),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_816),
.B(n_813),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_804),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_841),
.B(n_817),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_830),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_840),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_841),
.B(n_843),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_836),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_846),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_836),
.Y(n_853)
);

BUFx12f_ASAP7_75t_L g854 ( 
.A(n_837),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_830),
.Y(n_855)
);

INVx5_ASAP7_75t_L g856 ( 
.A(n_835),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_844),
.B(n_813),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_833),
.B(n_821),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_845),
.B(n_810),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_844),
.B(n_813),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_831),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_828),
.B(n_826),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_850),
.B(n_843),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_857),
.B(n_845),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_857),
.B(n_845),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_849),
.Y(n_866)
);

INVx3_ASAP7_75t_SL g867 ( 
.A(n_851),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_850),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_847),
.B(n_832),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_860),
.B(n_845),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_848),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_853),
.B(n_847),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_852),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_860),
.B(n_852),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_862),
.B(n_842),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_855),
.B(n_832),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_867),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_867),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_864),
.B(n_859),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_868),
.B(n_855),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_864),
.B(n_859),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_871),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_872),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_863),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_876),
.Y(n_885)
);

OAI22xp33_ASAP7_75t_L g886 ( 
.A1(n_874),
.A2(n_858),
.B1(n_854),
.B2(n_833),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_873),
.B(n_859),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_863),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_876),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_885),
.Y(n_890)
);

AOI21xp33_ASAP7_75t_L g891 ( 
.A1(n_878),
.A2(n_866),
.B(n_834),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_885),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_889),
.B(n_869),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_883),
.B(n_869),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_879),
.B(n_865),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_889),
.B(n_875),
.Y(n_896)
);

AOI221x1_ASAP7_75t_L g897 ( 
.A1(n_884),
.A2(n_829),
.B1(n_820),
.B2(n_839),
.C(n_861),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_877),
.A2(n_858),
.B(n_823),
.C(n_827),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_877),
.A2(n_802),
.B1(n_829),
.B2(n_838),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_886),
.A2(n_859),
.B1(n_870),
.B2(n_865),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_882),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_890),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_892),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_894),
.B(n_888),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_891),
.B(n_879),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_893),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_898),
.A2(n_827),
.B(n_754),
.C(n_742),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_906),
.B(n_899),
.Y(n_908)
);

AOI321xp33_ASAP7_75t_L g909 ( 
.A1(n_907),
.A2(n_899),
.A3(n_898),
.B1(n_905),
.B2(n_900),
.C(n_903),
.Y(n_909)
);

OAI221xp5_ASAP7_75t_L g910 ( 
.A1(n_905),
.A2(n_896),
.B1(n_880),
.B2(n_901),
.C(n_882),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_904),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_902),
.A2(n_897),
.B(n_887),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_907),
.B(n_854),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_904),
.Y(n_914)
);

NOR3xp33_ASAP7_75t_L g915 ( 
.A(n_913),
.B(n_791),
.C(n_749),
.Y(n_915)
);

NOR3xp33_ASAP7_75t_L g916 ( 
.A(n_913),
.B(n_796),
.C(n_800),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_914),
.Y(n_917)
);

XNOR2xp5_ASAP7_75t_L g918 ( 
.A(n_908),
.B(n_887),
.Y(n_918)
);

OA22x2_ASAP7_75t_L g919 ( 
.A1(n_909),
.A2(n_887),
.B1(n_895),
.B2(n_881),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_910),
.B(n_756),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_917),
.Y(n_921)
);

OAI21xp33_ASAP7_75t_L g922 ( 
.A1(n_919),
.A2(n_912),
.B(n_911),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_920),
.B(n_807),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_L g924 ( 
.A(n_916),
.B(n_762),
.C(n_757),
.Y(n_924)
);

NOR2x1p5_ASAP7_75t_L g925 ( 
.A(n_915),
.B(n_807),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_SL g926 ( 
.A(n_922),
.B(n_918),
.C(n_807),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_921),
.B(n_901),
.Y(n_927)
);

AND2x2_ASAP7_75t_SL g928 ( 
.A(n_923),
.B(n_769),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_925),
.B(n_856),
.Y(n_929)
);

NOR2x1_ASAP7_75t_L g930 ( 
.A(n_924),
.B(n_780),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_927),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_SL g932 ( 
.A(n_926),
.B(n_928),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_931),
.Y(n_933)
);

OAI222xp33_ASAP7_75t_L g934 ( 
.A1(n_932),
.A2(n_930),
.B1(n_929),
.B2(n_837),
.C1(n_822),
.C2(n_765),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_933),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_933),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_935),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_937),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_937),
.A2(n_936),
.B1(n_934),
.B2(n_777),
.Y(n_939)
);

OAI221xp5_ASAP7_75t_L g940 ( 
.A1(n_938),
.A2(n_784),
.B1(n_814),
.B2(n_755),
.C(n_765),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_940),
.A2(n_939),
.B1(n_777),
.B2(n_837),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_941),
.B(n_811),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_942),
.A2(n_782),
.B(n_779),
.Y(n_943)
);


endmodule