module fake_jpeg_13487_n_37 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_37);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

OA22x2_ASAP7_75t_SL g17 ( 
.A1(n_15),
.A2(n_5),
.B1(n_7),
.B2(n_6),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_18),
.B(n_20),
.Y(n_21)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_16),
.B(n_0),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_14),
.C(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_23),
.B(n_24),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_4),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_2),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_3),
.Y(n_33)
);

FAx1_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_34),
.CI(n_26),
.CON(n_35),
.SN(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_32),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_35),
.B(n_12),
.Y(n_37)
);


endmodule