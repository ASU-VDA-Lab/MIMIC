module fake_aes_1889_n_1305 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1305);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1305;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1130;
wire n_584;
wire n_1042;
wire n_912;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1219;
wire n_1120;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g277 ( .A(n_60), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_118), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_187), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_163), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_30), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_164), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_208), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_223), .Y(n_284) );
INVxp33_ASAP7_75t_L g285 ( .A(n_213), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_62), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_24), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_11), .Y(n_288) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_126), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_9), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_205), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_190), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_176), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_61), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_0), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_177), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_133), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_91), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_75), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_3), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_171), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_197), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_193), .Y(n_303) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_215), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_247), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_86), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_84), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_8), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_214), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_263), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_220), .Y(n_311) );
INVxp33_ASAP7_75t_SL g312 ( .A(n_230), .Y(n_312) );
NOR2xp67_ASAP7_75t_L g313 ( .A(n_199), .B(n_61), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_259), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_4), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_200), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_112), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_142), .Y(n_318) );
INVxp33_ASAP7_75t_SL g319 ( .A(n_262), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_3), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_226), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_210), .Y(n_322) );
INVxp33_ASAP7_75t_L g323 ( .A(n_153), .Y(n_323) );
INVx4_ASAP7_75t_R g324 ( .A(n_149), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_179), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_160), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_76), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_231), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_232), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_261), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_140), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_182), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_266), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_34), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_68), .Y(n_335) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_79), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_93), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_155), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_198), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_98), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_138), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_85), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_203), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_162), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_172), .Y(n_345) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_70), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_83), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_136), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_116), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_229), .Y(n_350) );
BUFx10_ASAP7_75t_L g351 ( .A(n_170), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_265), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_151), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_13), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_183), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_25), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_242), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_216), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_204), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_28), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_159), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_189), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_71), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_107), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_49), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_224), .Y(n_366) );
INVxp67_ASAP7_75t_L g367 ( .A(n_194), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_254), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_120), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_123), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_16), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_212), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_175), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_89), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_110), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_73), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_34), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_28), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_77), .Y(n_379) );
INVxp33_ASAP7_75t_SL g380 ( .A(n_66), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_54), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_240), .Y(n_382) );
INVxp33_ASAP7_75t_L g383 ( .A(n_245), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_67), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_150), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_63), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_22), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_228), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_17), .B(n_239), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_62), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_41), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_100), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_211), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_249), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_38), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_244), .Y(n_396) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_92), .Y(n_397) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_173), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_206), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_269), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_8), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_49), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_47), .Y(n_403) );
CKINVDCx14_ASAP7_75t_R g404 ( .A(n_246), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_264), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_90), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_152), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_235), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_174), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_146), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_65), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_185), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_297), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_337), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_297), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_281), .Y(n_416) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_340), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_337), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_381), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_297), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_351), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_402), .B(n_0), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_286), .B(n_1), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_281), .Y(n_424) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_337), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_334), .Y(n_426) );
OAI22xp5_ASAP7_75t_SL g427 ( .A1(n_295), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_351), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_340), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_359), .B(n_2), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_295), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_396), .B(n_5), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_285), .B(n_6), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_351), .B(n_7), .Y(n_434) );
INVx3_ASAP7_75t_L g435 ( .A(n_402), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_334), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_278), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_337), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_350), .Y(n_439) );
AND2x6_ASAP7_75t_L g440 ( .A(n_280), .B(n_64), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_308), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_282), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_346), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_283), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_395), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_413), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_421), .B(n_285), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_437), .B(n_323), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_413), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_445), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_422), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_421), .B(n_323), .Y(n_453) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_431), .A2(n_403), .B1(n_388), .B2(n_392), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_445), .B(n_383), .Y(n_455) );
BUFx4f_ASAP7_75t_L g456 ( .A(n_440), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_433), .A2(n_287), .B1(n_288), .B2(n_277), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_413), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_415), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_414), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_421), .B(n_383), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_421), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_417), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_415), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_414), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_415), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_428), .B(n_279), .Y(n_467) );
AO22x2_ASAP7_75t_L g468 ( .A1(n_422), .A2(n_389), .B1(n_284), .B2(n_344), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_419), .B(n_290), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_419), .B(n_404), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_433), .B(n_404), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_437), .B(n_333), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_418), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_428), .B(n_279), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_418), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_428), .B(n_367), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_428), .B(n_298), .Y(n_477) );
BUFx4f_ASAP7_75t_L g478 ( .A(n_440), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_422), .B(n_294), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_440), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_442), .B(n_298), .Y(n_481) );
OAI22xp5_ASAP7_75t_SL g482 ( .A1(n_429), .A2(n_388), .B1(n_392), .B2(n_350), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_433), .B(n_307), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_422), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_439), .Y(n_485) );
AND2x6_ASAP7_75t_L g486 ( .A(n_420), .B(n_280), .Y(n_486) );
AO22x2_ASAP7_75t_L g487 ( .A1(n_420), .A2(n_344), .B1(n_355), .B2(n_333), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_448), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_462), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_457), .A2(n_431), .B1(n_432), .B2(n_443), .Y(n_490) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_480), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_448), .B(n_442), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_468), .A2(n_444), .B1(n_440), .B2(n_435), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_462), .Y(n_494) );
NAND2x1p5_ASAP7_75t_L g495 ( .A(n_471), .B(n_434), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_471), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_483), .B(n_432), .Y(n_497) );
HB1xp67_ASAP7_75t_SL g498 ( .A(n_463), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_447), .B(n_444), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_482), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_446), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_450), .B(n_423), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_483), .B(n_430), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_455), .B(n_435), .Y(n_504) );
NOR2x2_ASAP7_75t_L g505 ( .A(n_482), .B(n_427), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_451), .Y(n_506) );
AND2x6_ASAP7_75t_SL g507 ( .A(n_485), .B(n_300), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_446), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_468), .A2(n_440), .B1(n_435), .B2(n_424), .Y(n_509) );
INVx1_ASAP7_75t_SL g510 ( .A(n_450), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_449), .Y(n_511) );
OAI21xp33_ASAP7_75t_SL g512 ( .A1(n_451), .A2(n_424), .B(n_416), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_470), .A2(n_312), .B1(n_380), .B2(n_319), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_449), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_470), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_468), .A2(n_440), .B1(n_426), .B2(n_436), .Y(n_516) );
BUFx6f_ASAP7_75t_SL g517 ( .A(n_479), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_468), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_458), .Y(n_519) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_480), .Y(n_520) );
AND2x6_ASAP7_75t_SL g521 ( .A(n_455), .B(n_315), .Y(n_521) );
INVxp67_ASAP7_75t_L g522 ( .A(n_469), .Y(n_522) );
NOR2x1_ASAP7_75t_R g523 ( .A(n_453), .B(n_307), .Y(n_523) );
AND2x4_ASAP7_75t_SL g524 ( .A(n_479), .B(n_451), .Y(n_524) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_484), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_458), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_456), .B(n_314), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_469), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_459), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_477), .B(n_314), .Y(n_530) );
INVxp67_ASAP7_75t_SL g531 ( .A(n_484), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_459), .Y(n_532) );
AO22x1_ASAP7_75t_L g533 ( .A1(n_479), .A2(n_319), .B1(n_380), .B2(n_312), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_464), .Y(n_534) );
BUFx4f_ASAP7_75t_L g535 ( .A(n_479), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_464), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_481), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_476), .B(n_322), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_461), .B(n_322), .Y(n_539) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_480), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_456), .B(n_331), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_467), .B(n_416), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_478), .B(n_331), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_474), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_466), .Y(n_545) );
NAND3xp33_ASAP7_75t_SL g546 ( .A(n_472), .B(n_341), .C(n_332), .Y(n_546) );
NOR2xp67_ASAP7_75t_L g547 ( .A(n_472), .B(n_426), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_484), .B(n_332), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_478), .B(n_341), .Y(n_549) );
INVx3_ASAP7_75t_L g550 ( .A(n_484), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_466), .B(n_374), .Y(n_551) );
BUFx12f_ASAP7_75t_SL g552 ( .A(n_454), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_487), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_478), .B(n_375), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_487), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_487), .A2(n_440), .B1(n_436), .B2(n_320), .Y(n_556) );
CKINVDCx8_ASAP7_75t_R g557 ( .A(n_486), .Y(n_557) );
INVx3_ASAP7_75t_L g558 ( .A(n_486), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_486), .B(n_393), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_478), .B(n_393), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_486), .B(n_409), .Y(n_561) );
INVxp67_ASAP7_75t_SL g562 ( .A(n_486), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_486), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_486), .A2(n_440), .B1(n_354), .B2(n_360), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_465), .B(n_409), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_452), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_465), .B(n_411), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_452), .B(n_411), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_452), .A2(n_365), .B1(n_371), .B2(n_356), .Y(n_569) );
CKINVDCx11_ASAP7_75t_R g570 ( .A(n_465), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_460), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_460), .A2(n_440), .B1(n_377), .B2(n_386), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_488), .B(n_378), .Y(n_573) );
OAI22xp5_ASAP7_75t_SL g574 ( .A1(n_500), .A2(n_391), .B1(n_401), .B2(n_387), .Y(n_574) );
BUFx2_ASAP7_75t_L g575 ( .A(n_510), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_518), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_506), .Y(n_577) );
INVx4_ASAP7_75t_L g578 ( .A(n_517), .Y(n_578) );
BUFx2_ASAP7_75t_L g579 ( .A(n_528), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_525), .A2(n_304), .B(n_289), .Y(n_580) );
OR2x6_ASAP7_75t_L g581 ( .A(n_522), .B(n_313), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_547), .Y(n_582) );
A2O1A1Ixp33_ASAP7_75t_L g583 ( .A1(n_512), .A2(n_292), .B(n_296), .C(n_291), .Y(n_583) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_570), .Y(n_584) );
INVx3_ASAP7_75t_L g585 ( .A(n_518), .Y(n_585) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_491), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_497), .B(n_336), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_502), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_506), .Y(n_589) );
BUFx12f_ASAP7_75t_L g590 ( .A(n_507), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_550), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_535), .Y(n_592) );
CKINVDCx12_ASAP7_75t_R g593 ( .A(n_523), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_550), .Y(n_594) );
BUFx2_ASAP7_75t_L g595 ( .A(n_522), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_525), .A2(n_398), .B(n_397), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_497), .B(n_382), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_496), .Y(n_598) );
INVx2_ASAP7_75t_SL g599 ( .A(n_535), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_498), .Y(n_600) );
BUFx3_ASAP7_75t_L g601 ( .A(n_544), .Y(n_601) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_491), .Y(n_602) );
BUFx3_ASAP7_75t_L g603 ( .A(n_542), .Y(n_603) );
INVx3_ASAP7_75t_L g604 ( .A(n_524), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_542), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_531), .A2(n_301), .B(n_299), .Y(n_606) );
NOR2x1_ASAP7_75t_R g607 ( .A(n_515), .B(n_293), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_531), .A2(n_492), .B(n_503), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_548), .A2(n_303), .B(n_302), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_508), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_501), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_519), .Y(n_612) );
CKINVDCx11_ASAP7_75t_R g613 ( .A(n_521), .Y(n_613) );
INVxp67_ASAP7_75t_SL g614 ( .A(n_516), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_517), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_526), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_553), .A2(n_390), .B1(n_308), .B2(n_305), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_532), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_504), .Y(n_619) );
CKINVDCx11_ASAP7_75t_R g620 ( .A(n_498), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_490), .A2(n_306), .B(n_310), .C(n_309), .Y(n_621) );
INVx5_ASAP7_75t_L g622 ( .A(n_558), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_491), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_534), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_511), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_513), .B(n_311), .Y(n_626) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_491), .Y(n_627) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_520), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_555), .A2(n_316), .B(n_318), .C(n_317), .Y(n_629) );
BUFx2_ASAP7_75t_L g630 ( .A(n_552), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_514), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_533), .B(n_308), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_529), .Y(n_633) );
OR2x2_ASAP7_75t_SL g634 ( .A(n_505), .B(n_308), .Y(n_634) );
INVx3_ASAP7_75t_L g635 ( .A(n_557), .Y(n_635) );
OR2x6_ASAP7_75t_SL g636 ( .A(n_537), .B(n_324), .Y(n_636) );
OAI22x1_ASAP7_75t_L g637 ( .A1(n_495), .A2(n_325), .B1(n_326), .B2(n_321), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_536), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_545), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_495), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_562), .B(n_327), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_489), .Y(n_642) );
AO32x2_ASAP7_75t_L g643 ( .A1(n_516), .A2(n_425), .A3(n_418), .B1(n_347), .B2(n_353), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_493), .B(n_328), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_499), .B(n_390), .Y(n_645) );
INVx5_ASAP7_75t_L g646 ( .A(n_558), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_530), .A2(n_330), .B(n_329), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_527), .A2(n_339), .B(n_338), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_569), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_546), .A2(n_343), .B1(n_345), .B2(n_342), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_551), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_538), .A2(n_390), .B1(n_335), .B2(n_349), .Y(n_652) );
AO21x1_ASAP7_75t_L g653 ( .A1(n_562), .A2(n_352), .B(n_348), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_493), .B(n_357), .Y(n_654) );
BUFx10_ASAP7_75t_L g655 ( .A(n_554), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_494), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_559), .Y(n_657) );
AND2x4_ASAP7_75t_L g658 ( .A(n_539), .B(n_358), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_541), .A2(n_362), .B(n_361), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_563), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_546), .B(n_363), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_520), .Y(n_662) );
BUFx3_ASAP7_75t_L g663 ( .A(n_561), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_509), .B(n_364), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g665 ( .A1(n_509), .A2(n_368), .B(n_369), .C(n_366), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_556), .B(n_10), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_543), .A2(n_372), .B(n_370), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_556), .B(n_373), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_520), .Y(n_669) );
INVx3_ASAP7_75t_SL g670 ( .A(n_565), .Y(n_670) );
NAND2x1_ASAP7_75t_L g671 ( .A(n_564), .B(n_405), .Y(n_671) );
BUFx2_ASAP7_75t_L g672 ( .A(n_540), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_567), .Y(n_673) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_540), .Y(n_674) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_540), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_549), .A2(n_379), .B(n_376), .Y(n_676) );
BUFx2_ASAP7_75t_L g677 ( .A(n_540), .Y(n_677) );
INVx3_ASAP7_75t_L g678 ( .A(n_571), .Y(n_678) );
BUFx12f_ASAP7_75t_L g679 ( .A(n_564), .Y(n_679) );
INVx2_ASAP7_75t_SL g680 ( .A(n_568), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_560), .B(n_384), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_572), .B(n_385), .Y(n_682) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_566), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_566), .Y(n_684) );
INVx1_ASAP7_75t_SL g685 ( .A(n_572), .Y(n_685) );
AO32x1_ASAP7_75t_L g686 ( .A1(n_518), .A2(n_438), .A3(n_394), .B1(n_399), .B2(n_408), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g687 ( .A1(n_512), .A2(n_412), .B(n_407), .C(n_410), .Y(n_687) );
INVx3_ASAP7_75t_L g688 ( .A(n_518), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_510), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_522), .A2(n_406), .B(n_441), .C(n_335), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_506), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_506), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_506), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_518), .A2(n_406), .B1(n_349), .B2(n_441), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_506), .Y(n_695) );
AND2x4_ASAP7_75t_L g696 ( .A(n_488), .B(n_10), .Y(n_696) );
BUFx2_ASAP7_75t_L g697 ( .A(n_510), .Y(n_697) );
INVx3_ASAP7_75t_L g698 ( .A(n_576), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_575), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_597), .A2(n_353), .B(n_347), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_611), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_611), .Y(n_702) );
BUFx12f_ASAP7_75t_L g703 ( .A(n_620), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_696), .B(n_347), .Y(n_704) );
BUFx3_ASAP7_75t_L g705 ( .A(n_584), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_598), .Y(n_706) );
OR2x2_ASAP7_75t_L g707 ( .A(n_697), .B(n_11), .Y(n_707) );
BUFx12f_ASAP7_75t_L g708 ( .A(n_584), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_588), .A2(n_441), .B1(n_400), .B2(n_353), .C(n_425), .Y(n_709) );
INVx1_ASAP7_75t_SL g710 ( .A(n_689), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_649), .B(n_12), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_595), .B(n_12), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_639), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_608), .A2(n_475), .B(n_473), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_679), .A2(n_400), .B1(n_353), .B2(n_425), .Y(n_715) );
BUFx6f_ASAP7_75t_L g716 ( .A(n_586), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_579), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_626), .A2(n_425), .B1(n_465), .B2(n_15), .C(n_16), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_696), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_719) );
NOR2xp67_ASAP7_75t_SL g720 ( .A(n_584), .B(n_14), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_612), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_634), .Y(n_722) );
INVx1_ASAP7_75t_SL g723 ( .A(n_601), .Y(n_723) );
AO31x2_ASAP7_75t_L g724 ( .A1(n_653), .A2(n_17), .A3(n_18), .B(n_19), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_612), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_616), .Y(n_726) );
AO21x2_ASAP7_75t_L g727 ( .A1(n_583), .A2(n_465), .B(n_72), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_616), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_618), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_619), .B(n_18), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g731 ( .A1(n_621), .A2(n_465), .B(n_20), .C(n_21), .Y(n_731) );
BUFx12f_ASAP7_75t_L g732 ( .A(n_613), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_618), .Y(n_733) );
OAI21x1_ASAP7_75t_L g734 ( .A1(n_660), .A2(n_74), .B(n_69), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_624), .Y(n_735) );
BUFx8_ASAP7_75t_SL g736 ( .A(n_590), .Y(n_736) );
OA21x2_ASAP7_75t_L g737 ( .A1(n_687), .A2(n_80), .B(n_78), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_624), .Y(n_738) );
OAI21x1_ASAP7_75t_SL g739 ( .A1(n_638), .A2(n_19), .B(n_20), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_638), .Y(n_740) );
OAI21x1_ASAP7_75t_L g741 ( .A1(n_660), .A2(n_82), .B(n_81), .Y(n_741) );
AND2x4_ASAP7_75t_L g742 ( .A(n_578), .B(n_21), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_683), .Y(n_743) );
INVxp67_ASAP7_75t_L g744 ( .A(n_607), .Y(n_744) );
BUFx2_ASAP7_75t_L g745 ( .A(n_578), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_573), .Y(n_746) );
NOR2xp67_ASAP7_75t_L g747 ( .A(n_600), .B(n_22), .Y(n_747) );
O2A1O1Ixp33_ASAP7_75t_L g748 ( .A1(n_661), .A2(n_23), .B(n_24), .C(n_25), .Y(n_748) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_576), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_614), .A2(n_23), .B1(n_26), .B2(n_27), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_651), .A2(n_88), .B(n_87), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_668), .A2(n_27), .B1(n_29), .B2(n_30), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_586), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_658), .B(n_29), .Y(n_754) );
BUFx3_ASAP7_75t_L g755 ( .A(n_672), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_630), .B(n_31), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_658), .B(n_31), .Y(n_757) );
BUFx12f_ASAP7_75t_L g758 ( .A(n_640), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_668), .A2(n_32), .B1(n_33), .B2(n_35), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_609), .A2(n_95), .B(n_94), .Y(n_760) );
OAI21x1_ASAP7_75t_L g761 ( .A1(n_662), .A2(n_97), .B(n_96), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_647), .A2(n_101), .B(n_99), .Y(n_762) );
OA21x2_ASAP7_75t_L g763 ( .A1(n_665), .A2(n_154), .B(n_275), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_656), .Y(n_764) );
OAI21x1_ASAP7_75t_L g765 ( .A1(n_669), .A2(n_148), .B(n_274), .Y(n_765) );
OAI21x1_ASAP7_75t_L g766 ( .A1(n_678), .A2(n_147), .B(n_273), .Y(n_766) );
OAI21x1_ASAP7_75t_L g767 ( .A1(n_678), .A2(n_145), .B(n_272), .Y(n_767) );
AO21x2_ASAP7_75t_L g768 ( .A1(n_632), .A2(n_144), .B(n_271), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_586), .Y(n_769) );
INVxp67_ASAP7_75t_SL g770 ( .A(n_585), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_603), .B(n_32), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_605), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_645), .A2(n_143), .B(n_270), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_666), .A2(n_33), .B1(n_35), .B2(n_36), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_587), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_602), .B(n_102), .Y(n_776) );
OAI21x1_ASAP7_75t_L g777 ( .A1(n_671), .A2(n_158), .B(n_268), .Y(n_777) );
AO21x2_ASAP7_75t_L g778 ( .A1(n_644), .A2(n_157), .B(n_267), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_685), .A2(n_37), .B1(n_39), .B2(n_40), .Y(n_779) );
BUFx3_ASAP7_75t_L g780 ( .A(n_677), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_592), .B(n_39), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_574), .A2(n_40), .B1(n_41), .B2(n_42), .Y(n_782) );
OAI21x1_ASAP7_75t_L g783 ( .A1(n_694), .A2(n_161), .B(n_260), .Y(n_783) );
OAI222xp33_ASAP7_75t_L g784 ( .A1(n_581), .A2(n_42), .B1(n_43), .B2(n_44), .C1(n_45), .C2(n_46), .Y(n_784) );
AO21x2_ASAP7_75t_L g785 ( .A1(n_654), .A2(n_156), .B(n_258), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_642), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_604), .B(n_43), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g788 ( .A1(n_606), .A2(n_165), .B(n_257), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_593), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_650), .B(n_44), .Y(n_790) );
OA21x2_ASAP7_75t_L g791 ( .A1(n_664), .A2(n_141), .B(n_256), .Y(n_791) );
OAI21x1_ASAP7_75t_L g792 ( .A1(n_690), .A2(n_139), .B(n_255), .Y(n_792) );
NAND2x1p5_ASAP7_75t_L g793 ( .A(n_585), .B(n_688), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_673), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_610), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_625), .Y(n_796) );
NAND2xp5_ASAP7_75t_SL g797 ( .A(n_602), .B(n_103), .Y(n_797) );
OAI21x1_ASAP7_75t_L g798 ( .A1(n_648), .A2(n_166), .B(n_253), .Y(n_798) );
AO21x2_ASAP7_75t_L g799 ( .A1(n_682), .A2(n_137), .B(n_252), .Y(n_799) );
OAI21x1_ASAP7_75t_L g800 ( .A1(n_659), .A2(n_135), .B(n_251), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_688), .A2(n_45), .B1(n_46), .B2(n_47), .Y(n_801) );
BUFx2_ASAP7_75t_R g802 ( .A(n_636), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_631), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_641), .A2(n_48), .B1(n_50), .B2(n_51), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_604), .B(n_50), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_580), .A2(n_168), .B(n_250), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_599), .B(n_51), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_633), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_581), .B(n_52), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_637), .B(n_53), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_582), .B(n_53), .Y(n_811) );
OAI21x1_ASAP7_75t_L g812 ( .A1(n_667), .A2(n_178), .B(n_248), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_680), .B(n_54), .Y(n_813) );
OA21x2_ASAP7_75t_L g814 ( .A1(n_617), .A2(n_169), .B(n_243), .Y(n_814) );
OAI21x1_ASAP7_75t_L g815 ( .A1(n_676), .A2(n_167), .B(n_241), .Y(n_815) );
INVx8_ASAP7_75t_L g816 ( .A(n_615), .Y(n_816) );
BUFx2_ASAP7_75t_SL g817 ( .A(n_615), .Y(n_817) );
OAI22xp33_ASAP7_75t_L g818 ( .A1(n_681), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_818) );
OA21x2_ASAP7_75t_L g819 ( .A1(n_686), .A2(n_134), .B(n_238), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_684), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_602), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_623), .Y(n_822) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_655), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_823) );
OA21x2_ASAP7_75t_L g824 ( .A1(n_686), .A2(n_181), .B(n_237), .Y(n_824) );
OR2x2_ASAP7_75t_L g825 ( .A(n_670), .B(n_58), .Y(n_825) );
OAI21x1_ASAP7_75t_L g826 ( .A1(n_629), .A2(n_180), .B(n_236), .Y(n_826) );
INVxp67_ASAP7_75t_L g827 ( .A(n_641), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_657), .B(n_58), .Y(n_828) );
OAI21x1_ASAP7_75t_L g829 ( .A1(n_577), .A2(n_132), .B(n_234), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_623), .Y(n_830) );
AO21x2_ASAP7_75t_L g831 ( .A1(n_686), .A2(n_131), .B(n_233), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_577), .B(n_59), .Y(n_832) );
AOI221xp5_ASAP7_75t_L g833 ( .A1(n_746), .A2(n_596), .B1(n_652), .B2(n_591), .C(n_693), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_722), .A2(n_655), .B1(n_663), .B2(n_591), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_719), .A2(n_675), .B1(n_623), .B2(n_628), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_719), .A2(n_675), .B1(n_627), .B2(n_628), .Y(n_836) );
OAI21xp5_ASAP7_75t_L g837 ( .A1(n_731), .A2(n_693), .B(n_594), .Y(n_837) );
AOI21xp33_ASAP7_75t_R g838 ( .A1(n_747), .A2(n_635), .B(n_643), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_711), .A2(n_695), .B1(n_692), .B2(n_691), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_710), .B(n_589), .Y(n_840) );
NAND3xp33_ASAP7_75t_SL g841 ( .A(n_794), .B(n_643), .C(n_60), .Y(n_841) );
AOI221xp5_ASAP7_75t_L g842 ( .A1(n_711), .A2(n_635), .B1(n_622), .B2(n_646), .C(n_674), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_701), .B(n_646), .Y(n_843) );
AOI221xp5_ASAP7_75t_L g844 ( .A1(n_712), .A2(n_646), .B1(n_622), .B2(n_628), .C(n_627), .Y(n_844) );
AOI222xp33_ASAP7_75t_L g845 ( .A1(n_809), .A2(n_706), .B1(n_712), .B2(n_713), .C1(n_784), .C2(n_756), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_764), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_702), .A2(n_674), .B1(n_643), .B2(n_622), .Y(n_847) );
INVx3_ASAP7_75t_L g848 ( .A(n_793), .Y(n_848) );
OAI211xp5_ASAP7_75t_L g849 ( .A1(n_782), .A2(n_59), .B(n_63), .C(n_104), .Y(n_849) );
AOI21xp33_ASAP7_75t_L g850 ( .A1(n_704), .A2(n_105), .B(n_106), .Y(n_850) );
BUFx3_ASAP7_75t_L g851 ( .A(n_708), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_702), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_794), .A2(n_108), .B1(n_109), .B2(n_111), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_726), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_743), .B(n_117), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_743), .B(n_119), .Y(n_856) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_699), .A2(n_774), .B1(n_818), .B2(n_820), .C(n_828), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_726), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_786), .Y(n_859) );
OAI221xp5_ASAP7_75t_L g860 ( .A1(n_699), .A2(n_121), .B1(n_122), .B2(n_124), .C(n_125), .Y(n_860) );
BUFx2_ASAP7_75t_L g861 ( .A(n_717), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_707), .B(n_127), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g863 ( .A1(n_714), .A2(n_128), .B(n_129), .Y(n_863) );
AOI222xp33_ASAP7_75t_L g864 ( .A1(n_744), .A2(n_130), .B1(n_184), .B2(n_186), .C1(n_188), .C2(n_191), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_721), .Y(n_865) );
INVx4_ASAP7_75t_L g866 ( .A(n_708), .Y(n_866) );
AOI221xp5_ASAP7_75t_SL g867 ( .A1(n_731), .A2(n_192), .B1(n_195), .B2(n_196), .C(n_201), .Y(n_867) );
AOI21xp5_ASAP7_75t_L g868 ( .A1(n_704), .A2(n_202), .B(n_207), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_725), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_729), .Y(n_870) );
OR2x6_ASAP7_75t_L g871 ( .A(n_703), .B(n_209), .Y(n_871) );
OAI21xp5_ASAP7_75t_L g872 ( .A1(n_832), .A2(n_217), .B(n_218), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_728), .Y(n_873) );
A2O1A1Ixp33_ASAP7_75t_SL g874 ( .A1(n_720), .A2(n_219), .B(n_221), .C(n_222), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_735), .Y(n_875) );
CKINVDCx5p33_ASAP7_75t_R g876 ( .A(n_736), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_828), .A2(n_225), .B1(n_227), .B2(n_276), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_723), .B(n_827), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_728), .B(n_733), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_790), .A2(n_781), .B1(n_832), .B2(n_754), .Y(n_880) );
AND2x4_ASAP7_75t_SL g881 ( .A(n_742), .B(n_733), .Y(n_881) );
AOI222xp33_ASAP7_75t_L g882 ( .A1(n_703), .A2(n_740), .B1(n_742), .B2(n_732), .C1(n_752), .C2(n_759), .Y(n_882) );
NAND2x1_ASAP7_75t_L g883 ( .A(n_738), .B(n_698), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_781), .A2(n_757), .B1(n_771), .B2(n_742), .Y(n_884) );
OAI221xp5_ASAP7_75t_L g885 ( .A1(n_775), .A2(n_752), .B1(n_759), .B2(n_804), .C(n_810), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_730), .A2(n_738), .B1(n_813), .B2(n_787), .Y(n_886) );
AO31x2_ASAP7_75t_L g887 ( .A1(n_750), .A2(n_753), .A3(n_830), .B(n_769), .Y(n_887) );
OAI21xp5_ASAP7_75t_L g888 ( .A1(n_792), .A2(n_826), .B(n_783), .Y(n_888) );
AOI222xp33_ASAP7_75t_L g889 ( .A1(n_732), .A2(n_818), .B1(n_804), .B2(n_775), .C1(n_789), .C2(n_772), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_805), .A2(n_823), .B1(n_807), .B2(n_780), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_755), .A2(n_780), .B1(n_811), .B2(n_705), .Y(n_891) );
OA21x2_ASAP7_75t_L g892 ( .A1(n_777), .A2(n_792), .B(n_826), .Y(n_892) );
OAI21xp5_ASAP7_75t_L g893 ( .A1(n_783), .A2(n_806), .B(n_762), .Y(n_893) );
AND2x4_ASAP7_75t_L g894 ( .A(n_705), .B(n_770), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_825), .B(n_795), .Y(n_895) );
NAND2xp33_ASAP7_75t_R g896 ( .A(n_789), .B(n_745), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_796), .B(n_808), .Y(n_897) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_758), .B(n_817), .Y(n_898) );
OAI221xp5_ASAP7_75t_L g899 ( .A1(n_718), .A2(n_748), .B1(n_715), .B2(n_700), .C(n_779), .Y(n_899) );
OR2x6_ASAP7_75t_L g900 ( .A(n_816), .B(n_758), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_803), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_739), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_801), .A2(n_770), .B1(n_816), .B2(n_737), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_755), .A2(n_749), .B1(n_816), .B2(n_698), .Y(n_904) );
OR2x2_ASAP7_75t_L g905 ( .A(n_724), .B(n_749), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_724), .Y(n_906) );
OAI22xp33_ASAP7_75t_L g907 ( .A1(n_793), .A2(n_802), .B1(n_788), .B2(n_737), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_715), .A2(n_709), .B1(n_737), .B2(n_727), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_814), .A2(n_791), .B1(n_763), .B2(n_716), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_724), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_753), .Y(n_911) );
A2O1A1Ixp33_ASAP7_75t_L g912 ( .A1(n_760), .A2(n_751), .B(n_773), .C(n_800), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_724), .Y(n_913) );
INVx3_ASAP7_75t_L g914 ( .A(n_716), .Y(n_914) );
OAI21xp5_ASAP7_75t_L g915 ( .A1(n_798), .A2(n_815), .B(n_812), .Y(n_915) );
BUFx3_ASAP7_75t_L g916 ( .A(n_736), .Y(n_916) );
HB1xp67_ASAP7_75t_L g917 ( .A(n_769), .Y(n_917) );
INVx3_ASAP7_75t_L g918 ( .A(n_716), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_829), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_766), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_727), .A2(n_814), .B1(n_830), .B2(n_822), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_821), .A2(n_822), .B1(n_785), .B2(n_778), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_821), .B(n_831), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_776), .A2(n_797), .B1(n_785), .B2(n_778), .C(n_799), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_716), .B(n_799), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_831), .A2(n_768), .B1(n_819), .B2(n_824), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_768), .A2(n_824), .B1(n_819), .B2(n_767), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_824), .A2(n_734), .B1(n_741), .B2(n_761), .Y(n_928) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_765), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_722), .A2(n_552), .B1(n_482), .B2(n_630), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_743), .B(n_588), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_722), .A2(n_552), .B1(n_482), .B2(n_630), .Y(n_932) );
AND2x2_ASAP7_75t_L g933 ( .A(n_743), .B(n_588), .Y(n_933) );
AOI332xp33_ASAP7_75t_L g934 ( .A1(n_782), .A2(n_431), .A3(n_505), .B1(n_457), .B2(n_598), .B3(n_290), .C1(n_294), .C2(n_287), .Y(n_934) );
AOI22xp33_ASAP7_75t_SL g935 ( .A1(n_722), .A2(n_417), .B1(n_439), .B2(n_429), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_722), .A2(n_552), .B1(n_482), .B2(n_630), .Y(n_936) );
OAI211xp5_ASAP7_75t_L g937 ( .A1(n_782), .A2(n_722), .B(n_823), .C(n_711), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_701), .Y(n_938) );
AOI221xp5_ASAP7_75t_L g939 ( .A1(n_746), .A2(n_454), .B1(n_522), .B2(n_490), .C(n_528), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_713), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g941 ( .A1(n_746), .A2(n_454), .B1(n_522), .B2(n_490), .C(n_528), .Y(n_941) );
INVxp67_ASAP7_75t_L g942 ( .A(n_699), .Y(n_942) );
A2O1A1Ixp33_ASAP7_75t_L g943 ( .A1(n_711), .A2(n_746), .B(n_629), .C(n_608), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_722), .A2(n_552), .B1(n_482), .B2(n_630), .Y(n_944) );
OAI22xp33_ASAP7_75t_L g945 ( .A1(n_722), .A2(n_429), .B1(n_439), .B2(n_417), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_722), .A2(n_552), .B1(n_482), .B2(n_630), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g947 ( .A1(n_746), .A2(n_454), .B1(n_522), .B2(n_490), .C(n_528), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_719), .A2(n_518), .B1(n_696), .B2(n_701), .Y(n_948) );
AOI22xp33_ASAP7_75t_SL g949 ( .A1(n_722), .A2(n_417), .B1(n_439), .B2(n_429), .Y(n_949) );
OAI22xp5_ASAP7_75t_SL g950 ( .A1(n_794), .A2(n_634), .B1(n_482), .B2(n_429), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_743), .B(n_588), .Y(n_951) );
BUFx2_ASAP7_75t_L g952 ( .A(n_894), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_879), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_879), .Y(n_954) );
INVxp67_ASAP7_75t_R g955 ( .A(n_950), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_852), .B(n_858), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_873), .B(n_938), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_906), .B(n_910), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_913), .Y(n_959) );
BUFx2_ASAP7_75t_L g960 ( .A(n_894), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_865), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_897), .B(n_881), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_869), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_889), .A2(n_882), .B1(n_845), .B2(n_948), .Y(n_964) );
BUFx3_ASAP7_75t_L g965 ( .A(n_900), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_870), .Y(n_966) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_835), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_875), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_943), .B(n_940), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_905), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_846), .B(n_859), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_901), .B(n_931), .Y(n_972) );
OR2x2_ASAP7_75t_L g973 ( .A(n_948), .B(n_933), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_951), .B(n_895), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_902), .B(n_835), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_880), .B(n_857), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_855), .B(n_856), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_923), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_911), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_917), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_920), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_848), .B(n_843), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_847), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_848), .B(n_843), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_847), .Y(n_985) );
OAI22xp33_ASAP7_75t_L g986 ( .A1(n_885), .A2(n_871), .B1(n_836), .B2(n_872), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_884), .B(n_862), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_919), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_836), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_839), .B(n_886), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_883), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_942), .B(n_837), .Y(n_992) );
AND2x4_ASAP7_75t_L g993 ( .A(n_914), .B(n_918), .Y(n_993) );
BUFx3_ASAP7_75t_L g994 ( .A(n_900), .Y(n_994) );
INVx2_ASAP7_75t_L g995 ( .A(n_892), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_837), .B(n_903), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_872), .B(n_861), .Y(n_997) );
NAND2xp5_ASAP7_75t_SL g998 ( .A(n_907), .B(n_864), .Y(n_998) );
INVx4_ASAP7_75t_R g999 ( .A(n_851), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_885), .B(n_833), .Y(n_1000) );
INVx5_ASAP7_75t_L g1001 ( .A(n_900), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_925), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_891), .B(n_941), .Y(n_1003) );
BUFx2_ASAP7_75t_SL g1004 ( .A(n_866), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_939), .B(n_947), .Y(n_1005) );
INVx3_ASAP7_75t_L g1006 ( .A(n_914), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_925), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_929), .Y(n_1008) );
INVx2_ASAP7_75t_L g1009 ( .A(n_918), .Y(n_1009) );
OR2x6_ASAP7_75t_L g1010 ( .A(n_888), .B(n_909), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_904), .B(n_890), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_887), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_840), .B(n_871), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_871), .B(n_867), .Y(n_1014) );
INVxp67_ASAP7_75t_SL g1015 ( .A(n_921), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_887), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_937), .B(n_854), .Y(n_1017) );
AND2x4_ASAP7_75t_L g1018 ( .A(n_915), .B(n_893), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_854), .Y(n_1019) );
INVx3_ASAP7_75t_L g1020 ( .A(n_866), .Y(n_1020) );
INVx2_ASAP7_75t_L g1021 ( .A(n_860), .Y(n_1021) );
OR2x2_ASAP7_75t_SL g1022 ( .A(n_841), .B(n_838), .Y(n_1022) );
NOR2xp33_ASAP7_75t_L g1023 ( .A(n_945), .B(n_930), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_928), .Y(n_1024) );
INVx2_ASAP7_75t_L g1025 ( .A(n_899), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_834), .B(n_849), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_927), .Y(n_1027) );
BUFx3_ASAP7_75t_L g1028 ( .A(n_898), .Y(n_1028) );
HB1xp67_ASAP7_75t_L g1029 ( .A(n_844), .Y(n_1029) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_878), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_926), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_932), .B(n_946), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_842), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_936), .B(n_944), .Y(n_1034) );
BUFx3_ASAP7_75t_L g1035 ( .A(n_853), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_899), .A2(n_949), .B1(n_935), .B2(n_934), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_971), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_971), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_953), .B(n_922), .Y(n_1039) );
NOR3xp33_ASAP7_75t_L g1040 ( .A(n_1023), .B(n_876), .C(n_916), .Y(n_1040) );
OR2x2_ASAP7_75t_L g1041 ( .A(n_970), .B(n_908), .Y(n_1041) );
OR2x2_ASAP7_75t_L g1042 ( .A(n_970), .B(n_877), .Y(n_1042) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_973), .B(n_850), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_974), .B(n_868), .Y(n_1044) );
OAI22xp5_ASAP7_75t_SL g1045 ( .A1(n_1004), .A2(n_896), .B1(n_850), .B2(n_874), .Y(n_1045) );
INVx2_ASAP7_75t_SL g1046 ( .A(n_1001), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_961), .Y(n_1047) );
OAI31xp33_ASAP7_75t_SL g1048 ( .A1(n_986), .A2(n_924), .A3(n_863), .B(n_912), .Y(n_1048) );
INVx3_ASAP7_75t_SL g1049 ( .A(n_1001), .Y(n_1049) );
BUFx2_ASAP7_75t_L g1050 ( .A(n_952), .Y(n_1050) );
HB1xp67_ASAP7_75t_L g1051 ( .A(n_953), .Y(n_1051) );
OR2x2_ASAP7_75t_L g1052 ( .A(n_973), .B(n_980), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_953), .B(n_958), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_958), .B(n_974), .Y(n_1054) );
BUFx2_ASAP7_75t_L g1055 ( .A(n_965), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_961), .Y(n_1056) );
INVx5_ASAP7_75t_L g1057 ( .A(n_1001), .Y(n_1057) );
OR2x2_ASAP7_75t_L g1058 ( .A(n_980), .B(n_1031), .Y(n_1058) );
BUFx3_ASAP7_75t_L g1059 ( .A(n_1001), .Y(n_1059) );
AND2x4_ASAP7_75t_L g1060 ( .A(n_958), .B(n_959), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_996), .B(n_1031), .Y(n_1061) );
INVx5_ASAP7_75t_L g1062 ( .A(n_1001), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_972), .B(n_976), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_963), .Y(n_1064) );
BUFx3_ASAP7_75t_L g1065 ( .A(n_1001), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_972), .B(n_976), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_996), .B(n_978), .Y(n_1067) );
NAND2xp33_ASAP7_75t_L g1068 ( .A(n_1014), .B(n_1001), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_964), .A2(n_1034), .B1(n_998), .B2(n_1032), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_996), .B(n_978), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_963), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_966), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_995), .Y(n_1073) );
OR2x2_ASAP7_75t_L g1074 ( .A(n_954), .B(n_959), .Y(n_1074) );
NAND4xp25_ASAP7_75t_L g1075 ( .A(n_964), .B(n_1036), .C(n_1032), .D(n_1034), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_978), .B(n_954), .Y(n_1076) );
INVx4_ASAP7_75t_L g1077 ( .A(n_965), .Y(n_1077) );
AOI22xp5_ASAP7_75t_L g1078 ( .A1(n_1036), .A2(n_1005), .B1(n_1011), .B2(n_1003), .Y(n_1078) );
OR2x2_ASAP7_75t_L g1079 ( .A(n_1027), .B(n_952), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1027), .B(n_956), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_966), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_968), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_956), .B(n_957), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_957), .B(n_992), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_968), .Y(n_1085) );
BUFx2_ASAP7_75t_L g1086 ( .A(n_965), .Y(n_1086) );
AND2x6_ASAP7_75t_L g1087 ( .A(n_975), .B(n_1019), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_979), .Y(n_1088) );
INVx3_ASAP7_75t_L g1089 ( .A(n_1006), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_979), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1005), .B(n_1003), .Y(n_1091) );
INVx3_ASAP7_75t_L g1092 ( .A(n_1006), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1011), .B(n_962), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_962), .B(n_990), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_990), .B(n_987), .Y(n_1095) );
NOR3xp33_ASAP7_75t_L g1096 ( .A(n_1020), .B(n_1013), .C(n_1026), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_992), .B(n_1024), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_981), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_987), .B(n_1025), .Y(n_1099) );
BUFx3_ASAP7_75t_L g1100 ( .A(n_994), .Y(n_1100) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_960), .Y(n_1101) );
AOI211xp5_ASAP7_75t_L g1102 ( .A1(n_986), .A2(n_955), .B(n_1017), .C(n_1014), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_982), .Y(n_1103) );
INVx1_ASAP7_75t_SL g1104 ( .A(n_1004), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1025), .B(n_1030), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_982), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_984), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1024), .B(n_975), .Y(n_1108) );
BUFx2_ASAP7_75t_L g1109 ( .A(n_1051), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1047), .Y(n_1110) );
AND2x4_ASAP7_75t_SL g1111 ( .A(n_1077), .B(n_1020), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1067), .B(n_975), .Y(n_1112) );
AOI33xp33_ASAP7_75t_L g1113 ( .A1(n_1069), .A2(n_1013), .A3(n_1017), .B1(n_997), .B2(n_1026), .B3(n_1025), .Y(n_1113) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1073), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1056), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1070), .B(n_1002), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_1054), .B(n_1002), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_1054), .B(n_1007), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1037), .B(n_997), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1070), .B(n_1007), .Y(n_1120) );
INVx3_ASAP7_75t_L g1121 ( .A(n_1057), .Y(n_1121) );
AND2x6_ASAP7_75t_SL g1122 ( .A(n_1091), .B(n_955), .Y(n_1122) );
AND2x4_ASAP7_75t_L g1123 ( .A(n_1060), .B(n_1018), .Y(n_1123) );
INVx2_ASAP7_75t_SL g1124 ( .A(n_1057), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1038), .B(n_1000), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1053), .B(n_1018), .Y(n_1126) );
INVx3_ASAP7_75t_L g1127 ( .A(n_1057), .Y(n_1127) );
OAI221xp5_ASAP7_75t_L g1128 ( .A1(n_1078), .A2(n_1030), .B1(n_1000), .B2(n_1028), .C(n_1033), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1053), .B(n_1018), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1098), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1074), .Y(n_1131) );
O2A1O1Ixp33_ASAP7_75t_L g1132 ( .A1(n_1075), .A2(n_1033), .B(n_1020), .C(n_1030), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1108), .B(n_1018), .Y(n_1133) );
AND2x4_ASAP7_75t_L g1134 ( .A(n_1060), .B(n_1012), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1108), .B(n_985), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1084), .B(n_985), .Y(n_1136) );
NOR2xp33_ASAP7_75t_L g1137 ( .A(n_1093), .B(n_1028), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1074), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1084), .B(n_983), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1083), .B(n_969), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1061), .B(n_983), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1083), .B(n_969), .Y(n_1142) );
OR2x6_ASAP7_75t_L g1143 ( .A(n_1050), .B(n_1010), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1061), .B(n_989), .Y(n_1144) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_1052), .B(n_988), .Y(n_1145) );
OAI21xp33_ASAP7_75t_L g1146 ( .A1(n_1102), .A2(n_1035), .B(n_1015), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1064), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1097), .B(n_989), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1097), .B(n_1016), .Y(n_1149) );
AND2x4_ASAP7_75t_L g1150 ( .A(n_1060), .B(n_1012), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1080), .B(n_1016), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1071), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1080), .B(n_1015), .Y(n_1153) );
NOR2xp33_ASAP7_75t_L g1154 ( .A(n_1063), .B(n_1028), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1076), .B(n_1010), .Y(n_1155) );
NAND2xp5_ASAP7_75t_SL g1156 ( .A(n_1104), .B(n_994), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1076), .B(n_1010), .Y(n_1157) );
AND2x2_ASAP7_75t_SL g1158 ( .A(n_1068), .B(n_960), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1039), .B(n_1010), .Y(n_1159) );
HB1xp67_ASAP7_75t_L g1160 ( .A(n_1050), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1072), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1081), .Y(n_1162) );
OR2x2_ASAP7_75t_L g1163 ( .A(n_1058), .B(n_1008), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1039), .B(n_1010), .Y(n_1164) );
AND2x4_ASAP7_75t_L g1165 ( .A(n_1087), .B(n_1010), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_1131), .B(n_1095), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1130), .Y(n_1167) );
INVx3_ASAP7_75t_L g1168 ( .A(n_1121), .Y(n_1168) );
NAND2x1_ASAP7_75t_L g1169 ( .A(n_1121), .B(n_999), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1130), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1161), .Y(n_1171) );
NOR3xp33_ASAP7_75t_SL g1172 ( .A(n_1128), .B(n_1045), .C(n_1044), .Y(n_1172) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1114), .Y(n_1173) );
BUFx2_ASAP7_75t_L g1174 ( .A(n_1121), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1133), .B(n_1112), .Y(n_1175) );
NOR2xp33_ASAP7_75t_L g1176 ( .A(n_1122), .B(n_1066), .Y(n_1176) );
INVx1_ASAP7_75t_SL g1177 ( .A(n_1111), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1126), .B(n_1101), .Y(n_1178) );
INVx1_ASAP7_75t_SL g1179 ( .A(n_1111), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1126), .B(n_1129), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1131), .B(n_1103), .Y(n_1181) );
NOR2xp33_ASAP7_75t_SL g1182 ( .A(n_1124), .B(n_1057), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1129), .B(n_1101), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1117), .B(n_1079), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1133), .B(n_1087), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1117), .B(n_1079), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1161), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1162), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1162), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1110), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1115), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1138), .B(n_1136), .Y(n_1192) );
AOI221xp5_ASAP7_75t_L g1193 ( .A1(n_1154), .A2(n_1094), .B1(n_1082), .B2(n_1085), .C(n_1096), .Y(n_1193) );
AND2x2_ASAP7_75t_SL g1194 ( .A(n_1158), .B(n_1068), .Y(n_1194) );
OAI22xp33_ASAP7_75t_L g1195 ( .A1(n_1127), .A2(n_1057), .B1(n_1062), .B2(n_1049), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1138), .B(n_1106), .Y(n_1196) );
NOR2xp33_ASAP7_75t_L g1197 ( .A(n_1132), .B(n_1099), .Y(n_1197) );
NAND2xp5_ASAP7_75t_SL g1198 ( .A(n_1158), .B(n_1062), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1112), .B(n_1087), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1118), .B(n_1058), .Y(n_1200) );
AND2x4_ASAP7_75t_L g1201 ( .A(n_1165), .B(n_1087), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1136), .B(n_1107), .Y(n_1202) );
O2A1O1Ixp33_ASAP7_75t_L g1203 ( .A1(n_1146), .A2(n_1040), .B(n_1020), .C(n_1029), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1147), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1152), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1163), .Y(n_1206) );
OAI21xp33_ASAP7_75t_L g1207 ( .A1(n_1113), .A2(n_1048), .B(n_1105), .Y(n_1207) );
OAI211xp5_ASAP7_75t_L g1208 ( .A1(n_1137), .A2(n_994), .B(n_1077), .C(n_1062), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1163), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1139), .B(n_1088), .Y(n_1210) );
AOI221x1_ASAP7_75t_L g1211 ( .A1(n_1176), .A2(n_1127), .B1(n_1077), .B2(n_1089), .C(n_1092), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g1212 ( .A1(n_1207), .A2(n_1125), .B1(n_1142), .B2(n_1140), .C(n_1139), .Y(n_1212) );
AOI21xp5_ASAP7_75t_L g1213 ( .A1(n_1198), .A2(n_1124), .B(n_1156), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1214 ( .A(n_1174), .Y(n_1214) );
INVx2_ASAP7_75t_L g1215 ( .A(n_1173), .Y(n_1215) );
NOR2x1_ASAP7_75t_L g1216 ( .A(n_1169), .B(n_1127), .Y(n_1216) );
OAI321xp33_ASAP7_75t_L g1217 ( .A1(n_1198), .A2(n_1143), .A3(n_1153), .B1(n_1119), .B2(n_1164), .C(n_1159), .Y(n_1217) );
NOR2xp33_ASAP7_75t_L g1218 ( .A(n_1176), .B(n_1145), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1190), .Y(n_1219) );
AOI21xp33_ASAP7_75t_SL g1220 ( .A1(n_1194), .A2(n_1049), .B(n_1046), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1191), .Y(n_1221) );
AOI21xp5_ASAP7_75t_L g1222 ( .A1(n_1194), .A2(n_1062), .B(n_1046), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1206), .B(n_1135), .Y(n_1223) );
NOR2xp33_ASAP7_75t_L g1224 ( .A(n_1197), .B(n_1145), .Y(n_1224) );
INVx2_ASAP7_75t_SL g1225 ( .A(n_1177), .Y(n_1225) );
NOR4xp75_ASAP7_75t_L g1226 ( .A(n_1168), .B(n_1153), .C(n_999), .D(n_1164), .Y(n_1226) );
OR2x2_ASAP7_75t_L g1227 ( .A(n_1184), .B(n_1118), .Y(n_1227) );
AOI321xp33_ASAP7_75t_L g1228 ( .A1(n_1197), .A2(n_1159), .A3(n_1141), .B1(n_1144), .B2(n_1148), .C(n_1135), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1175), .B(n_1155), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1204), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1175), .B(n_1155), .Y(n_1231) );
NAND2xp5_ASAP7_75t_SL g1232 ( .A(n_1195), .B(n_1109), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1205), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1180), .B(n_1157), .Y(n_1234) );
INVxp67_ASAP7_75t_L g1235 ( .A(n_1179), .Y(n_1235) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_1193), .A2(n_1143), .B1(n_1062), .B2(n_1123), .Y(n_1236) );
NOR3xp33_ASAP7_75t_SL g1237 ( .A(n_1203), .B(n_1090), .C(n_991), .Y(n_1237) );
AOI21xp33_ASAP7_75t_SL g1238 ( .A1(n_1195), .A2(n_1143), .B(n_1165), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1167), .Y(n_1239) );
INVxp67_ASAP7_75t_L g1240 ( .A(n_1209), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1227), .B(n_1192), .Y(n_1241) );
NAND2x1p5_ASAP7_75t_L g1242 ( .A(n_1216), .B(n_1168), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1219), .Y(n_1243) );
OAI211xp5_ASAP7_75t_SL g1244 ( .A1(n_1212), .A2(n_1172), .B(n_1166), .C(n_1210), .Y(n_1244) );
INVxp67_ASAP7_75t_SL g1245 ( .A(n_1214), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1221), .Y(n_1246) );
OAI21xp33_ASAP7_75t_L g1247 ( .A1(n_1224), .A2(n_1172), .B(n_1199), .Y(n_1247) );
OAI221xp5_ASAP7_75t_SL g1248 ( .A1(n_1228), .A2(n_1199), .B1(n_1143), .B2(n_1185), .C(n_1208), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1224), .B(n_1202), .Y(n_1249) );
NAND3xp33_ASAP7_75t_L g1250 ( .A(n_1237), .B(n_1160), .C(n_1168), .Y(n_1250) );
NAND3xp33_ASAP7_75t_L g1251 ( .A(n_1232), .B(n_1182), .C(n_1170), .Y(n_1251) );
AOI221xp5_ASAP7_75t_L g1252 ( .A1(n_1218), .A2(n_1181), .B1(n_1196), .B2(n_1189), .C(n_1171), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1229), .B(n_1201), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1230), .Y(n_1254) );
NAND2x1_ASAP7_75t_L g1255 ( .A(n_1225), .B(n_1201), .Y(n_1255) );
HB1xp67_ASAP7_75t_L g1256 ( .A(n_1225), .Y(n_1256) );
AOI22xp5_ASAP7_75t_L g1257 ( .A1(n_1236), .A2(n_1201), .B1(n_1185), .B2(n_1087), .Y(n_1257) );
NOR4xp25_ASAP7_75t_L g1258 ( .A(n_1232), .B(n_1188), .C(n_1187), .D(n_984), .Y(n_1258) );
OAI221xp5_ASAP7_75t_L g1259 ( .A1(n_1238), .A2(n_1186), .B1(n_1200), .B2(n_1035), .C(n_1029), .Y(n_1259) );
AOI321xp33_ASAP7_75t_L g1260 ( .A1(n_1217), .A2(n_1148), .A3(n_1141), .B1(n_1144), .B2(n_1178), .C(n_1183), .Y(n_1260) );
OAI22xp5_ASAP7_75t_L g1261 ( .A1(n_1248), .A2(n_1235), .B1(n_1220), .B2(n_1218), .Y(n_1261) );
NAND5xp2_ASAP7_75t_L g1262 ( .A(n_1260), .B(n_1222), .C(n_1213), .D(n_977), .E(n_1055), .Y(n_1262) );
CKINVDCx5p33_ASAP7_75t_R g1263 ( .A(n_1256), .Y(n_1263) );
NOR3xp33_ASAP7_75t_L g1264 ( .A(n_1251), .B(n_1240), .C(n_1233), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1243), .Y(n_1265) );
OAI31xp33_ASAP7_75t_L g1266 ( .A1(n_1247), .A2(n_1231), .A3(n_1229), .B(n_1234), .Y(n_1266) );
AOI221xp5_ASAP7_75t_L g1267 ( .A1(n_1258), .A2(n_1223), .B1(n_1239), .B2(n_1231), .C(n_1234), .Y(n_1267) );
AOI322xp5_ASAP7_75t_L g1268 ( .A1(n_1249), .A2(n_1157), .A3(n_1149), .B1(n_1165), .B2(n_1151), .C1(n_1120), .C2(n_1116), .Y(n_1268) );
OAI211xp5_ASAP7_75t_L g1269 ( .A1(n_1258), .A2(n_1211), .B(n_1035), .C(n_1086), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1246), .Y(n_1270) );
INVx2_ASAP7_75t_L g1271 ( .A(n_1242), .Y(n_1271) );
NOR2xp33_ASAP7_75t_R g1272 ( .A(n_1254), .B(n_1059), .Y(n_1272) );
OAI21xp33_ASAP7_75t_L g1273 ( .A1(n_1244), .A2(n_1123), .B(n_1149), .Y(n_1273) );
AOI22xp5_ASAP7_75t_L g1274 ( .A1(n_1261), .A2(n_1259), .B1(n_1257), .B2(n_1245), .Y(n_1274) );
INVxp67_ASAP7_75t_L g1275 ( .A(n_1263), .Y(n_1275) );
OAI211xp5_ASAP7_75t_SL g1276 ( .A1(n_1266), .A2(n_1252), .B(n_1250), .C(n_1241), .Y(n_1276) );
AOI21xp5_ASAP7_75t_L g1277 ( .A1(n_1262), .A2(n_1255), .B(n_1242), .Y(n_1277) );
OAI211xp5_ASAP7_75t_SL g1278 ( .A1(n_1267), .A2(n_1043), .B(n_1042), .C(n_1041), .Y(n_1278) );
NAND2xp5_ASAP7_75t_SL g1279 ( .A(n_1272), .B(n_1253), .Y(n_1279) );
O2A1O1Ixp33_ASAP7_75t_L g1280 ( .A1(n_1264), .A2(n_1021), .B(n_1042), .C(n_977), .Y(n_1280) );
XOR2xp5_ASAP7_75t_L g1281 ( .A(n_1265), .B(n_1134), .Y(n_1281) );
A2O1A1Ixp33_ASAP7_75t_L g1282 ( .A1(n_1269), .A2(n_1123), .B(n_1065), .C(n_1059), .Y(n_1282) );
NOR3xp33_ASAP7_75t_SL g1283 ( .A(n_1276), .B(n_1273), .C(n_1270), .Y(n_1283) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1275), .Y(n_1284) );
NOR3x2_ASAP7_75t_L g1285 ( .A(n_1277), .B(n_1272), .C(n_1271), .Y(n_1285) );
NAND3xp33_ASAP7_75t_SL g1286 ( .A(n_1274), .B(n_1268), .C(n_1271), .Y(n_1286) );
OAI21xp5_ASAP7_75t_L g1287 ( .A1(n_1282), .A2(n_1021), .B(n_1043), .Y(n_1287) );
NOR3xp33_ASAP7_75t_SL g1288 ( .A(n_1278), .B(n_1226), .C(n_991), .Y(n_1288) );
AOI22xp5_ASAP7_75t_L g1289 ( .A1(n_1286), .A2(n_1279), .B1(n_1281), .B2(n_1087), .Y(n_1289) );
AND2x4_ASAP7_75t_L g1290 ( .A(n_1284), .B(n_1134), .Y(n_1290) );
O2A1O1Ixp33_ASAP7_75t_L g1291 ( .A1(n_1283), .A2(n_1280), .B(n_1021), .C(n_1019), .Y(n_1291) );
NAND3xp33_ASAP7_75t_L g1292 ( .A(n_1288), .B(n_1215), .C(n_1009), .Y(n_1292) );
AND2x4_ASAP7_75t_L g1293 ( .A(n_1287), .B(n_1150), .Y(n_1293) );
OR3x2_ASAP7_75t_L g1294 ( .A(n_1289), .B(n_1285), .C(n_1041), .Y(n_1294) );
BUFx2_ASAP7_75t_L g1295 ( .A(n_1290), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1292), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1291), .Y(n_1297) );
OAI22xp5_ASAP7_75t_SL g1298 ( .A1(n_1297), .A2(n_1293), .B1(n_1022), .B2(n_1065), .Y(n_1298) );
INVx2_ASAP7_75t_L g1299 ( .A(n_1295), .Y(n_1299) );
OAI22xp5_ASAP7_75t_SL g1300 ( .A1(n_1296), .A2(n_1022), .B1(n_1100), .B2(n_967), .Y(n_1300) );
AOI22xp5_ASAP7_75t_L g1301 ( .A1(n_1299), .A2(n_1294), .B1(n_1298), .B2(n_1300), .Y(n_1301) );
XNOR2xp5_ASAP7_75t_L g1302 ( .A(n_1299), .B(n_1294), .Y(n_1302) );
AOI21xp5_ASAP7_75t_L g1303 ( .A1(n_1302), .A2(n_993), .B(n_1009), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1303), .B(n_1301), .Y(n_1304) );
AOI21xp5_ASAP7_75t_L g1305 ( .A1(n_1304), .A2(n_993), .B(n_1009), .Y(n_1305) );
endmodule