module fake_ibex_569_n_998 (n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_998);

input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_998;

wire n_151;
wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_992;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_947;
wire n_981;
wire n_972;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_153;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_317;
wire n_375;
wire n_280;
wire n_340;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_154;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_158;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_732;
wire n_673;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_982;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_968;
wire n_625;
wire n_953;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_607;
wire n_427;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_689;
wire n_960;
wire n_793;
wire n_167;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_648;
wire n_229;
wire n_209;
wire n_472;
wire n_571;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_444;
wire n_200;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_379;
wire n_320;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_858;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_164;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_890;
wire n_874;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_21),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_50),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_43),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g162 ( 
.A(n_58),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_2),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g164 ( 
.A(n_53),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_137),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_73),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_49),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_75),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_38),
.B(n_34),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_86),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_62),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_41),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_23),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_48),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_29),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_11),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_52),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_111),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_57),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_84),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_89),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_31),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_61),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_0),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_18),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_28),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_17),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_149),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_82),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_22),
.Y(n_198)
);

INVxp33_ASAP7_75t_SL g199 ( 
.A(n_17),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_56),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_72),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_35),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_88),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_100),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_114),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_78),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g209 ( 
.A(n_6),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_67),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_101),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_8),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_12),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_10),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_32),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_92),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_7),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_104),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_22),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_37),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_106),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_24),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_51),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_4),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_54),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_96),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_144),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_36),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_68),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_109),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_116),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_135),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_40),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_18),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_12),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_7),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_125),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_123),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_20),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_117),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_115),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_19),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g243 ( 
.A(n_13),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_85),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_30),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_19),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_133),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_1),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g250 ( 
.A(n_42),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_6),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_131),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_174),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_217),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_174),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_159),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_175),
.Y(n_257)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_0),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_175),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_212),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_183),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_159),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_226),
.Y(n_264)
);

AND2x6_ASAP7_75t_L g265 ( 
.A(n_173),
.B(n_27),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_183),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_206),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_153),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_155),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_213),
.B(n_1),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_245),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

AND3x2_ASAP7_75t_L g277 ( 
.A(n_172),
.B(n_2),
.C(n_3),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_211),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_169),
.B(n_3),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_183),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_150),
.Y(n_281)
);

CKINVDCx8_ASAP7_75t_R g282 ( 
.A(n_156),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_183),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_151),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_152),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_197),
.B(n_4),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_154),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_157),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_244),
.B(n_8),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_178),
.B(n_9),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_158),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_221),
.B(n_9),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_153),
.B(n_10),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_186),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_160),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_167),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_168),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_L g299 ( 
.A(n_156),
.B(n_148),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_170),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_177),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_179),
.B(n_11),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_180),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_183),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_181),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_163),
.B(n_13),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_182),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_184),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_172),
.B(n_14),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_163),
.B(n_214),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_185),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_214),
.B(n_14),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_187),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_219),
.B(n_15),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_219),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_224),
.B(n_15),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_224),
.B(n_16),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_186),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_234),
.B(n_16),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_188),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_189),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_190),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_200),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_202),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_234),
.B(n_20),
.Y(n_325)
);

OA21x2_ASAP7_75t_L g326 ( 
.A1(n_203),
.A2(n_215),
.B(n_207),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_196),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_204),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_251),
.B(n_21),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_236),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_205),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_208),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_192),
.B(n_23),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_216),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_309),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_260),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_315),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_271),
.B(n_161),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

AND2x6_ASAP7_75t_L g341 ( 
.A(n_273),
.B(n_173),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_253),
.A2(n_198),
.B1(n_222),
.B2(n_249),
.Y(n_342)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_265),
.Y(n_343)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_265),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_309),
.Y(n_345)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_265),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_309),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_193),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_253),
.B(n_218),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_333),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_269),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_254),
.B(n_251),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_255),
.B(n_220),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_270),
.B(n_165),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_265),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_279),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_273),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_255),
.B(n_225),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_260),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_260),
.Y(n_361)
);

AND2x2_ASAP7_75t_SL g362 ( 
.A(n_273),
.B(n_236),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_265),
.B(n_196),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_265),
.Y(n_364)
);

AND2x6_ASAP7_75t_L g365 ( 
.A(n_273),
.B(n_227),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_257),
.B(n_228),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_257),
.B(n_232),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_333),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_310),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_304),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_314),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_321),
.B(n_201),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_321),
.B(n_233),
.Y(n_375)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_265),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_279),
.B(n_165),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_259),
.B(n_241),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_259),
.B(n_281),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_282),
.B(n_223),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_256),
.Y(n_381)
);

BUFx10_ASAP7_75t_L g382 ( 
.A(n_264),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_304),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_256),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_287),
.B(n_195),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_256),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_260),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_295),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_263),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_263),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_263),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_287),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_260),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_318),
.B(n_223),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_268),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_327),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_266),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_266),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_268),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_266),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_281),
.B(n_292),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_314),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_276),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_276),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_293),
.B(n_248),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_304),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g407 ( 
.A(n_316),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_278),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_316),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_293),
.B(n_239),
.Y(n_410)
);

OAI21xp33_ASAP7_75t_L g411 ( 
.A1(n_292),
.A2(n_250),
.B(n_247),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_266),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_266),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_296),
.B(n_171),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_282),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_278),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_262),
.Y(n_417)
);

AO22x2_ASAP7_75t_L g418 ( 
.A1(n_296),
.A2(n_209),
.B1(n_243),
.B2(n_242),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_300),
.B(n_236),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_283),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_300),
.B(n_236),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_285),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_283),
.Y(n_423)
);

INVx8_ASAP7_75t_L g424 ( 
.A(n_262),
.Y(n_424)
);

NAND2x1p5_ASAP7_75t_L g425 ( 
.A(n_290),
.B(n_236),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_285),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_262),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_301),
.B(n_171),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_326),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_262),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_267),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_326),
.Y(n_432)
);

OR2x2_ASAP7_75t_SL g433 ( 
.A(n_294),
.B(n_199),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_326),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_288),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_267),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_288),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_288),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_289),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_301),
.B(n_194),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_289),
.Y(n_441)
);

BUFx10_ASAP7_75t_L g442 ( 
.A(n_307),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_306),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_307),
.B(n_194),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_313),
.B(n_231),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_312),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_421),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_419),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_442),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_442),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_365),
.A2(n_326),
.B1(n_328),
.B2(n_289),
.Y(n_451)
);

AND2x2_ASAP7_75t_SL g452 ( 
.A(n_363),
.B(n_299),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_435),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_422),
.B(n_231),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_379),
.B(n_285),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_395),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_379),
.B(n_313),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_392),
.B(n_317),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_437),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_320),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_395),
.Y(n_461)
);

BUFx4f_ASAP7_75t_L g462 ( 
.A(n_362),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_446),
.B(n_250),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_403),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_338),
.B(n_319),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_440),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_338),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_415),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_388),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_439),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_344),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_R g473 ( 
.A(n_380),
.B(n_237),
.Y(n_473)
);

NAND3xp33_ASAP7_75t_L g474 ( 
.A(n_339),
.B(n_325),
.C(n_329),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_403),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_441),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_371),
.B(n_320),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_341),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_401),
.Y(n_480)
);

BUFx12f_ASAP7_75t_L g481 ( 
.A(n_382),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_373),
.B(n_291),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_373),
.B(n_322),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_446),
.B(n_322),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_402),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_404),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_404),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_382),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_341),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_385),
.B(n_323),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_401),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_362),
.B(n_323),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_344),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_341),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_409),
.B(n_324),
.Y(n_495)
);

BUFx4f_ASAP7_75t_SL g496 ( 
.A(n_341),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_385),
.B(n_324),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_339),
.B(n_331),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_357),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_357),
.B(n_331),
.Y(n_500)
);

CKINVDCx14_ASAP7_75t_R g501 ( 
.A(n_394),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_399),
.Y(n_502)
);

CKINVDCx14_ASAP7_75t_R g503 ( 
.A(n_396),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_410),
.B(n_348),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_414),
.B(n_332),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_352),
.A2(n_199),
.B1(n_240),
.B2(n_238),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_407),
.B(n_332),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_408),
.Y(n_508)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_400),
.Y(n_510)
);

O2A1O1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_349),
.A2(n_274),
.B(n_261),
.C(n_272),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_356),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_400),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_335),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_354),
.Y(n_515)
);

AND3x1_ASAP7_75t_L g516 ( 
.A(n_380),
.B(n_258),
.C(n_334),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_343),
.B(n_286),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_343),
.B(n_286),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_416),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_414),
.B(n_297),
.Y(n_520)
);

NAND2x1p5_ASAP7_75t_L g521 ( 
.A(n_377),
.B(n_302),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_407),
.B(n_334),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_420),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_443),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_423),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_381),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_428),
.B(n_328),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_433),
.B(n_297),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_418),
.A2(n_237),
.B1(n_240),
.B2(n_238),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_443),
.Y(n_530)
);

AO22x1_ASAP7_75t_L g531 ( 
.A1(n_405),
.A2(n_258),
.B1(n_164),
.B2(n_166),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_434),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_348),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_384),
.Y(n_534)
);

CKINVDCx11_ASAP7_75t_R g535 ( 
.A(n_410),
.Y(n_535)
);

O2A1O1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_349),
.A2(n_275),
.B(n_272),
.C(n_261),
.Y(n_536)
);

INVx3_ASAP7_75t_SL g537 ( 
.A(n_405),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_386),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_428),
.B(n_298),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_389),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_390),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_391),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_351),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_445),
.B(n_277),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_445),
.Y(n_545)
);

BUFx12f_ASAP7_75t_L g546 ( 
.A(n_425),
.Y(n_546)
);

BUFx12f_ASAP7_75t_L g547 ( 
.A(n_425),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_335),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_358),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_434),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_405),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_468),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_480),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_491),
.B(n_405),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_481),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_472),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_535),
.Y(n_557)
);

OAI21x1_ASAP7_75t_SL g558 ( 
.A1(n_479),
.A2(n_364),
.B(n_356),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_532),
.A2(n_364),
.B(n_376),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_514),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_545),
.B(n_405),
.Y(n_561)
);

OR2x6_ASAP7_75t_L g562 ( 
.A(n_488),
.B(n_450),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_545),
.B(n_484),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_457),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_524),
.B(n_418),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_450),
.B(n_449),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_469),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_514),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_524),
.B(n_376),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_457),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_548),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_548),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_468),
.Y(n_573)
);

INVx3_ASAP7_75t_SL g574 ( 
.A(n_543),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_509),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_549),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_479),
.B(n_418),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_550),
.A2(n_346),
.B(n_343),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_447),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_472),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_447),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_550),
.A2(n_346),
.B(n_343),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_544),
.B(n_490),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_530),
.B(n_411),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_473),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_485),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_483),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_483),
.Y(n_588)
);

BUFx12f_ASAP7_75t_L g589 ( 
.A(n_470),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_515),
.B(n_363),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_490),
.Y(n_591)
);

AOI221xp5_ASAP7_75t_L g592 ( 
.A1(n_500),
.A2(n_342),
.B1(n_275),
.B2(n_274),
.C(n_353),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_509),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_509),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_484),
.B(n_350),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_472),
.Y(n_596)
);

BUFx4f_ASAP7_75t_SL g597 ( 
.A(n_546),
.Y(n_597)
);

O2A1O1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_498),
.A2(n_485),
.B(n_499),
.C(n_500),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_493),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_529),
.B(n_353),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_489),
.B(n_358),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_489),
.B(n_529),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_493),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_505),
.A2(n_432),
.B(n_429),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_547),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_497),
.Y(n_606)
);

OAI221xp5_ASAP7_75t_L g607 ( 
.A1(n_498),
.A2(n_342),
.B1(n_366),
.B2(n_368),
.C(n_367),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_493),
.A2(n_370),
.B(n_369),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_466),
.B(n_366),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_494),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_505),
.B(n_341),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_503),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_504),
.B(n_467),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_504),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_512),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_537),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_520),
.A2(n_365),
.B1(n_347),
.B2(n_345),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_497),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_462),
.A2(n_365),
.B1(n_347),
.B2(n_345),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_462),
.A2(n_365),
.B1(n_432),
.B2(n_429),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_455),
.A2(n_537),
.B1(n_451),
.B2(n_527),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_507),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_501),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_482),
.B(n_374),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_482),
.A2(n_365),
.B1(n_375),
.B2(n_374),
.Y(n_625)
);

BUFx4f_ASAP7_75t_L g626 ( 
.A(n_533),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_492),
.A2(n_375),
.B1(n_359),
.B2(n_378),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_551),
.B(n_368),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_464),
.B(n_458),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_494),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_455),
.A2(n_328),
.B1(n_378),
.B2(n_359),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_522),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_544),
.A2(n_426),
.B1(n_346),
.B2(n_308),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_506),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_495),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_512),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_534),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_448),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_541),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_525),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_502),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_527),
.A2(n_424),
.B(n_360),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_477),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_494),
.Y(n_644)
);

BUFx12f_ASAP7_75t_L g645 ( 
.A(n_528),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_L g646 ( 
.A1(n_496),
.A2(n_311),
.B1(n_298),
.B2(n_303),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_486),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_496),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_477),
.B(n_303),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_508),
.Y(n_650)
);

NOR2xp67_ASAP7_75t_SL g651 ( 
.A(n_494),
.B(n_305),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_519),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_523),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_486),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_460),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_451),
.A2(n_305),
.B1(n_308),
.B2(n_311),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_512),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_460),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_478),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_487),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_487),
.Y(n_661)
);

O2A1O1Ixp33_ASAP7_75t_SL g662 ( 
.A1(n_517),
.A2(n_162),
.B(n_176),
.C(n_191),
.Y(n_662)
);

AOI221xp5_ASAP7_75t_L g663 ( 
.A1(n_655),
.A2(n_536),
.B1(n_511),
.B2(n_539),
.C(n_520),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_657),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_563),
.A2(n_458),
.B1(n_516),
.B2(n_474),
.Y(n_665)
);

INVx6_ASAP7_75t_L g666 ( 
.A(n_657),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_553),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_564),
.A2(n_452),
.B1(n_539),
.B2(n_540),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_SL g669 ( 
.A1(n_577),
.A2(n_452),
.B1(n_521),
.B2(n_471),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_570),
.A2(n_542),
.B1(n_538),
.B2(n_526),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_563),
.A2(n_459),
.B1(n_453),
.B2(n_463),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_638),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_609),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_552),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_577),
.A2(n_476),
.B1(n_521),
.B2(n_465),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_641),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_607),
.A2(n_536),
.B1(n_511),
.B2(n_456),
.Y(n_677)
);

AO31x2_ASAP7_75t_L g678 ( 
.A1(n_621),
.A2(n_604),
.A3(n_656),
.B(n_631),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_597),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_573),
.Y(n_680)
);

O2A1O1Ixp33_ASAP7_75t_SL g681 ( 
.A1(n_595),
.A2(n_518),
.B(n_454),
.C(n_230),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_658),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_555),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_650),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_586),
.B(n_461),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_607),
.A2(n_475),
.B1(n_210),
.B2(n_246),
.Y(n_686)
);

OAI221xp5_ASAP7_75t_L g687 ( 
.A1(n_598),
.A2(n_267),
.B1(n_280),
.B2(n_284),
.C(n_330),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_565),
.B(n_531),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_652),
.Y(n_689)
);

AO21x2_ASAP7_75t_L g690 ( 
.A1(n_604),
.A2(n_398),
.B(n_361),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_L g691 ( 
.A(n_621),
.B(n_510),
.Y(n_691)
);

AOI221xp5_ASAP7_75t_L g692 ( 
.A1(n_635),
.A2(n_267),
.B1(n_284),
.B2(n_280),
.C(n_330),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_653),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_622),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_624),
.B(n_24),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_591),
.Y(n_696)
);

AO22x2_ASAP7_75t_L g697 ( 
.A1(n_600),
.A2(n_25),
.B1(n_26),
.B2(n_413),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_640),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_577),
.A2(n_280),
.B1(n_284),
.B2(n_330),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_602),
.A2(n_280),
.B1(n_284),
.B2(n_330),
.Y(n_700)
);

NOR2xp67_ASAP7_75t_L g701 ( 
.A(n_589),
.B(n_25),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_606),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_617),
.A2(n_513),
.B1(n_424),
.B2(n_412),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_595),
.B(n_397),
.Y(n_704)
);

CKINVDCx6p67_ASAP7_75t_R g705 ( 
.A(n_574),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_637),
.Y(n_706)
);

AOI221xp5_ASAP7_75t_L g707 ( 
.A1(n_592),
.A2(n_436),
.B1(n_431),
.B2(n_430),
.C(n_427),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_632),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_659),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_639),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_587),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_617),
.A2(n_393),
.B1(n_387),
.B2(n_336),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_611),
.A2(n_430),
.B1(n_427),
.B2(n_417),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_576),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_605),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_562),
.Y(n_716)
);

AO31x2_ASAP7_75t_L g717 ( 
.A1(n_656),
.A2(n_26),
.A3(n_406),
.B(n_383),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_611),
.A2(n_430),
.B1(n_427),
.B2(n_417),
.Y(n_718)
);

AO21x2_ASAP7_75t_L g719 ( 
.A1(n_642),
.A2(n_406),
.B(n_383),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_657),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_602),
.A2(n_430),
.B1(n_427),
.B2(n_417),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_602),
.A2(n_417),
.B1(n_406),
.B2(n_383),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_579),
.Y(n_723)
);

OAI221xp5_ASAP7_75t_L g724 ( 
.A1(n_592),
.A2(n_406),
.B1(n_383),
.B2(n_372),
.C(n_355),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_588),
.A2(n_372),
.B1(n_355),
.B2(n_340),
.Y(n_725)
);

CKINVDCx11_ASAP7_75t_R g726 ( 
.A(n_557),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_581),
.Y(n_727)
);

AO31x2_ASAP7_75t_L g728 ( 
.A1(n_631),
.A2(n_372),
.A3(n_355),
.B(n_340),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_556),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_556),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_556),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_649),
.B(n_33),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_612),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_566),
.B(n_39),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_562),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_585),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_736)
);

BUFx8_ASAP7_75t_L g737 ( 
.A(n_645),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_610),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_562),
.B(n_372),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_580),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_580),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_557),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_613),
.Y(n_743)
);

NAND2x1p5_ASAP7_75t_L g744 ( 
.A(n_616),
.B(n_355),
.Y(n_744)
);

OAI211xp5_ASAP7_75t_L g745 ( 
.A1(n_584),
.A2(n_340),
.B(n_337),
.C(n_59),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_580),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_628),
.A2(n_340),
.B1(n_337),
.B2(n_60),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_596),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_628),
.A2(n_337),
.B1(n_55),
.B2(n_63),
.Y(n_749)
);

INVx3_ASAP7_75t_SL g750 ( 
.A(n_583),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_554),
.A2(n_337),
.B(n_64),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_583),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_567),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_596),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_590),
.A2(n_629),
.B1(n_554),
.B2(n_643),
.Y(n_755)
);

BUFx4f_ASAP7_75t_SL g756 ( 
.A(n_648),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_626),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_618),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_578),
.A2(n_47),
.B(n_65),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_614),
.Y(n_760)
);

OAI221xp5_ASAP7_75t_L g761 ( 
.A1(n_625),
.A2(n_70),
.B1(n_71),
.B2(n_76),
.C(n_77),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_566),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_634),
.B(n_79),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_623),
.B(n_80),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_643),
.A2(n_81),
.B1(n_83),
.B2(n_87),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_596),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_561),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_561),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_SL g769 ( 
.A1(n_626),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_569),
.B(n_143),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_654),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_599),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_616),
.B(n_110),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_661),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_569),
.B(n_140),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_628),
.B(n_112),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_647),
.Y(n_777)
);

BUFx4f_ASAP7_75t_SL g778 ( 
.A(n_594),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_594),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_599),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_610),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_599),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_619),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_660),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_646),
.B(n_124),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_627),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_679),
.Y(n_787)
);

OA21x2_ASAP7_75t_L g788 ( 
.A1(n_745),
.A2(n_620),
.B(n_582),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_666),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_SL g790 ( 
.A1(n_697),
.A2(n_601),
.B1(n_644),
.B2(n_630),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_SL g791 ( 
.A1(n_697),
.A2(n_601),
.B1(n_644),
.B2(n_630),
.Y(n_791)
);

OAI21xp33_ASAP7_75t_SL g792 ( 
.A1(n_732),
.A2(n_601),
.B(n_608),
.Y(n_792)
);

AO21x2_ASAP7_75t_L g793 ( 
.A1(n_724),
.A2(n_558),
.B(n_559),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_673),
.Y(n_794)
);

AOI221xp5_ASAP7_75t_L g795 ( 
.A1(n_743),
.A2(n_662),
.B1(n_633),
.B2(n_572),
.C(n_571),
.Y(n_795)
);

AOI21xp33_ASAP7_75t_L g796 ( 
.A1(n_668),
.A2(n_560),
.B(n_568),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_751),
.A2(n_593),
.B(n_575),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_682),
.B(n_593),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_666),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_SL g800 ( 
.A1(n_697),
.A2(n_734),
.B1(n_716),
.B2(n_778),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_669),
.A2(n_575),
.B1(n_636),
.B2(n_615),
.Y(n_801)
);

OAI21x1_ASAP7_75t_L g802 ( 
.A1(n_751),
.A2(n_603),
.B(n_636),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_779),
.A2(n_603),
.B1(n_636),
.B2(n_615),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_672),
.Y(n_804)
);

OAI22xp33_ASAP7_75t_L g805 ( 
.A1(n_665),
.A2(n_603),
.B1(n_615),
.B2(n_651),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_715),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_667),
.B(n_663),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_669),
.A2(n_132),
.B1(n_134),
.B2(n_138),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_676),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_674),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_734),
.B(n_139),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_695),
.A2(n_671),
.B1(n_674),
.B2(n_755),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_724),
.A2(n_721),
.B1(n_747),
.B2(n_675),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_716),
.B(n_770),
.Y(n_814)
);

OA21x2_ASAP7_75t_L g815 ( 
.A1(n_745),
.A2(n_759),
.B(n_722),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_SL g816 ( 
.A1(n_778),
.A2(n_770),
.B1(n_775),
.B2(n_761),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_757),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_755),
.A2(n_663),
.B1(n_688),
.B2(n_680),
.Y(n_818)
);

OAI221xp5_ASAP7_75t_L g819 ( 
.A1(n_762),
.A2(n_675),
.B1(n_752),
.B2(n_694),
.C(n_708),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_684),
.Y(n_820)
);

AOI221xp5_ASAP7_75t_L g821 ( 
.A1(n_686),
.A2(n_709),
.B1(n_677),
.B2(n_696),
.C(n_702),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_775),
.B(n_689),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_685),
.B(n_750),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_693),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_688),
.A2(n_687),
.B1(n_670),
.B2(n_735),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_687),
.A2(n_760),
.B1(n_763),
.B2(n_750),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_721),
.A2(n_747),
.B1(n_749),
.B2(n_700),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_785),
.A2(n_776),
.B1(n_707),
.B2(n_692),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_705),
.A2(n_742),
.B1(n_733),
.B2(n_758),
.Y(n_829)
);

CKINVDCx11_ASAP7_75t_R g830 ( 
.A(n_726),
.Y(n_830)
);

BUFx12f_ASAP7_75t_L g831 ( 
.A(n_737),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_698),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_771),
.B(n_774),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_707),
.A2(n_692),
.B1(n_710),
.B2(n_706),
.Y(n_834)
);

AOI222xp33_ASAP7_75t_L g835 ( 
.A1(n_701),
.A2(n_711),
.B1(n_756),
.B2(n_737),
.C1(n_761),
.C2(n_753),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_700),
.A2(n_699),
.B1(n_714),
.B2(n_739),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_756),
.B(n_683),
.Y(n_837)
);

OAI22xp33_ASAP7_75t_L g838 ( 
.A1(n_764),
.A2(n_739),
.B1(n_749),
.B2(n_664),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_699),
.A2(n_739),
.B1(n_732),
.B2(n_769),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_777),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_769),
.A2(n_765),
.B1(n_704),
.B2(n_767),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_664),
.A2(n_720),
.B1(n_666),
.B2(n_727),
.Y(n_842)
);

OR2x6_ASAP7_75t_L g843 ( 
.A(n_720),
.B(n_723),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_784),
.A2(n_738),
.B1(n_781),
.B2(n_691),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_765),
.A2(n_704),
.B1(n_767),
.B2(n_768),
.Y(n_845)
);

OAI22xp33_ASAP7_75t_L g846 ( 
.A1(n_783),
.A2(n_738),
.B1(n_781),
.B2(n_703),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_713),
.A2(n_718),
.B1(n_690),
.B2(n_773),
.Y(n_847)
);

AOI21xp33_ASAP7_75t_L g848 ( 
.A1(n_736),
.A2(n_719),
.B(n_768),
.Y(n_848)
);

OAI21xp33_ASAP7_75t_SL g849 ( 
.A1(n_786),
.A2(n_725),
.B(n_782),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_681),
.B(n_740),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_717),
.B(n_741),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_786),
.A2(n_731),
.B1(n_772),
.B2(n_766),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_SL g853 ( 
.A1(n_744),
.A2(n_729),
.B1(n_754),
.B2(n_748),
.Y(n_853)
);

OAI211xp5_ASAP7_75t_L g854 ( 
.A1(n_725),
.A2(n_780),
.B(n_746),
.C(n_730),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_678),
.A2(n_712),
.B1(n_717),
.B2(n_728),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_719),
.A2(n_678),
.B1(n_717),
.B2(n_728),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_717),
.Y(n_857)
);

AOI221xp5_ASAP7_75t_L g858 ( 
.A1(n_678),
.A2(n_673),
.B1(n_524),
.B2(n_622),
.C(n_635),
.Y(n_858)
);

AND2x4_ASAP7_75t_SL g859 ( 
.A(n_728),
.B(n_705),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_728),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_671),
.A2(n_570),
.B1(n_564),
.B2(n_563),
.Y(n_861)
);

NAND2x1p5_ASAP7_75t_L g862 ( 
.A(n_716),
.B(n_664),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_682),
.B(n_564),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_673),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_679),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_673),
.B(n_524),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_673),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_804),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_835),
.A2(n_816),
.B1(n_861),
.B2(n_826),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_809),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_L g871 ( 
.A(n_835),
.B(n_791),
.C(n_790),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_859),
.B(n_814),
.Y(n_872)
);

OAI211xp5_ASAP7_75t_L g873 ( 
.A1(n_800),
.A2(n_812),
.B(n_818),
.C(n_858),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_SL g874 ( 
.A1(n_861),
.A2(n_839),
.B1(n_811),
.B2(n_814),
.Y(n_874)
);

OAI211xp5_ASAP7_75t_L g875 ( 
.A1(n_819),
.A2(n_829),
.B(n_842),
.C(n_821),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_L g876 ( 
.A(n_856),
.B(n_855),
.C(n_860),
.Y(n_876)
);

BUFx2_ASAP7_75t_SL g877 ( 
.A(n_811),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_807),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_820),
.B(n_824),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_807),
.B(n_863),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_857),
.Y(n_881)
);

OAI221xp5_ASAP7_75t_L g882 ( 
.A1(n_825),
.A2(n_828),
.B1(n_839),
.B2(n_863),
.C(n_795),
.Y(n_882)
);

NAND4xp25_ASAP7_75t_SL g883 ( 
.A(n_830),
.B(n_823),
.C(n_801),
.D(n_866),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_SL g884 ( 
.A1(n_827),
.A2(n_813),
.B1(n_822),
.B2(n_841),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_806),
.Y(n_885)
);

BUFx4f_ASAP7_75t_SL g886 ( 
.A(n_831),
.Y(n_886)
);

AO21x2_ASAP7_75t_L g887 ( 
.A1(n_855),
.A2(n_848),
.B(n_813),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_794),
.B(n_864),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_SL g889 ( 
.A1(n_827),
.A2(n_822),
.B1(n_841),
.B2(n_845),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_838),
.A2(n_845),
.B1(n_810),
.B2(n_867),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_843),
.B(n_840),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_851),
.Y(n_892)
);

AOI221xp5_ASAP7_75t_L g893 ( 
.A1(n_796),
.A2(n_798),
.B1(n_848),
.B2(n_817),
.C(n_834),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_836),
.A2(n_844),
.B1(n_843),
.B2(n_846),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_SL g895 ( 
.A1(n_862),
.A2(n_792),
.B1(n_815),
.B2(n_849),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_862),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_843),
.A2(n_808),
.B1(n_852),
.B2(n_803),
.Y(n_897)
);

OAI33xp33_ASAP7_75t_L g898 ( 
.A1(n_805),
.A2(n_832),
.A3(n_796),
.B1(n_798),
.B2(n_850),
.B3(n_799),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_802),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_833),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_797),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_789),
.B(n_799),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_SL g903 ( 
.A1(n_815),
.A2(n_854),
.B1(n_789),
.B2(n_799),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_793),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_789),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_793),
.Y(n_906)
);

OAI33xp33_ASAP7_75t_L g907 ( 
.A1(n_837),
.A2(n_847),
.A3(n_787),
.B1(n_865),
.B2(n_853),
.B3(n_788),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_788),
.Y(n_908)
);

OAI33xp33_ASAP7_75t_L g909 ( 
.A1(n_810),
.A2(n_529),
.A3(n_794),
.B1(n_864),
.B2(n_867),
.B3(n_861),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_859),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_892),
.B(n_889),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_892),
.B(n_884),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_885),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_L g914 ( 
.A(n_875),
.B(n_871),
.C(n_883),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_877),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_880),
.B(n_878),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_900),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_878),
.B(n_880),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_890),
.B(n_868),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_908),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_910),
.B(n_881),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_881),
.Y(n_922)
);

OAI33xp33_ASAP7_75t_L g923 ( 
.A1(n_888),
.A2(n_868),
.A3(n_871),
.B1(n_894),
.B2(n_904),
.B3(n_891),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_870),
.B(n_879),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_870),
.B(n_879),
.Y(n_925)
);

INVxp67_ASAP7_75t_SL g926 ( 
.A(n_910),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_901),
.A2(n_899),
.B(n_874),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_887),
.B(n_904),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_877),
.B(n_900),
.Y(n_929)
);

AOI211xp5_ASAP7_75t_L g930 ( 
.A1(n_873),
.A2(n_882),
.B(n_894),
.C(n_896),
.Y(n_930)
);

OAI33xp33_ASAP7_75t_L g931 ( 
.A1(n_888),
.A2(n_891),
.A3(n_876),
.B1(n_897),
.B2(n_906),
.B3(n_909),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_922),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_914),
.A2(n_869),
.B1(n_911),
.B2(n_912),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_921),
.B(n_876),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_924),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_913),
.B(n_886),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_917),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_924),
.B(n_925),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_920),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_921),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_929),
.B(n_927),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_SL g942 ( 
.A1(n_915),
.A2(n_872),
.B1(n_897),
.B2(n_887),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_925),
.B(n_872),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_912),
.B(n_872),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_935),
.B(n_928),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_932),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_937),
.B(n_911),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_938),
.B(n_919),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_940),
.B(n_932),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_939),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_933),
.B(n_919),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_936),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_944),
.B(n_918),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_942),
.A2(n_930),
.B(n_915),
.Y(n_954)
);

AND3x2_ASAP7_75t_L g955 ( 
.A(n_940),
.B(n_930),
.C(n_926),
.Y(n_955)
);

AND4x1_ASAP7_75t_L g956 ( 
.A(n_943),
.B(n_923),
.C(n_893),
.D(n_931),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_939),
.B(n_916),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_945),
.B(n_957),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_945),
.B(n_928),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_947),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_946),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_951),
.B(n_918),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_949),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_949),
.Y(n_964)
);

NAND2x1_ASAP7_75t_L g965 ( 
.A(n_954),
.B(n_941),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_950),
.B(n_934),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_950),
.B(n_934),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_948),
.B(n_916),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_957),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_958),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_963),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_960),
.B(n_934),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_965),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_964),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_SL g975 ( 
.A(n_968),
.B(n_929),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_960),
.B(n_962),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_961),
.Y(n_977)
);

XOR2x2_ASAP7_75t_L g978 ( 
.A(n_969),
.B(n_952),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_959),
.B(n_956),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_966),
.B(n_953),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_979),
.A2(n_967),
.B1(n_966),
.B2(n_955),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_977),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_980),
.B(n_967),
.Y(n_983)
);

BUFx4f_ASAP7_75t_SL g984 ( 
.A(n_973),
.Y(n_984)
);

NAND5xp2_ASAP7_75t_L g985 ( 
.A(n_981),
.B(n_895),
.C(n_927),
.D(n_903),
.E(n_976),
.Y(n_985)
);

NAND4xp25_ASAP7_75t_SL g986 ( 
.A(n_984),
.B(n_978),
.C(n_970),
.D(n_973),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_SL g987 ( 
.A1(n_984),
.A2(n_973),
.B1(n_978),
.B2(n_872),
.Y(n_987)
);

NAND4xp25_ASAP7_75t_L g988 ( 
.A(n_985),
.B(n_975),
.C(n_972),
.D(n_982),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_986),
.B(n_974),
.Y(n_989)
);

OR3x1_ASAP7_75t_L g990 ( 
.A(n_988),
.B(n_987),
.C(n_931),
.Y(n_990)
);

NOR4xp25_ASAP7_75t_L g991 ( 
.A(n_989),
.B(n_971),
.C(n_972),
.D(n_983),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_990),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_L g993 ( 
.A(n_991),
.B(n_975),
.C(n_907),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_992),
.A2(n_941),
.B1(n_898),
.B2(n_921),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_993),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_995),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_996),
.Y(n_997)
);

AOI221xp5_ASAP7_75t_L g998 ( 
.A1(n_997),
.A2(n_994),
.B1(n_905),
.B2(n_902),
.C(n_921),
.Y(n_998)
);


endmodule