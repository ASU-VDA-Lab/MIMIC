module fake_jpeg_879_n_93 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx12_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_25),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_26),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_32),
.B1(n_27),
.B2(n_24),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_23),
.B(n_2),
.C(n_3),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_0),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_29),
.B1(n_27),
.B2(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_40),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_7),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_57),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_64),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_53),
.A3(n_57),
.B1(n_4),
.B2(n_5),
.Y(n_63)
);

AO21x1_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_65),
.B(n_8),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_70),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_42),
.B1(n_11),
.B2(n_12),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_73),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_9),
.C(n_13),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_14),
.C(n_16),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_77),
.B1(n_73),
.B2(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_87),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_85),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_80),
.B(n_79),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_82),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_82),
.Y(n_93)
);


endmodule