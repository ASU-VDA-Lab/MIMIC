module fake_netlist_1_10834_n_663 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_663);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_663;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_476;
wire n_617;
wire n_227;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx4_ASAP7_75t_R g77 ( .A(n_53), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_10), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_63), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_29), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_9), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_17), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_38), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_39), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_52), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_30), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_18), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_31), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_21), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_9), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_75), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_61), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_76), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_16), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_34), .Y(n_95) );
BUFx3_ASAP7_75t_L g96 ( .A(n_44), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_1), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_45), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_43), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_55), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_72), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_35), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_48), .Y(n_103) );
INVxp33_ASAP7_75t_SL g104 ( .A(n_19), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_71), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_15), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_54), .Y(n_108) );
INVxp33_ASAP7_75t_L g109 ( .A(n_23), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_28), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_47), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_50), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_16), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_41), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_3), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_7), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_73), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_67), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_58), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_79), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_82), .B(n_0), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_93), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_79), .Y(n_123) );
BUFx12f_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_82), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_104), .B(n_0), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_97), .B(n_1), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g129 ( .A(n_115), .B(n_2), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_119), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_93), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_109), .B(n_3), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_83), .B(n_4), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_99), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_87), .B(n_4), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_84), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_94), .B(n_5), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_96), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_94), .B(n_5), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_96), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_88), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_107), .B(n_6), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_89), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_107), .B(n_6), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_99), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_95), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_95), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_102), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_91), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_116), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_102), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_103), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_100), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_149), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_125), .B(n_78), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g160 ( .A1(n_132), .A2(n_81), .B1(n_106), .B2(n_113), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_139), .B(n_113), .Y(n_161) );
INVx5_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
BUFx3_ASAP7_75t_L g163 ( .A(n_140), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_149), .Y(n_164) );
AND2x6_ASAP7_75t_L g165 ( .A(n_139), .B(n_118), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_125), .B(n_118), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_133), .B(n_103), .Y(n_167) );
OR2x6_ASAP7_75t_L g168 ( .A(n_127), .B(n_111), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_133), .B(n_105), .Y(n_169) );
INVx1_ASAP7_75t_SL g170 ( .A(n_127), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_149), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_132), .B(n_92), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
OR2x2_ASAP7_75t_L g175 ( .A(n_132), .B(n_90), .Y(n_175) );
INVx5_ASAP7_75t_L g176 ( .A(n_140), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_120), .B(n_110), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_155), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
NAND2xp33_ASAP7_75t_SL g182 ( .A(n_137), .B(n_117), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_120), .B(n_114), .Y(n_183) );
AND2x6_ASAP7_75t_L g184 ( .A(n_139), .B(n_111), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_137), .B(n_108), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_137), .B(n_108), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_148), .B(n_105), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_148), .A2(n_85), .B1(n_101), .B2(n_98), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_148), .Y(n_190) );
OR2x6_ASAP7_75t_L g191 ( .A(n_129), .B(n_77), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_123), .B(n_112), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_123), .B(n_86), .Y(n_194) );
INVx6_ASAP7_75t_L g195 ( .A(n_140), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_155), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_154), .Y(n_197) );
INVxp33_ASAP7_75t_L g198 ( .A(n_126), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_140), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_146), .B(n_147), .Y(n_200) );
INVxp67_ASAP7_75t_L g201 ( .A(n_130), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_146), .B(n_7), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_140), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_155), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_200), .B(n_144), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_200), .B(n_144), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_163), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_185), .B(n_146), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_165), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_173), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_181), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_159), .B(n_150), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_173), .Y(n_213) );
O2A1O1Ixp5_ASAP7_75t_L g214 ( .A1(n_194), .A2(n_148), .B(n_142), .C(n_138), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_185), .B(n_150), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_186), .B(n_151), .Y(n_216) );
INVx5_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_180), .Y(n_218) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_170), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_186), .B(n_128), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_181), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_163), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_168), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_165), .A2(n_128), .B1(n_156), .B2(n_138), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_172), .B(n_156), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_180), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_190), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_190), .A2(n_142), .B(n_135), .C(n_145), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_192), .B(n_135), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_196), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_189), .B(n_124), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_168), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_165), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_190), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_161), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_198), .B(n_124), .Y(n_237) );
OR2x6_ASAP7_75t_L g238 ( .A(n_168), .B(n_121), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_161), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_175), .A2(n_121), .B(n_141), .C(n_151), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_197), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_161), .A2(n_145), .B(n_147), .Y(n_242) );
OAI22xp33_ASAP7_75t_L g243 ( .A1(n_168), .A2(n_157), .B1(n_153), .B2(n_141), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_196), .Y(n_244) );
INVx4_ASAP7_75t_L g245 ( .A(n_165), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_178), .A2(n_142), .B(n_122), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_183), .B(n_142), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_199), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_166), .B(n_124), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_202), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_202), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_204), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_167), .B(n_134), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_165), .B(n_152), .Y(n_254) );
NAND3xp33_ASAP7_75t_SL g255 ( .A(n_160), .B(n_152), .C(n_136), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_184), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_169), .A2(n_175), .B(n_193), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_184), .B(n_152), .Y(n_258) );
NOR3xp33_ASAP7_75t_SL g259 ( .A(n_182), .B(n_8), .C(n_10), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_184), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_184), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_211), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_219), .Y(n_263) );
INVx3_ASAP7_75t_SL g264 ( .A(n_241), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_223), .Y(n_265) );
NAND3xp33_ASAP7_75t_L g266 ( .A(n_259), .B(n_143), .C(n_176), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_245), .B(n_182), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_240), .A2(n_191), .B(n_201), .C(n_131), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_238), .A2(n_122), .B1(n_136), .B2(n_131), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_208), .B(n_191), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_212), .A2(n_174), .B(n_171), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_122), .B(n_131), .C(n_136), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_238), .A2(n_191), .B1(n_184), .B2(n_188), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_245), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_208), .B(n_188), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_241), .Y(n_276) );
AO32x1_ASAP7_75t_L g277 ( .A1(n_250), .A2(n_204), .A3(n_158), .B1(n_164), .B2(n_171), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_220), .Y(n_278) );
BUFx12f_ASAP7_75t_L g279 ( .A(n_223), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_211), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_238), .A2(n_184), .B1(n_188), .B2(n_191), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_245), .Y(n_282) );
NAND2x1p5_ASAP7_75t_L g283 ( .A(n_217), .B(n_203), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_220), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_236), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_238), .A2(n_188), .B1(n_143), .B2(n_195), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_209), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_233), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_217), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_215), .B(n_188), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_216), .B(n_188), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_225), .A2(n_158), .B(n_193), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_221), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_236), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_250), .A2(n_143), .B1(n_199), .B2(n_203), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_237), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_209), .B(n_197), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_205), .B(n_143), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_206), .B(n_143), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_221), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_239), .A2(n_143), .B1(n_195), .B2(n_162), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_251), .Y(n_302) );
INVx4_ASAP7_75t_L g303 ( .A(n_217), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_247), .A2(n_164), .B(n_187), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_251), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g306 ( .A1(n_257), .A2(n_187), .B(n_174), .C(n_176), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_254), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_254), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_254), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_230), .A2(n_179), .B(n_177), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_226), .A2(n_179), .B(n_177), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_226), .A2(n_179), .B(n_177), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_263), .Y(n_313) );
NAND2x1p5_ASAP7_75t_L g314 ( .A(n_274), .B(n_217), .Y(n_314) );
BUFx12f_ASAP7_75t_L g315 ( .A(n_279), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_262), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_270), .B(n_217), .Y(n_317) );
AO31x2_ASAP7_75t_L g318 ( .A1(n_269), .A2(n_229), .A3(n_246), .B(n_253), .Y(n_318) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_297), .A2(n_243), .B1(n_249), .B2(n_239), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
BUFx4f_ASAP7_75t_L g321 ( .A(n_274), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_280), .Y(n_322) );
OAI21xp5_ASAP7_75t_L g323 ( .A1(n_290), .A2(n_235), .B(n_228), .Y(n_323) );
AO21x2_ASAP7_75t_L g324 ( .A1(n_310), .A2(n_255), .B(n_258), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_293), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_278), .B(n_232), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_268), .A2(n_214), .B(n_228), .C(n_235), .Y(n_327) );
INVx5_ASAP7_75t_L g328 ( .A(n_274), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_270), .B(n_234), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_281), .A2(n_224), .B1(n_234), .B2(n_258), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_294), .Y(n_331) );
OAI21x1_ASAP7_75t_L g332 ( .A1(n_311), .A2(n_312), .B(n_269), .Y(n_332) );
NOR2xp67_ASAP7_75t_L g333 ( .A(n_281), .B(n_261), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_295), .A2(n_292), .B(n_271), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_284), .B(n_261), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_265), .B(n_256), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_265), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_300), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_295), .A2(n_256), .B(n_260), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_297), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g341 ( .A1(n_291), .A2(n_213), .B(n_210), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_286), .A2(n_195), .B1(n_248), .B2(n_207), .Y(n_342) );
O2A1O1Ixp33_ASAP7_75t_L g343 ( .A1(n_275), .A2(n_252), .B(n_244), .C(n_231), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_302), .B(n_207), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_304), .A2(n_252), .B(n_210), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_319), .A2(n_276), .B1(n_296), .B2(n_273), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_315), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_340), .A2(n_305), .B1(n_266), .B2(n_297), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_327), .A2(n_306), .B(n_273), .Y(n_349) );
OAI22xp5_ASAP7_75t_SL g350 ( .A1(n_315), .A2(n_264), .B1(n_288), .B2(n_266), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_338), .A2(n_286), .B1(n_299), .B2(n_309), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_315), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_337), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_342), .A2(n_277), .B(n_298), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_338), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_313), .B(n_307), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_320), .A2(n_267), .B1(n_272), .B2(n_308), .C(n_301), .Y(n_357) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_326), .A2(n_299), .B(n_244), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_326), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_320), .B(n_299), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_316), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_316), .A2(n_282), .B1(n_287), .B2(n_283), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_331), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_330), .A2(n_282), .B1(n_287), .B2(n_289), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_330), .A2(n_282), .B1(n_287), .B2(n_289), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_329), .B(n_303), .Y(n_366) );
OAI322xp33_ASAP7_75t_L g367 ( .A1(n_331), .A2(n_177), .A3(n_179), .B1(n_12), .B2(n_13), .C1(n_14), .C2(n_15), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_321), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_334), .A2(n_283), .B(n_213), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_316), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_332), .A2(n_277), .B(n_218), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_329), .B(n_303), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_370), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_361), .B(n_318), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_346), .A2(n_333), .B1(n_329), .B2(n_336), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_361), .B(n_333), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_371), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_355), .B(n_322), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_369), .B(n_328), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_363), .B(n_322), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_360), .B(n_322), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_365), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_359), .B(n_325), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_366), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_353), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_367), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_364), .B(n_325), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_366), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_358), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_366), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_351), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_368), .Y(n_392) );
BUFx2_ASAP7_75t_L g393 ( .A(n_368), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_362), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_372), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_349), .B(n_325), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_372), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_354), .Y(n_398) );
INVx2_ASAP7_75t_SL g399 ( .A(n_356), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_357), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_348), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_348), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_350), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_386), .A2(n_352), .B1(n_335), .B2(n_342), .C(n_323), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_384), .Y(n_405) );
NAND2x1_ASAP7_75t_L g406 ( .A(n_379), .B(n_344), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_381), .B(n_318), .Y(n_407) );
AO21x2_ASAP7_75t_L g408 ( .A1(n_398), .A2(n_332), .B(n_334), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_374), .B(n_318), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_381), .B(n_378), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_374), .B(n_318), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_374), .B(n_318), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_403), .B(n_347), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g414 ( .A1(n_386), .A2(n_335), .B1(n_344), .B2(n_343), .C(n_347), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_377), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_381), .B(n_318), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_377), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_378), .B(n_324), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_399), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_378), .B(n_324), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_399), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_401), .B(n_324), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_379), .B(n_324), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_379), .Y(n_424) );
AO21x2_ASAP7_75t_L g425 ( .A1(n_398), .A2(n_345), .B(n_339), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_401), .B(n_8), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_393), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_379), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g429 ( .A1(n_403), .A2(n_321), .B(n_317), .C(n_336), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_373), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_380), .B(n_328), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_373), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_396), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_399), .B(n_317), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_377), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_383), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_380), .B(n_402), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_383), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_402), .B(n_336), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_396), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_379), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_380), .B(n_336), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g443 ( .A1(n_400), .A2(n_375), .B1(n_385), .B2(n_395), .C(n_397), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_396), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_384), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_383), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_376), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_409), .B(n_391), .Y(n_448) );
NAND2x1p5_ASAP7_75t_L g449 ( .A(n_406), .B(n_384), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_407), .B(n_391), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_419), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_443), .A2(n_400), .B1(n_397), .B2(n_395), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_421), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_407), .B(n_391), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_430), .Y(n_455) );
NOR3xp33_ASAP7_75t_L g456 ( .A(n_413), .B(n_385), .C(n_392), .Y(n_456) );
NAND2x1p5_ASAP7_75t_L g457 ( .A(n_406), .B(n_384), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_430), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_431), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_432), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_416), .B(n_387), .Y(n_461) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_431), .B(n_384), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_432), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_436), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_409), .B(n_382), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_416), .B(n_410), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_411), .B(n_382), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_410), .B(n_387), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_411), .B(n_389), .Y(n_469) );
CKINVDCx8_ASAP7_75t_R g470 ( .A(n_445), .Y(n_470) );
NAND4xp75_ASAP7_75t_L g471 ( .A(n_434), .B(n_392), .C(n_388), .D(n_390), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_447), .B(n_387), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_415), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_433), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_418), .B(n_389), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_438), .Y(n_476) );
NAND2xp33_ASAP7_75t_SL g477 ( .A(n_427), .B(n_384), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_446), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_418), .B(n_376), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_415), .Y(n_480) );
BUFx3_ASAP7_75t_L g481 ( .A(n_445), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_437), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_404), .B(n_384), .C(n_397), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_412), .B(n_395), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_415), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_412), .B(n_390), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_433), .B(n_390), .Y(n_487) );
NAND3xp33_ASAP7_75t_L g488 ( .A(n_404), .B(n_388), .C(n_394), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_437), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_420), .B(n_376), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_417), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_417), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_420), .B(n_376), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_426), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_426), .B(n_388), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_439), .B(n_376), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_442), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_440), .B(n_394), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_442), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_440), .B(n_394), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_440), .B(n_339), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_447), .B(n_392), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_439), .B(n_393), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_473), .Y(n_504) );
INVx3_ASAP7_75t_SL g505 ( .A(n_502), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_482), .B(n_444), .Y(n_506) );
CKINVDCx14_ASAP7_75t_R g507 ( .A(n_477), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_489), .B(n_444), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_455), .Y(n_509) );
NAND3xp33_ASAP7_75t_L g510 ( .A(n_456), .B(n_414), .C(n_443), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_451), .Y(n_511) );
NAND2x1_ASAP7_75t_L g512 ( .A(n_451), .B(n_424), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_494), .B(n_414), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_473), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_453), .B(n_429), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_466), .B(n_444), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_480), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_466), .B(n_422), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_480), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_459), .B(n_424), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_464), .B(n_422), .Y(n_522) );
OR2x6_ASAP7_75t_L g523 ( .A(n_449), .B(n_441), .Y(n_523) );
INVx4_ASAP7_75t_L g524 ( .A(n_449), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_468), .B(n_441), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_460), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_468), .B(n_428), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_479), .B(n_428), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_463), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_476), .B(n_405), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_478), .B(n_405), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_497), .B(n_408), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_SL g533 ( .A1(n_452), .A2(n_435), .B(n_417), .C(n_323), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_474), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_474), .Y(n_535) );
AND2x4_ASAP7_75t_SL g536 ( .A(n_502), .B(n_423), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_475), .B(n_423), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_485), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_475), .B(n_423), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_499), .B(n_408), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_461), .B(n_408), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_465), .B(n_423), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_465), .B(n_11), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_461), .B(n_408), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_467), .B(n_435), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_485), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_450), .B(n_435), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_487), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_467), .B(n_11), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_483), .B(n_488), .C(n_477), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_486), .B(n_425), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_486), .B(n_425), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_450), .B(n_425), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_491), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_479), .B(n_490), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_487), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_490), .B(n_425), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_484), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_509), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g560 ( .A1(n_510), .A2(n_471), .B(n_449), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_514), .A2(n_503), .B1(n_472), .B2(n_495), .C(n_493), .Y(n_561) );
AOI322xp5_ASAP7_75t_L g562 ( .A1(n_514), .A2(n_454), .A3(n_472), .B1(n_493), .B2(n_496), .C1(n_498), .C2(n_500), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_548), .B(n_469), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_513), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_526), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_517), .B(n_519), .Y(n_566) );
AOI211xp5_ASAP7_75t_L g567 ( .A1(n_543), .A2(n_502), .B(n_469), .C(n_484), .Y(n_567) );
OAI22xp5_ASAP7_75t_SL g568 ( .A1(n_507), .A2(n_470), .B1(n_457), .B2(n_462), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_516), .A2(n_472), .B1(n_471), .B2(n_454), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_533), .A2(n_457), .B(n_462), .C(n_448), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_516), .A2(n_448), .B1(n_462), .B2(n_481), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_556), .B(n_500), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_529), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_543), .A2(n_498), .B1(n_481), .B2(n_501), .Y(n_574) );
OAI22xp33_ASAP7_75t_SL g575 ( .A1(n_512), .A2(n_470), .B1(n_457), .B2(n_491), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_511), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_555), .B(n_12), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_534), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_533), .A2(n_492), .B(n_501), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_557), .A2(n_492), .B1(n_317), .B2(n_329), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_535), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_555), .B(n_13), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_558), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_549), .A2(n_177), .B1(n_179), .B2(n_317), .C(n_176), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_506), .Y(n_585) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_505), .A2(n_328), .B1(n_321), .B2(n_314), .Y(n_586) );
OAI321xp33_ASAP7_75t_L g587 ( .A1(n_550), .A2(n_341), .A3(n_314), .B1(n_18), .B2(n_19), .C(n_14), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_508), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_530), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g591 ( .A1(n_507), .A2(n_321), .B(n_328), .C(n_345), .Y(n_591) );
AO21x1_ASAP7_75t_L g592 ( .A1(n_524), .A2(n_17), .B(n_314), .Y(n_592) );
O2A1O1Ixp5_ASAP7_75t_L g593 ( .A1(n_524), .A2(n_341), .B(n_277), .C(n_328), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_522), .Y(n_594) );
NOR2x1p5_ASAP7_75t_L g595 ( .A(n_524), .B(n_20), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_525), .Y(n_596) );
INVx5_ASAP7_75t_L g597 ( .A(n_523), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_549), .A2(n_328), .B1(n_195), .B2(n_162), .Y(n_598) );
NAND4xp25_ASAP7_75t_L g599 ( .A(n_577), .B(n_541), .C(n_553), .D(n_540), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_575), .A2(n_523), .B(n_532), .Y(n_600) );
XNOR2xp5_ASAP7_75t_L g601 ( .A(n_582), .B(n_527), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g602 ( .A1(n_562), .A2(n_544), .B(n_537), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_566), .B(n_547), .Y(n_603) );
OAI322xp33_ASAP7_75t_L g604 ( .A1(n_594), .A2(n_590), .A3(n_589), .B1(n_574), .B2(n_563), .C1(n_588), .C2(n_585), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_596), .B(n_505), .Y(n_605) );
OAI21xp5_ASAP7_75t_SL g606 ( .A1(n_560), .A2(n_536), .B(n_521), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_559), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_572), .B(n_544), .Y(n_608) );
OAI21xp33_ASAP7_75t_L g609 ( .A1(n_571), .A2(n_537), .B(n_539), .Y(n_609) );
OAI211xp5_ASAP7_75t_L g610 ( .A1(n_567), .A2(n_552), .B(n_551), .C(n_539), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_561), .A2(n_528), .B1(n_542), .B2(n_536), .C(n_545), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_583), .B(n_554), .Y(n_612) );
NOR2x1_ASAP7_75t_L g613 ( .A(n_595), .B(n_523), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_569), .A2(n_554), .B1(n_546), .B2(n_538), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_576), .B(n_573), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_567), .A2(n_546), .B1(n_538), .B2(n_520), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_597), .A2(n_520), .B1(n_518), .B2(n_515), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g618 ( .A(n_587), .B(n_518), .C(n_515), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g619 ( .A1(n_591), .A2(n_504), .B(n_176), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_564), .B(n_504), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_565), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_578), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_581), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_611), .A2(n_592), .B1(n_568), .B2(n_598), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_606), .A2(n_570), .B1(n_584), .B2(n_580), .C(n_597), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_622), .Y(n_626) );
INVxp33_ASAP7_75t_SL g627 ( .A(n_613), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_623), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_605), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_604), .A2(n_579), .B1(n_586), .B2(n_593), .C(n_597), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_601), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g632 ( .A1(n_602), .A2(n_597), .B1(n_176), .B2(n_162), .C(n_26), .Y(n_632) );
NOR2xp67_ASAP7_75t_L g633 ( .A(n_610), .B(n_22), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_603), .Y(n_634) );
NAND4xp25_ASAP7_75t_L g635 ( .A(n_619), .B(n_24), .C(n_25), .D(n_27), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_600), .A2(n_162), .B(n_33), .Y(n_636) );
OAI321xp33_ASAP7_75t_L g637 ( .A1(n_599), .A2(n_32), .A3(n_36), .B1(n_37), .B2(n_40), .C(n_42), .Y(n_637) );
AOI31xp33_ASAP7_75t_L g638 ( .A1(n_609), .A2(n_46), .A3(n_49), .B(n_51), .Y(n_638) );
OAI211xp5_ASAP7_75t_SL g639 ( .A1(n_624), .A2(n_614), .B(n_621), .C(n_616), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_627), .A2(n_599), .B1(n_615), .B2(n_607), .C(n_618), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_626), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g642 ( .A1(n_625), .A2(n_617), .B(n_620), .C(n_612), .Y(n_642) );
AOI222xp33_ASAP7_75t_L g643 ( .A1(n_627), .A2(n_608), .B1(n_162), .B2(n_222), .C1(n_207), .C2(n_248), .Y(n_643) );
OAI211xp5_ASAP7_75t_SL g644 ( .A1(n_632), .A2(n_231), .B(n_227), .C(n_218), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_631), .A2(n_248), .B1(n_222), .B2(n_207), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_628), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_630), .A2(n_56), .B1(n_57), .B2(n_59), .C(n_60), .Y(n_647) );
NOR2x1_ASAP7_75t_L g648 ( .A(n_647), .B(n_635), .Y(n_648) );
NAND3xp33_ASAP7_75t_SL g649 ( .A(n_640), .B(n_636), .C(n_629), .Y(n_649) );
AND2x4_ASAP7_75t_L g650 ( .A(n_641), .B(n_634), .Y(n_650) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_639), .A2(n_633), .B1(n_638), .B2(n_637), .C(n_66), .Y(n_651) );
NOR3xp33_ASAP7_75t_L g652 ( .A(n_642), .B(n_227), .C(n_64), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g653 ( .A(n_648), .B(n_643), .C(n_645), .D(n_644), .Y(n_653) );
INVx3_ASAP7_75t_L g654 ( .A(n_650), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_649), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_654), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_655), .A2(n_652), .B1(n_651), .B2(n_646), .Y(n_657) );
OAI22xp5_ASAP7_75t_SL g658 ( .A1(n_657), .A2(n_653), .B1(n_65), .B2(n_68), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_656), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_659), .Y(n_660) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_660), .A2(n_658), .B1(n_69), .B2(n_70), .C1(n_74), .C2(n_62), .Y(n_661) );
AOI22x1_ASAP7_75t_L g662 ( .A1(n_661), .A2(n_207), .B1(n_222), .B2(n_248), .Y(n_662) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_662), .A2(n_222), .B1(n_248), .B2(n_655), .Y(n_663) );
endmodule