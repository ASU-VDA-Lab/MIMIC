module fake_jpeg_31080_n_288 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_225;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_154;
wire n_76;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_46),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_36),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_17),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_56),
.B(n_58),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_37),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_21),
.B1(n_28),
.B2(n_39),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_64),
.B1(n_86),
.B2(n_20),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_65),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_21),
.B1(n_28),
.B2(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_66),
.B(n_77),
.Y(n_94)
);

NAND2x1_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_46),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_27),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_75),
.Y(n_124)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_36),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_49),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_29),
.Y(n_101)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_44),
.B(n_23),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_35),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_32),
.B1(n_29),
.B2(n_39),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_92),
.B(n_101),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_57),
.A2(n_24),
.B(n_35),
.C(n_23),
.Y(n_95)
);

NOR2x1_ASAP7_75t_R g131 ( 
.A(n_95),
.B(n_90),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_116),
.B1(n_126),
.B2(n_74),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_99),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_33),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_113),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_33),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_28),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_123),
.C(n_82),
.Y(n_141)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_122),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_21),
.B1(n_31),
.B2(n_32),
.Y(n_116)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_56),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_30),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_77),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_78),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_129),
.B(n_136),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_130),
.A2(n_137),
.B1(n_99),
.B2(n_2),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_84),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_142),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_15),
.C(n_14),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_12),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_90),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_87),
.B1(n_88),
.B2(n_81),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_14),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_31),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_154),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_89),
.B1(n_59),
.B2(n_64),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_112),
.B1(n_98),
.B2(n_115),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_0),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_100),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_82),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_150),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_76),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_76),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_118),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_25),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_156),
.A2(n_95),
.B(n_108),
.C(n_104),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_157),
.A2(n_160),
.B1(n_181),
.B2(n_156),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_141),
.B1(n_155),
.B2(n_143),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_112),
.B1(n_109),
.B2(n_103),
.Y(n_160)
);

AO21x2_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_110),
.B(n_111),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_162),
.A2(n_182),
.B(n_186),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_121),
.B1(n_125),
.B2(n_108),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_104),
.C(n_123),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_174),
.C(n_155),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_93),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_172),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_123),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_173),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_125),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_147),
.C(n_145),
.Y(n_195)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_25),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_179),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_1),
.B(n_2),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_133),
.B(n_5),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_128),
.A2(n_5),
.B(n_6),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_148),
.B(n_9),
.Y(n_208)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_151),
.A2(n_7),
.B(n_8),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_189),
.A2(n_162),
.B(n_171),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_190),
.B(n_206),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_195),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_147),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_205),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_153),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_159),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_134),
.B(n_146),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_162),
.B(n_166),
.Y(n_211)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_210),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_217),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_173),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_228),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_207),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_162),
.B(n_161),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_219),
.B(n_220),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_197),
.B(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_167),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_224),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_202),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_194),
.B(n_168),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_191),
.B1(n_197),
.B2(n_196),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_200),
.B1(n_160),
.B2(n_210),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_227),
.A2(n_230),
.B1(n_187),
.B2(n_201),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_187),
.A2(n_157),
.B1(n_162),
.B2(n_167),
.Y(n_230)
);

INVx11_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_243),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_215),
.B1(n_229),
.B2(n_226),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_235),
.A2(n_238),
.B1(n_227),
.B2(n_211),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_216),
.B1(n_158),
.B2(n_186),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_209),
.B1(n_208),
.B2(n_198),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_214),
.A2(n_205),
.B1(n_204),
.B2(n_190),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_241),
.B1(n_231),
.B2(n_226),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_193),
.C(n_192),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_244),
.C(n_245),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_192),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_188),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_158),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_249),
.B1(n_252),
.B2(n_243),
.Y(n_259)
);

BUFx12_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_235),
.A2(n_223),
.B1(n_215),
.B2(n_219),
.Y(n_249)
);

A2O1A1O1Ixp25_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_221),
.B(n_212),
.C(n_229),
.D(n_220),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_256),
.B(n_254),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_193),
.C(n_222),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_254),
.C(n_234),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_222),
.C(n_188),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_257),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_253),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_127),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_263),
.B1(n_250),
.B2(n_249),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_234),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_262),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_216),
.Y(n_262)
);

AOI21x1_ASAP7_75t_SL g265 ( 
.A1(n_251),
.A2(n_238),
.B(n_245),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_248),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_250),
.Y(n_269)
);

NAND4xp25_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_248),
.C(n_238),
.D(n_247),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_272),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_271),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_270),
.B(n_273),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_158),
.CI(n_127),
.CON(n_273),
.SN(n_273)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_266),
.C(n_258),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_269),
.B(n_144),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_264),
.B(n_146),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_277),
.B(n_273),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_276),
.B(n_264),
.Y(n_279)
);

OAI21x1_ASAP7_75t_L g284 ( 
.A1(n_279),
.A2(n_281),
.B(n_144),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g283 ( 
.A1(n_280),
.A2(n_282),
.B(n_278),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_270),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_283),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_284),
.C(n_9),
.Y(n_286)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_216),
.C1(n_285),
.C2(n_217),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_10),
.Y(n_288)
);


endmodule