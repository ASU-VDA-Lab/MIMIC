module fake_netlist_6_4936_n_2377 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2377);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2377;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2301;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_400;
wire n_739;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g233 ( 
.A(n_65),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_40),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_89),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_25),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_113),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_103),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_152),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_133),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_74),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_106),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_36),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_195),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_160),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_150),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_154),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_153),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_175),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_70),
.Y(n_252)
);

CKINVDCx11_ASAP7_75t_R g253 ( 
.A(n_120),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_223),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_38),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_164),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_97),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_177),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_30),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_40),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_156),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_207),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_155),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_9),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_108),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_109),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_99),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_134),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_55),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_101),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_22),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_137),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_216),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_118),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_56),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_11),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_123),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_102),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_112),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_15),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_219),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_14),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_6),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_222),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_227),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_200),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_47),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_183),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_173),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_34),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_14),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_111),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_147),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_171),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_52),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_17),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_101),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_36),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_6),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_192),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_64),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_31),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_108),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_226),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_76),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_208),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_104),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_38),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_107),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_189),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_131),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_165),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_196),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_64),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_187),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_70),
.Y(n_317)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_140),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_135),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_221),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_54),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_142),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_78),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_205),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_65),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_23),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_7),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_50),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_166),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_220),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_37),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_190),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_107),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_19),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_232),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_98),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_117),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_144),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_50),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_168),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_212),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_218),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_124),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_139),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_97),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_201),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_89),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_209),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_114),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_215),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_61),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_83),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_2),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_149),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_151),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_69),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_27),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_214),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_206),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_24),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_186),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_43),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_3),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_28),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_68),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_58),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_82),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_37),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_94),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_19),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_31),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_90),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_174),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_63),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_106),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_53),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_18),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_56),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_96),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_9),
.Y(n_380)
);

BUFx2_ASAP7_75t_SL g381 ( 
.A(n_197),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_43),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_51),
.Y(n_383)
);

BUFx2_ASAP7_75t_SL g384 ( 
.A(n_1),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_121),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_170),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_182),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_176),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_71),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_62),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_161),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_20),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_47),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_23),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_125),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_24),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_30),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_25),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_87),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_119),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_230),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_194),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_0),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_141),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_80),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_5),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_71),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_33),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_96),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_26),
.Y(n_410)
);

BUFx10_ASAP7_75t_L g411 ( 
.A(n_128),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_122),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_92),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_185),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_167),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_8),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_211),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_11),
.Y(n_418)
);

BUFx10_ASAP7_75t_L g419 ( 
.A(n_86),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_66),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_32),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_72),
.Y(n_422)
);

HB1xp67_ASAP7_75t_SL g423 ( 
.A(n_157),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_45),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_63),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_67),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_115),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_129),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_188),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_103),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_42),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_78),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_73),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_5),
.Y(n_434)
);

BUFx5_ASAP7_75t_L g435 ( 
.A(n_143),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_58),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_69),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_105),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_203),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_2),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_99),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_60),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_162),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_0),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_42),
.Y(n_445)
);

BUFx8_ASAP7_75t_SL g446 ( 
.A(n_172),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_109),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_83),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_180),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_94),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_159),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_132),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_181),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_92),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_136),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_57),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_274),
.B(n_1),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_446),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_280),
.Y(n_460)
);

INVxp33_ASAP7_75t_SL g461 ( 
.A(n_234),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_282),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_253),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_326),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_238),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_326),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_245),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_326),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_349),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_326),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_354),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_326),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_326),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_247),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_248),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_336),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_336),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_249),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_250),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_251),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_427),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_254),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_256),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_258),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_336),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_336),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_336),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_261),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_336),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_339),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_439),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_262),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_297),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_339),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_339),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_339),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_339),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_263),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_364),
.B(n_3),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_339),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_275),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_362),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_362),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_278),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_306),
.B(n_4),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_285),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_287),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_362),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_290),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_293),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_301),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_305),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_362),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_312),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_274),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_313),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_362),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_314),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_362),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_320),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_318),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_322),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_329),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_332),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_335),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_338),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_456),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_456),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_340),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_342),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_244),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_346),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_350),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_456),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_233),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_233),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_267),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_244),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_387),
.B(n_4),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_267),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_323),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_358),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_361),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_323),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_415),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_327),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_373),
.Y(n_548)
);

INVxp33_ASAP7_75t_SL g549 ( 
.A(n_235),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_327),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_388),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_390),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_364),
.B(n_7),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_400),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_387),
.B(n_8),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_390),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_243),
.B(n_10),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_325),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_415),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_402),
.Y(n_560)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_415),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_243),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_271),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_424),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_325),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_417),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_424),
.Y(n_567)
);

NOR2xp67_ASAP7_75t_L g568 ( 
.A(n_306),
.B(n_10),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_431),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_443),
.B(n_12),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_428),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_431),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_444),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_449),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_452),
.Y(n_575)
);

NOR2xp67_ASAP7_75t_L g576 ( 
.A(n_370),
.B(n_12),
.Y(n_576)
);

NOR2xp67_ASAP7_75t_L g577 ( 
.A(n_370),
.B(n_13),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_444),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_271),
.Y(n_579)
);

NOR2xp67_ASAP7_75t_L g580 ( 
.A(n_447),
.B(n_13),
.Y(n_580)
);

NAND2x1_ASAP7_75t_L g581 ( 
.A(n_465),
.B(n_443),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_466),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_465),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_460),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_468),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_467),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_467),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_558),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_546),
.B(n_561),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_469),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_559),
.B(n_455),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_469),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_494),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_471),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_475),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_471),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_473),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_473),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_462),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_565),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_476),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_464),
.B(n_436),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_474),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_470),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_500),
.B(n_240),
.Y(n_605)
);

INVxp33_ASAP7_75t_SL g606 ( 
.A(n_459),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_SL g607 ( 
.A(n_500),
.B(n_360),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_474),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_479),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_559),
.B(n_453),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_477),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_539),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_477),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_480),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_540),
.B(n_436),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_532),
.B(n_411),
.Y(n_616)
);

OA21x2_ASAP7_75t_L g617 ( 
.A1(n_478),
.A2(n_241),
.B(n_237),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_478),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_472),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_522),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_482),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_553),
.B(n_559),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_R g623 ( 
.A(n_505),
.B(n_423),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_486),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_492),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_539),
.B(n_321),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_553),
.B(n_364),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_486),
.B(n_426),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_487),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_487),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_488),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_570),
.B(n_307),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_488),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_490),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_490),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_491),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_555),
.B(n_412),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_522),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_532),
.B(n_411),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_491),
.B(n_426),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_481),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_483),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_511),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_522),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_495),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_495),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_484),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_485),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_496),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_489),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_R g651 ( 
.A(n_521),
.B(n_236),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_496),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_497),
.Y(n_653)
);

BUFx8_ASAP7_75t_L g654 ( 
.A(n_557),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_493),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_497),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_527),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_498),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_498),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_501),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_501),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_503),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_506),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_503),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_499),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_544),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_504),
.B(n_426),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_502),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_506),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_504),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_509),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_509),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_507),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_508),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_510),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_514),
.B(n_237),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_554),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_622),
.B(n_512),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_638),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_583),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_638),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_638),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_583),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_629),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_622),
.B(n_513),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_629),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_622),
.B(n_515),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_632),
.B(n_517),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_638),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_628),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_629),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_589),
.B(n_557),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_615),
.A2(n_516),
.B1(n_566),
.B2(n_560),
.Y(n_693)
);

AND2x6_ASAP7_75t_L g694 ( 
.A(n_605),
.B(n_295),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_587),
.Y(n_695)
);

CKINVDCx16_ASAP7_75t_R g696 ( 
.A(n_623),
.Y(n_696)
);

NAND2x1p5_ASAP7_75t_L g697 ( 
.A(n_617),
.B(n_241),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_583),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_638),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_587),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_SL g701 ( 
.A(n_626),
.B(n_458),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_627),
.B(n_528),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_627),
.B(n_528),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_638),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_596),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_637),
.B(n_461),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_638),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_596),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_632),
.B(n_519),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_612),
.B(n_457),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_598),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_637),
.B(n_549),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_589),
.B(n_523),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_598),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_627),
.B(n_529),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_586),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_615),
.B(n_524),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_591),
.B(n_525),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_644),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_651),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_591),
.B(n_526),
.Y(n_721)
);

INVx5_ASAP7_75t_L g722 ( 
.A(n_644),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_586),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_582),
.B(n_530),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_608),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_626),
.B(n_463),
.C(n_531),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_663),
.Y(n_727)
);

AO22x2_ASAP7_75t_L g728 ( 
.A1(n_616),
.A2(n_570),
.B1(n_284),
.B2(n_288),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_586),
.Y(n_729)
);

INVx6_ASAP7_75t_L g730 ( 
.A(n_605),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_610),
.B(n_533),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_610),
.B(n_534),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_605),
.B(n_543),
.Y(n_733)
);

AND2x6_ASAP7_75t_L g734 ( 
.A(n_605),
.B(n_295),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_590),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_628),
.B(n_529),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_585),
.B(n_548),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_644),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_590),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_590),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_595),
.B(n_551),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_644),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_628),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_608),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_663),
.B(n_571),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_624),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_643),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_676),
.B(n_640),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_644),
.Y(n_749)
);

AND2x6_ASAP7_75t_L g750 ( 
.A(n_676),
.B(n_295),
.Y(n_750)
);

AND2x6_ASAP7_75t_L g751 ( 
.A(n_676),
.B(n_295),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_669),
.B(n_574),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_624),
.Y(n_753)
);

INVx6_ASAP7_75t_L g754 ( 
.A(n_644),
.Y(n_754)
);

OR2x6_ASAP7_75t_L g755 ( 
.A(n_655),
.B(n_381),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_601),
.B(n_575),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_669),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_631),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_592),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_640),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_607),
.A2(n_576),
.B1(n_577),
.B2(n_568),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_592),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_667),
.B(n_535),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_581),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_581),
.Y(n_765)
);

AND2x2_ASAP7_75t_SL g766 ( 
.A(n_655),
.B(n_240),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_592),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_631),
.B(n_633),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_639),
.A2(n_580),
.B1(n_576),
.B2(n_577),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_588),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_667),
.B(n_535),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_644),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_594),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_633),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_588),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_609),
.B(n_568),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_584),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_634),
.B(n_514),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_634),
.B(n_518),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_635),
.B(n_649),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_654),
.Y(n_781)
);

BUFx4f_ASAP7_75t_L g782 ( 
.A(n_617),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_614),
.B(n_562),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_635),
.B(n_246),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_649),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_656),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_594),
.Y(n_787)
);

AND2x6_ASAP7_75t_L g788 ( 
.A(n_620),
.B(n_295),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_654),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_656),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_658),
.B(n_536),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_658),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_594),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_603),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_659),
.B(n_246),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_659),
.B(n_295),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_660),
.B(n_518),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_660),
.B(n_536),
.Y(n_798)
);

INVx5_ASAP7_75t_L g799 ( 
.A(n_652),
.Y(n_799)
);

AO22x2_ASAP7_75t_L g800 ( 
.A1(n_600),
.A2(n_284),
.B1(n_288),
.B2(n_272),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_661),
.B(n_264),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_661),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_620),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_603),
.Y(n_804)
);

INVx4_ASAP7_75t_SL g805 ( 
.A(n_652),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_657),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_662),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_599),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_597),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_662),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_671),
.B(n_672),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_671),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_597),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_620),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_597),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_672),
.B(n_520),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_641),
.B(n_411),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_642),
.B(n_411),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_611),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_604),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_620),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_602),
.B(n_381),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_611),
.B(n_264),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_647),
.B(n_563),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_603),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_603),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_611),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_603),
.B(n_520),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_603),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_648),
.B(n_579),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_652),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_613),
.B(n_269),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_613),
.B(n_269),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_618),
.Y(n_834)
);

INVxp33_ASAP7_75t_SL g835 ( 
.A(n_650),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_600),
.A2(n_580),
.B1(n_242),
.B2(n_252),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_618),
.B(n_273),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_665),
.B(n_321),
.Y(n_838)
);

BUFx6f_ASAP7_75t_SL g839 ( 
.A(n_766),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_713),
.B(n_668),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_695),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_760),
.B(n_673),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_706),
.B(n_674),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_695),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_718),
.B(n_675),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_712),
.A2(n_416),
.B1(n_433),
.B2(n_368),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_721),
.B(n_654),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_748),
.B(n_654),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_748),
.B(n_617),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_690),
.Y(n_850)
);

OR2x6_ASAP7_75t_L g851 ( 
.A(n_781),
.B(n_593),
.Y(n_851)
);

NOR2x2_ASAP7_75t_L g852 ( 
.A(n_822),
.B(n_330),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_763),
.B(n_617),
.Y(n_853)
);

OAI22xp33_ASAP7_75t_L g854 ( 
.A1(n_701),
.A2(n_769),
.B1(n_822),
.B2(n_709),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_748),
.A2(n_617),
.B1(n_355),
.B2(n_385),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_700),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_690),
.B(n_618),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_743),
.B(n_618),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_766),
.B(n_606),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_688),
.B(n_311),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_743),
.A2(n_355),
.B1(n_385),
.B2(n_330),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_727),
.B(n_311),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_731),
.B(n_618),
.Y(n_863)
);

NAND3xp33_ASAP7_75t_L g864 ( 
.A(n_761),
.B(n_255),
.C(n_239),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_700),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_732),
.B(n_618),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_705),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_763),
.B(n_537),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_730),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_705),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_728),
.A2(n_273),
.B1(n_289),
.B2(n_286),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_752),
.B(n_783),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_730),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_708),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_728),
.A2(n_289),
.B1(n_294),
.B2(n_286),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_728),
.A2(n_294),
.B1(n_319),
.B2(n_316),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_708),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_730),
.B(n_636),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_824),
.B(n_593),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_711),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_730),
.Y(n_881)
);

NOR2x2_ASAP7_75t_L g882 ( 
.A(n_822),
.B(n_321),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_710),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_814),
.B(n_636),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_684),
.B(n_636),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_686),
.B(n_636),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_711),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_728),
.A2(n_316),
.B1(n_324),
.B2(n_319),
.Y(n_888)
);

AND2x6_ASAP7_75t_SL g889 ( 
.A(n_822),
.B(n_272),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_714),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_727),
.B(n_311),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_757),
.B(n_311),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_714),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_L g894 ( 
.A(n_697),
.B(n_318),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_725),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_782),
.A2(n_630),
.B(n_613),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_702),
.B(n_537),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_764),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_715),
.A2(n_337),
.B1(n_341),
.B2(n_324),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_830),
.B(n_757),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_710),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_745),
.B(n_311),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_678),
.B(n_666),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_692),
.A2(n_337),
.B1(n_343),
.B2(n_341),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_725),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_775),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_691),
.B(n_636),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_744),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_733),
.B(n_311),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_774),
.B(n_636),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_692),
.A2(n_343),
.B1(n_348),
.B2(n_344),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_782),
.A2(n_687),
.B(n_685),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_774),
.B(n_652),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_744),
.Y(n_914)
);

INVx8_ASAP7_75t_L g915 ( 
.A(n_692),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_786),
.B(n_652),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_786),
.B(n_652),
.Y(n_917)
);

O2A1O1Ixp5_ASAP7_75t_L g918 ( 
.A1(n_782),
.A2(n_812),
.B(n_810),
.C(n_746),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_775),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_746),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_702),
.B(n_538),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_703),
.B(n_652),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_753),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_753),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_703),
.B(n_653),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_720),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_692),
.A2(n_348),
.B1(n_359),
.B2(n_344),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_758),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_771),
.B(n_653),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_758),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_771),
.B(n_715),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_785),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_771),
.B(n_653),
.Y(n_933)
);

OR2x6_ASAP7_75t_L g934 ( 
.A(n_781),
.B(n_359),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_715),
.B(n_736),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_736),
.B(n_538),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_693),
.B(n_391),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_694),
.A2(n_386),
.B1(n_401),
.B2(n_395),
.Y(n_938)
);

BUFx12f_ASAP7_75t_L g939 ( 
.A(n_777),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_785),
.B(n_790),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_790),
.B(n_653),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_792),
.B(n_653),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_770),
.Y(n_943)
);

NAND2xp33_ASAP7_75t_L g944 ( 
.A(n_697),
.B(n_318),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_792),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_802),
.B(n_653),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_717),
.B(n_391),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_800),
.A2(n_395),
.B1(n_401),
.B2(n_386),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_802),
.Y(n_949)
);

AO22x1_ASAP7_75t_L g950 ( 
.A1(n_784),
.A2(n_414),
.B1(n_404),
.B2(n_303),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_807),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_807),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_803),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_803),
.B(n_653),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_803),
.B(n_670),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_821),
.Y(n_956)
);

AND2x6_ASAP7_75t_SL g957 ( 
.A(n_755),
.B(n_298),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_821),
.B(n_670),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_821),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_768),
.B(n_670),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_724),
.B(n_677),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_800),
.A2(n_414),
.B1(n_404),
.B2(n_259),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_827),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_777),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_694),
.A2(n_391),
.B1(n_451),
.B2(n_429),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_784),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_680),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_827),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_784),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_737),
.B(n_619),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_741),
.B(n_621),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_756),
.B(n_625),
.Y(n_972)
);

NAND3xp33_ASAP7_75t_L g973 ( 
.A(n_726),
.B(n_260),
.C(n_257),
.Y(n_973)
);

OAI22xp33_ASAP7_75t_L g974 ( 
.A1(n_755),
.A2(n_303),
.B1(n_351),
.B2(n_298),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_755),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_764),
.B(n_351),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_780),
.B(n_670),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_791),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_828),
.A2(n_645),
.B(n_630),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_776),
.B(n_817),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_811),
.B(n_670),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_680),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_765),
.B(n_670),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_755),
.A2(n_391),
.B1(n_429),
.B2(n_451),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_754),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_683),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_791),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_765),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_679),
.B(n_670),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_818),
.B(n_265),
.Y(n_990)
);

OR2x6_ASAP7_75t_L g991 ( 
.A(n_789),
.B(n_356),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_694),
.A2(n_391),
.B1(n_429),
.B2(n_451),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_679),
.B(n_630),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_682),
.Y(n_994)
);

OAI22xp33_ASAP7_75t_L g995 ( 
.A1(n_836),
.A2(n_392),
.B1(n_356),
.B2(n_357),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_679),
.B(n_645),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_808),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_720),
.B(n_391),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_681),
.B(n_664),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_696),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_681),
.B(n_664),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_795),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_835),
.B(n_429),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_800),
.A2(n_291),
.B1(n_454),
.B2(n_450),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_835),
.B(n_429),
.Y(n_1005)
);

AOI221xp5_ASAP7_75t_L g1006 ( 
.A1(n_800),
.A2(n_357),
.B1(n_365),
.B2(n_372),
.C(n_377),
.Y(n_1006)
);

OAI221xp5_ASAP7_75t_L g1007 ( 
.A1(n_798),
.A2(n_365),
.B1(n_372),
.B2(n_442),
.C(n_437),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_683),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_795),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_789),
.B(n_429),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_698),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_926),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_872),
.B(n_795),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_841),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_898),
.B(n_801),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_873),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_R g1017 ( 
.A(n_1000),
.B(n_808),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_898),
.B(n_850),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_843),
.B(n_883),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_873),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_841),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_865),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_871),
.A2(n_694),
.B1(n_734),
.B2(n_801),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_865),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_906),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_867),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_SL g1027 ( 
.A1(n_839),
.A2(n_820),
.B1(n_806),
.B2(n_747),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_919),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_867),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_870),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_840),
.B(n_801),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_850),
.B(n_798),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_SL g1033 ( 
.A(n_995),
.B(n_820),
.C(n_268),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_988),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_900),
.B(n_697),
.Y(n_1035)
);

CKINVDCx16_ASAP7_75t_R g1036 ( 
.A(n_939),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_943),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_870),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_873),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_976),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_874),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_926),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_845),
.B(n_681),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_868),
.Y(n_1044)
);

AND3x1_ASAP7_75t_SL g1045 ( 
.A(n_1007),
.B(n_379),
.C(n_377),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_901),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_1000),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_874),
.Y(n_1048)
);

INVx5_ASAP7_75t_L g1049 ( 
.A(n_994),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_SL g1050 ( 
.A(n_974),
.B(n_270),
.C(n_266),
.Y(n_1050)
);

BUFx4_ASAP7_75t_SL g1051 ( 
.A(n_957),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_R g1052 ( 
.A(n_939),
.B(n_276),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_877),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_854),
.A2(n_838),
.B1(n_734),
.B2(n_694),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_877),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_988),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_918),
.A2(n_707),
.B(n_689),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_966),
.B(n_823),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_890),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_912),
.B(n_682),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_988),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_890),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_988),
.B(n_682),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_895),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_988),
.Y(n_1065)
);

INVx5_ASAP7_75t_L g1066 ( 
.A(n_994),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_994),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_895),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_905),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_915),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_868),
.B(n_844),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_966),
.B(n_823),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_937),
.A2(n_837),
.B(n_779),
.C(n_797),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_905),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_928),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_873),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_994),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_R g1078 ( 
.A(n_847),
.B(n_879),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_869),
.B(n_682),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_964),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_844),
.B(n_856),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_842),
.B(n_689),
.Y(n_1082)
);

AND2x6_ASAP7_75t_SL g1083 ( 
.A(n_961),
.B(n_379),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_856),
.B(n_880),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_969),
.B(n_823),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_928),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_976),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_880),
.B(n_689),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_930),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_997),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_975),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_930),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_869),
.B(n_682),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_887),
.B(n_707),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_932),
.Y(n_1095)
);

BUFx12f_ASAP7_75t_L g1096 ( 
.A(n_851),
.Y(n_1096)
);

AND2x6_ASAP7_75t_L g1097 ( 
.A(n_853),
.B(n_707),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_851),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_873),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_932),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_969),
.B(n_832),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_839),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_887),
.B(n_699),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_945),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_1003),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_915),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1002),
.B(n_1009),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_851),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_SL g1109 ( 
.A(n_859),
.B(n_279),
.C(n_277),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_945),
.Y(n_1110)
);

AND2x6_ASAP7_75t_L g1111 ( 
.A(n_853),
.B(n_699),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1002),
.B(n_832),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_839),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_915),
.B(n_832),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_869),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_953),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_963),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_994),
.Y(n_1118)
);

INVxp67_ASAP7_75t_SL g1119 ( 
.A(n_881),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_881),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_875),
.A2(n_382),
.B(n_383),
.C(n_380),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_852),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_953),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_963),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_976),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_R g1126 ( 
.A(n_970),
.B(n_971),
.Y(n_1126)
);

OR2x2_ASAP7_75t_SL g1127 ( 
.A(n_864),
.B(n_380),
.Y(n_1127)
);

NAND3xp33_ASAP7_75t_SL g1128 ( 
.A(n_846),
.B(n_283),
.C(n_281),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_978),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_968),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_881),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_SL g1132 ( 
.A1(n_990),
.A2(n_980),
.B1(n_903),
.B2(n_972),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_L g1133 ( 
.A(n_846),
.B(n_296),
.C(n_292),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_968),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_1005),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_915),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_956),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_876),
.A2(n_694),
.B1(n_734),
.B2(n_833),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_967),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_967),
.Y(n_1140)
);

NOR2x2_ASAP7_75t_L g1141 ( 
.A(n_851),
.B(n_321),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_R g1142 ( 
.A(n_848),
.B(n_299),
.Y(n_1142)
);

BUFx2_ASAP7_75t_SL g1143 ( 
.A(n_978),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_956),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_959),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_893),
.B(n_699),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_985),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_959),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_893),
.B(n_699),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_908),
.B(n_699),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_985),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1009),
.B(n_833),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_987),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_982),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_889),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_931),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_914),
.B(n_704),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_987),
.B(n_935),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_985),
.Y(n_1159)
);

BUFx12f_ASAP7_75t_L g1160 ( 
.A(n_991),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_982),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_920),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_923),
.B(n_704),
.Y(n_1163)
);

BUFx12f_ASAP7_75t_L g1164 ( 
.A(n_991),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_897),
.A2(n_734),
.B1(n_751),
.B2(n_750),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_923),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_986),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_986),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1008),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_927),
.A2(n_816),
.B(n_778),
.C(n_833),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_888),
.A2(n_734),
.B1(n_751),
.B2(n_750),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_924),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_924),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_936),
.B(n_805),
.Y(n_1174)
);

NOR2x1_ASAP7_75t_L g1175 ( 
.A(n_973),
.B(n_825),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1008),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_897),
.B(n_419),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_949),
.B(n_738),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_949),
.B(n_704),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_921),
.A2(n_734),
.B1(n_751),
.B2(n_750),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_951),
.B(n_704),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_951),
.Y(n_1182)
);

BUFx4f_ASAP7_75t_L g1183 ( 
.A(n_991),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_849),
.B(n_704),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_952),
.B(n_719),
.Y(n_1185)
);

BUFx10_ASAP7_75t_L g1186 ( 
.A(n_934),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_952),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_940),
.B(n_719),
.Y(n_1188)
);

OR2x4_ASAP7_75t_L g1189 ( 
.A(n_882),
.B(n_382),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_983),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_921),
.A2(n_751),
.B1(n_750),
.B2(n_826),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_857),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_936),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_991),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1011),
.Y(n_1195)
);

NAND2xp33_ASAP7_75t_SL g1196 ( 
.A(n_855),
.B(n_451),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_922),
.B(n_719),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_934),
.B(n_805),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1004),
.B(n_738),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1011),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_925),
.B(n_863),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_947),
.A2(n_751),
.B1(n_750),
.B2(n_754),
.Y(n_1202)
);

INVxp67_ASAP7_75t_SL g1203 ( 
.A(n_929),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1132),
.A2(n_904),
.B1(n_911),
.B2(n_875),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_1143),
.B(n_934),
.Y(n_1205)
);

AO21x1_ASAP7_75t_L g1206 ( 
.A1(n_1199),
.A2(n_860),
.B(n_894),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_1199),
.A2(n_984),
.A3(n_896),
.B(n_866),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1019),
.B(n_1004),
.Y(n_1208)
);

O2A1O1Ixp5_ASAP7_75t_L g1209 ( 
.A1(n_1060),
.A2(n_902),
.B(n_909),
.C(n_862),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1057),
.A2(n_1060),
.B(n_1088),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1035),
.A2(n_933),
.B(n_894),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1201),
.A2(n_942),
.B(n_941),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1013),
.A2(n_858),
.B1(n_861),
.B2(n_878),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1094),
.A2(n_989),
.B(n_955),
.Y(n_1214)
);

NAND2x1p5_ASAP7_75t_L g1215 ( 
.A(n_1120),
.B(n_910),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1184),
.A2(n_944),
.B(n_960),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1025),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1156),
.B(n_913),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1197),
.A2(n_1184),
.B(n_1146),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1031),
.A2(n_1071),
.B(n_1203),
.Y(n_1220)
);

NOR2xp67_ASAP7_75t_L g1221 ( 
.A(n_1037),
.B(n_998),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1070),
.B(n_934),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1019),
.B(n_962),
.Y(n_1223)
);

OA21x2_ASAP7_75t_L g1224 ( 
.A1(n_1081),
.A2(n_946),
.B(n_977),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1196),
.A2(n_944),
.B(n_981),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1103),
.A2(n_958),
.B(n_954),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1149),
.A2(n_1157),
.B(n_1150),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1163),
.A2(n_886),
.B(n_885),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1079),
.A2(n_907),
.B(n_916),
.Y(n_1229)
);

NAND2x1p5_ASAP7_75t_L g1230 ( 
.A(n_1120),
.B(n_917),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1120),
.A2(n_749),
.B(n_738),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1080),
.B(n_891),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1196),
.A2(n_884),
.B(n_993),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1121),
.A2(n_979),
.A3(n_999),
.B(n_996),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1044),
.B(n_962),
.Y(n_1235)
);

O2A1O1Ixp5_ASAP7_75t_L g1236 ( 
.A1(n_1082),
.A2(n_892),
.B(n_1010),
.C(n_950),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1044),
.B(n_948),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1115),
.A2(n_1001),
.B(n_749),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1117),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1179),
.A2(n_716),
.B(n_698),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1193),
.A2(n_1006),
.B(n_948),
.C(n_899),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1177),
.B(n_899),
.Y(n_1242)
);

NAND2x1p5_ASAP7_75t_L g1243 ( 
.A(n_1120),
.B(n_749),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_SL g1244 ( 
.A(n_1012),
.B(n_419),
.Y(n_1244)
);

AOI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1079),
.A2(n_723),
.B(n_716),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1158),
.B(n_938),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1117),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1090),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1158),
.A2(n_992),
.B(n_965),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1124),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1067),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1158),
.B(n_723),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1181),
.A2(n_735),
.B(n_729),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1070),
.B(n_541),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1084),
.A2(n_754),
.B1(n_719),
.B2(n_742),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1032),
.B(n_729),
.Y(n_1256)
);

AOI21xp33_ASAP7_75t_L g1257 ( 
.A1(n_1133),
.A2(n_302),
.B(n_300),
.Y(n_1257)
);

AOI221x1_ASAP7_75t_L g1258 ( 
.A1(n_1128),
.A2(n_432),
.B1(n_437),
.B2(n_442),
.C(n_425),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1124),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1032),
.B(n_735),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1130),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1121),
.A2(n_383),
.B(n_392),
.C(n_403),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1130),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1087),
.A2(n_754),
.B1(n_750),
.B2(n_751),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1046),
.B(n_541),
.Y(n_1265)
);

NAND2x1_ASAP7_75t_L g1266 ( 
.A(n_1131),
.B(n_719),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1185),
.A2(n_740),
.B(n_739),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1131),
.B(n_804),
.Y(n_1268)
);

OAI21xp33_ASAP7_75t_L g1269 ( 
.A1(n_1078),
.A2(n_308),
.B(n_304),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1134),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_SL g1271 ( 
.A1(n_1131),
.A2(n_410),
.B(n_408),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1156),
.B(n_742),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1134),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1026),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1188),
.A2(n_740),
.B(n_739),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_SL g1276 ( 
.A(n_1186),
.Y(n_1276)
);

OR2x6_ASAP7_75t_L g1277 ( 
.A(n_1096),
.B(n_1098),
.Y(n_1277)
);

AND3x1_ASAP7_75t_SL g1278 ( 
.A(n_1083),
.B(n_421),
.C(n_418),
.Y(n_1278)
);

AOI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1093),
.A2(n_762),
.B(n_759),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1122),
.B(n_309),
.Y(n_1280)
);

NOR2xp67_ASAP7_75t_SL g1281 ( 
.A(n_1049),
.B(n_451),
.Y(n_1281)
);

BUFx12f_ASAP7_75t_L g1282 ( 
.A(n_1096),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1106),
.B(n_542),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1126),
.B(n_419),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1093),
.A2(n_762),
.B(n_759),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1032),
.B(n_767),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1091),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1129),
.B(n_767),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1126),
.B(n_419),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1087),
.A2(n_742),
.B1(n_772),
.B2(n_852),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1073),
.A2(n_787),
.B(n_773),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1178),
.A2(n_787),
.A3(n_793),
.B(n_819),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1082),
.A2(n_793),
.B(n_773),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1153),
.B(n_809),
.Y(n_1294)
);

NAND2x1p5_ASAP7_75t_L g1295 ( 
.A(n_1115),
.B(n_804),
.Y(n_1295)
);

BUFx12f_ASAP7_75t_L g1296 ( 
.A(n_1098),
.Y(n_1296)
);

AO21x1_ASAP7_75t_L g1297 ( 
.A1(n_1043),
.A2(n_1178),
.B(n_1054),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1018),
.B(n_809),
.Y(n_1298)
);

OA22x2_ASAP7_75t_L g1299 ( 
.A1(n_1028),
.A2(n_882),
.B1(n_399),
.B2(n_398),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1114),
.B(n_451),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1170),
.A2(n_815),
.B(n_813),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1125),
.B(n_542),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1026),
.Y(n_1303)
);

AO21x1_ASAP7_75t_L g1304 ( 
.A1(n_1162),
.A2(n_796),
.B(n_813),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_SL g1305 ( 
.A1(n_1119),
.A2(n_772),
.B(n_742),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1097),
.A2(n_819),
.B(n_815),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1041),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1067),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1012),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1156),
.B(n_742),
.Y(n_1310)
);

NOR2xp67_ASAP7_75t_SL g1311 ( 
.A(n_1049),
.B(n_772),
.Y(n_1311)
);

INVx5_ASAP7_75t_L g1312 ( 
.A(n_1111),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1115),
.A2(n_772),
.B(n_804),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1166),
.A2(n_772),
.B1(n_829),
.B2(n_834),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_1102),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1042),
.B(n_545),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1097),
.A2(n_829),
.B(n_796),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1078),
.B(n_545),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1063),
.A2(n_646),
.B(n_645),
.Y(n_1319)
);

NAND2xp33_ASAP7_75t_L g1320 ( 
.A(n_1111),
.B(n_318),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1172),
.A2(n_829),
.B1(n_834),
.B2(n_794),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1049),
.A2(n_834),
.B(n_794),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1041),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_1067),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1018),
.B(n_1173),
.Y(n_1325)
);

NAND3xp33_ASAP7_75t_L g1326 ( 
.A(n_1033),
.B(n_1109),
.C(n_1050),
.Y(n_1326)
);

AO32x2_ASAP7_75t_L g1327 ( 
.A1(n_1040),
.A2(n_15),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1018),
.B(n_834),
.Y(n_1328)
);

AO21x1_ASAP7_75t_L g1329 ( 
.A1(n_1182),
.A2(n_550),
.B(n_547),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1063),
.A2(n_664),
.B(n_646),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1048),
.Y(n_1331)
);

AOI21xp33_ASAP7_75t_L g1332 ( 
.A1(n_1105),
.A2(n_1135),
.B(n_1156),
.Y(n_1332)
);

BUFx8_ASAP7_75t_L g1333 ( 
.A(n_1108),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1139),
.A2(n_646),
.B(n_550),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1192),
.B(n_794),
.Y(n_1335)
);

CKINVDCx8_ASAP7_75t_R g1336 ( 
.A(n_1036),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1187),
.A2(n_567),
.A3(n_578),
.B(n_547),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1107),
.B(n_834),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1042),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1014),
.A2(n_1022),
.B(n_1021),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1194),
.B(n_552),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1139),
.A2(n_556),
.B(n_552),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1048),
.A2(n_1055),
.B(n_1053),
.Y(n_1343)
);

NAND2x1p5_ASAP7_75t_L g1344 ( 
.A(n_1061),
.B(n_794),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1192),
.B(n_794),
.Y(n_1345)
);

AO22x2_ASAP7_75t_L g1346 ( 
.A1(n_1116),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1053),
.A2(n_393),
.B(n_389),
.C(n_378),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1055),
.A2(n_569),
.A3(n_578),
.B(n_556),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1140),
.A2(n_572),
.B(n_564),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1192),
.B(n_318),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1049),
.A2(n_722),
.B(n_831),
.Y(n_1351)
);

A2O1A1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1074),
.A2(n_374),
.B(n_371),
.C(n_369),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1015),
.A2(n_1107),
.B1(n_1174),
.B2(n_1072),
.Y(n_1353)
);

NAND2x2_ASAP7_75t_L g1354 ( 
.A(n_1106),
.B(n_310),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1140),
.A2(n_572),
.B(n_564),
.Y(n_1355)
);

AOI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1024),
.A2(n_573),
.B(n_567),
.Y(n_1356)
);

OAI21xp33_ASAP7_75t_L g1357 ( 
.A1(n_1142),
.A2(n_1017),
.B(n_1027),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1074),
.A2(n_569),
.B(n_573),
.Y(n_1358)
);

AOI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1029),
.A2(n_805),
.B(n_722),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1154),
.A2(n_1167),
.B(n_1161),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1154),
.A2(n_805),
.B(n_722),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1066),
.A2(n_722),
.B(n_831),
.Y(n_1362)
);

AO21x2_ASAP7_75t_L g1363 ( 
.A1(n_1030),
.A2(n_1059),
.B(n_1038),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1160),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1107),
.B(n_315),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1161),
.A2(n_1168),
.B(n_1167),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1174),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1240),
.A2(n_1175),
.B(n_1095),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1223),
.B(n_1192),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1253),
.A2(n_1095),
.B(n_1089),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1312),
.Y(n_1371)
);

AO21x2_ASAP7_75t_L g1372 ( 
.A1(n_1297),
.A2(n_1301),
.B(n_1304),
.Y(n_1372)
);

AO21x2_ASAP7_75t_L g1373 ( 
.A1(n_1206),
.A2(n_1064),
.B(n_1062),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1353),
.B(n_1136),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1336),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1267),
.A2(n_1110),
.B(n_1089),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1223),
.B(n_1068),
.Y(n_1377)
);

NOR2x1_ASAP7_75t_L g1378 ( 
.A(n_1339),
.B(n_1047),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1208),
.B(n_1102),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1220),
.A2(n_1180),
.B(n_1165),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1239),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1343),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1312),
.B(n_1034),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1367),
.B(n_1136),
.Y(n_1384)
);

AO21x2_ASAP7_75t_L g1385 ( 
.A1(n_1291),
.A2(n_1075),
.B(n_1069),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1245),
.A2(n_1279),
.B(n_1226),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1367),
.B(n_1222),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1217),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1242),
.B(n_1110),
.Y(n_1389)
);

AO31x2_ASAP7_75t_L g1390 ( 
.A1(n_1329),
.A2(n_1104),
.A3(n_1100),
.B(n_1086),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1214),
.A2(n_1092),
.B(n_1168),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1287),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1219),
.A2(n_1176),
.B(n_1169),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1250),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1208),
.B(n_1113),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1305),
.A2(n_1066),
.B(n_1067),
.Y(n_1396)
);

NAND3xp33_ASAP7_75t_L g1397 ( 
.A(n_1257),
.B(n_1326),
.C(n_1204),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1210),
.A2(n_1176),
.B(n_1169),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1229),
.A2(n_1137),
.B(n_1123),
.Y(n_1399)
);

AOI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1225),
.A2(n_1200),
.B(n_1195),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1250),
.B(n_1015),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1318),
.B(n_1015),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1222),
.B(n_1061),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1309),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1284),
.A2(n_1144),
.B(n_1145),
.C(n_1148),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1312),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1309),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1324),
.Y(n_1408)
);

INVxp67_ASAP7_75t_L g1409 ( 
.A(n_1316),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1343),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_SL g1411 ( 
.A1(n_1271),
.A2(n_1099),
.B(n_1191),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1315),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1273),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1315),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1360),
.A2(n_1020),
.B(n_1016),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_SL g1416 ( 
.A1(n_1241),
.A2(n_1016),
.B(n_1020),
.C(n_1039),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1251),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1237),
.A2(n_1183),
.B1(n_1023),
.B2(n_1174),
.Y(n_1418)
);

NAND2x1p5_ASAP7_75t_L g1419 ( 
.A(n_1312),
.B(n_1034),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1235),
.B(n_1190),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1251),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1273),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1302),
.B(n_1190),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1251),
.Y(n_1424)
);

OAI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1244),
.A2(n_1183),
.B1(n_1155),
.B2(n_1113),
.C(n_1138),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1331),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1247),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1259),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1261),
.B(n_1058),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1209),
.A2(n_1202),
.B(n_1171),
.Y(n_1430)
);

NOR2x1_ASAP7_75t_R g1431 ( 
.A(n_1282),
.B(n_1160),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1324),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1236),
.A2(n_1072),
.B(n_1058),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1358),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1366),
.A2(n_1020),
.B(n_1016),
.Y(n_1435)
);

AOI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1225),
.A2(n_1072),
.B(n_1058),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1333),
.Y(n_1437)
);

NOR2xp67_ASAP7_75t_L g1438 ( 
.A(n_1232),
.B(n_1164),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1340),
.A2(n_1076),
.B(n_1039),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_SL g1440 ( 
.A1(n_1216),
.A2(n_1099),
.B(n_1159),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1331),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1289),
.A2(n_1047),
.B(n_1114),
.C(n_1112),
.Y(n_1442)
);

BUFx12f_ASAP7_75t_L g1443 ( 
.A(n_1282),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1357),
.A2(n_1085),
.B1(n_1112),
.B2(n_1152),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_SL g1445 ( 
.A1(n_1211),
.A2(n_1099),
.B(n_1159),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1334),
.A2(n_1076),
.B(n_1039),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1231),
.A2(n_1066),
.B(n_1077),
.Y(n_1447)
);

AO21x2_ASAP7_75t_L g1448 ( 
.A1(n_1233),
.A2(n_1142),
.B(n_1101),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1209),
.A2(n_1101),
.B(n_1085),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1358),
.Y(n_1450)
);

INVxp67_ASAP7_75t_SL g1451 ( 
.A(n_1311),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1333),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1263),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1270),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1274),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1358),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1296),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1303),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1241),
.B(n_1085),
.Y(n_1459)
);

NAND2x1p5_ASAP7_75t_L g1460 ( 
.A(n_1272),
.B(n_1034),
.Y(n_1460)
);

AO31x2_ASAP7_75t_L g1461 ( 
.A1(n_1213),
.A2(n_1159),
.A3(n_1045),
.B(n_1127),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1228),
.A2(n_1076),
.B(n_1147),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1307),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1248),
.Y(n_1464)
);

AOI32xp33_ASAP7_75t_L g1465 ( 
.A1(n_1346),
.A2(n_1155),
.A3(n_317),
.B1(n_409),
.B2(n_413),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1243),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1254),
.B(n_1114),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1293),
.A2(n_1236),
.B(n_1233),
.Y(n_1468)
);

BUFx8_ASAP7_75t_L g1469 ( 
.A(n_1276),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1254),
.B(n_1114),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_L g1471 ( 
.A(n_1258),
.B(n_331),
.C(n_328),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1323),
.Y(n_1472)
);

NOR2xp67_ASAP7_75t_L g1473 ( 
.A(n_1365),
.B(n_1164),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1325),
.B(n_1190),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1317),
.A2(n_1066),
.B(n_1077),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1243),
.Y(n_1476)
);

AOI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1269),
.A2(n_1052),
.B1(n_333),
.B2(n_434),
.C(n_334),
.Y(n_1477)
);

INVxp67_ASAP7_75t_SL g1478 ( 
.A(n_1251),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1361),
.A2(n_1151),
.B(n_1147),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1342),
.Y(n_1480)
);

AOI21xp33_ASAP7_75t_L g1481 ( 
.A1(n_1280),
.A2(n_1112),
.B(n_1101),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1283),
.B(n_1152),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1313),
.A2(n_1077),
.B(n_1118),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1332),
.B(n_1190),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1348),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1341),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1280),
.A2(n_1097),
.B1(n_1186),
.B2(n_1198),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1285),
.A2(n_1151),
.B(n_1147),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1227),
.A2(n_1330),
.B(n_1319),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1218),
.A2(n_1198),
.B(n_1111),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1299),
.A2(n_1097),
.B1(n_1186),
.B2(n_1198),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1348),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1348),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1238),
.A2(n_1151),
.B(n_1111),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1348),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_SL g1496 ( 
.A1(n_1359),
.A2(n_1097),
.B(n_1111),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1288),
.B(n_1034),
.Y(n_1497)
);

AO21x2_ASAP7_75t_L g1498 ( 
.A1(n_1218),
.A2(n_1017),
.B(n_1052),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1299),
.A2(n_1065),
.B1(n_1056),
.B2(n_318),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1252),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1238),
.A2(n_1056),
.B(n_1065),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1337),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1313),
.A2(n_1118),
.B(n_1077),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1349),
.Y(n_1504)
);

NOR2x1_ASAP7_75t_SL g1505 ( 
.A(n_1363),
.B(n_1118),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1308),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1249),
.A2(n_1056),
.B(n_1065),
.C(n_1118),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1265),
.B(n_1189),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1355),
.A2(n_1065),
.B(n_1056),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1350),
.A2(n_788),
.B(n_722),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1350),
.A2(n_788),
.B(n_407),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1337),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1278),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1364),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1283),
.Y(n_1515)
);

AOI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1356),
.A2(n_788),
.B(n_435),
.Y(n_1516)
);

INVx6_ASAP7_75t_L g1517 ( 
.A(n_1308),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1363),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1337),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1337),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1294),
.Y(n_1521)
);

BUFx10_ASAP7_75t_L g1522 ( 
.A(n_1276),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1234),
.Y(n_1523)
);

A2O1A1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1347),
.A2(n_405),
.B(n_345),
.C(n_347),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1275),
.A2(n_435),
.B(n_318),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1277),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1256),
.Y(n_1527)
);

AO21x2_ASAP7_75t_L g1528 ( 
.A1(n_1306),
.A2(n_318),
.B(n_435),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1322),
.A2(n_435),
.B(n_318),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1246),
.A2(n_1205),
.B1(n_1328),
.B2(n_1221),
.Y(n_1530)
);

O2A1O1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1347),
.A2(n_1141),
.B(n_1051),
.C(n_448),
.Y(n_1531)
);

O2A1O1Ixp33_ASAP7_75t_SL g1532 ( 
.A1(n_1352),
.A2(n_1141),
.B(n_435),
.C(n_229),
.Y(n_1532)
);

BUFx4f_ASAP7_75t_L g1533 ( 
.A(n_1308),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1322),
.A2(n_435),
.B(n_799),
.Y(n_1534)
);

AO31x2_ASAP7_75t_L g1535 ( 
.A1(n_1262),
.A2(n_435),
.A3(n_26),
.B(n_27),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1308),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1260),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1286),
.Y(n_1538)
);

A2O1A1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1352),
.A2(n_406),
.B(n_353),
.C(n_445),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1298),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1205),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1338),
.A2(n_788),
.B(n_352),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1212),
.B(n_1224),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1314),
.A2(n_435),
.B(n_799),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1234),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1234),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1234),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1321),
.A2(n_1362),
.B(n_1351),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1277),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1351),
.A2(n_435),
.B(n_799),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1427),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1397),
.A2(n_1346),
.B1(n_1354),
.B2(n_1205),
.Y(n_1552)
);

AO21x2_ASAP7_75t_L g1553 ( 
.A1(n_1436),
.A2(n_1320),
.B(n_1345),
.Y(n_1553)
);

INVx4_ASAP7_75t_L g1554 ( 
.A(n_1533),
.Y(n_1554)
);

AOI222xp33_ASAP7_75t_L g1555 ( 
.A1(n_1379),
.A2(n_1395),
.B1(n_1409),
.B2(n_1477),
.C1(n_1508),
.C2(n_1346),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1436),
.A2(n_1272),
.B(n_1310),
.Y(n_1556)
);

CKINVDCx6p67_ASAP7_75t_R g1557 ( 
.A(n_1443),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1388),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1533),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1428),
.Y(n_1560)
);

AOI332xp33_ASAP7_75t_L g1561 ( 
.A1(n_1465),
.A2(n_1278),
.A3(n_1327),
.B1(n_367),
.B2(n_375),
.B3(n_376),
.C1(n_394),
.C2(n_396),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1533),
.Y(n_1562)
);

BUFx8_ASAP7_75t_L g1563 ( 
.A(n_1443),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1507),
.A2(n_1396),
.B(n_1475),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1453),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1389),
.B(n_1212),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1403),
.B(n_1277),
.Y(n_1567)
);

NAND2x1p5_ASAP7_75t_L g1568 ( 
.A(n_1408),
.B(n_1310),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_SL g1569 ( 
.A1(n_1513),
.A2(n_1354),
.B1(n_1320),
.B2(n_1300),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1389),
.B(n_1212),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1403),
.B(n_1300),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1371),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1471),
.A2(n_366),
.B1(n_363),
.B2(n_397),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1453),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1369),
.B(n_1335),
.Y(n_1575)
);

CKINVDCx16_ASAP7_75t_R g1576 ( 
.A(n_1437),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1447),
.A2(n_1295),
.B(n_1268),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1402),
.B(n_1335),
.Y(n_1578)
);

NAND2x1p5_ASAP7_75t_L g1579 ( 
.A(n_1408),
.B(n_1345),
.Y(n_1579)
);

OR2x6_ASAP7_75t_L g1580 ( 
.A(n_1442),
.B(n_1300),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_SL g1581 ( 
.A(n_1531),
.B(n_420),
.C(n_422),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1422),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1459),
.A2(n_430),
.B1(n_441),
.B2(n_438),
.Y(n_1583)
);

OAI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1425),
.A2(n_1290),
.B1(n_440),
.B2(n_1264),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_SL g1585 ( 
.A1(n_1513),
.A2(n_1327),
.B1(n_1215),
.B2(n_1230),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1375),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1459),
.A2(n_1224),
.B1(n_1327),
.B2(n_1215),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1486),
.B(n_1327),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1380),
.A2(n_1295),
.B(n_1268),
.Y(n_1589)
);

NOR3xp33_ASAP7_75t_SL g1590 ( 
.A(n_1404),
.B(n_1255),
.C(n_1362),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1377),
.A2(n_1224),
.B1(n_1230),
.B2(n_1344),
.Y(n_1591)
);

NOR2xp67_ASAP7_75t_L g1592 ( 
.A(n_1392),
.B(n_110),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1522),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_1375),
.Y(n_1594)
);

CKINVDCx8_ASAP7_75t_R g1595 ( 
.A(n_1404),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1417),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1377),
.A2(n_1481),
.B1(n_1521),
.B2(n_1498),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1388),
.Y(n_1598)
);

OAI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1524),
.A2(n_1266),
.B1(n_1281),
.B2(n_1207),
.C(n_32),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1541),
.B(n_1374),
.Y(n_1600)
);

OAI22x1_ASAP7_75t_L g1601 ( 
.A1(n_1541),
.A2(n_1207),
.B1(n_1292),
.B2(n_29),
.Y(n_1601)
);

AOI21x1_ASAP7_75t_L g1602 ( 
.A1(n_1400),
.A2(n_1207),
.B(n_1292),
.Y(n_1602)
);

CKINVDCx6p67_ASAP7_75t_R g1603 ( 
.A(n_1437),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1464),
.B(n_1207),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1423),
.B(n_21),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1420),
.B(n_1292),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1403),
.B(n_1292),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_1469),
.Y(n_1608)
);

AO31x2_ASAP7_75t_L g1609 ( 
.A1(n_1502),
.A2(n_788),
.A3(n_29),
.B(n_33),
.Y(n_1609)
);

NOR2x1_ASAP7_75t_SL g1610 ( 
.A(n_1530),
.B(n_799),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1498),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1386),
.A2(n_831),
.B(n_799),
.Y(n_1612)
);

AOI21xp33_ASAP7_75t_L g1613 ( 
.A1(n_1405),
.A2(n_35),
.B(n_39),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1454),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1500),
.B(n_39),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1514),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1382),
.Y(n_1617)
);

OAI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1515),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_1618)
);

AOI222xp33_ASAP7_75t_L g1619 ( 
.A1(n_1438),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.C1(n_48),
.C2(n_49),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1517),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1444),
.A2(n_831),
.B1(n_48),
.B2(n_49),
.Y(n_1621)
);

AO21x2_ASAP7_75t_L g1622 ( 
.A1(n_1400),
.A2(n_788),
.B(n_184),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1387),
.B(n_46),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_SL g1624 ( 
.A1(n_1498),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1374),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1387),
.B(n_59),
.Y(n_1626)
);

INVx4_ASAP7_75t_SL g1627 ( 
.A(n_1517),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1454),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1484),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1374),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1401),
.B(n_62),
.Y(n_1631)
);

INVx4_ASAP7_75t_L g1632 ( 
.A(n_1417),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1378),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1527),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1371),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1455),
.Y(n_1636)
);

BUFx12f_ASAP7_75t_L g1637 ( 
.A(n_1412),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1371),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1517),
.Y(n_1639)
);

AO31x2_ASAP7_75t_L g1640 ( 
.A1(n_1502),
.A2(n_72),
.A3(n_73),
.B(n_74),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1455),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1500),
.B(n_75),
.Y(n_1642)
);

OAI222xp33_ASAP7_75t_L g1643 ( 
.A1(n_1418),
.A2(n_1474),
.B1(n_1499),
.B2(n_1487),
.C1(n_1491),
.C2(n_1538),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_1412),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1527),
.A2(n_1537),
.B1(n_1538),
.B2(n_1540),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1407),
.A2(n_831),
.B1(n_76),
.B2(n_77),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1537),
.B(n_75),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1514),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1467),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_1649)
);

AO31x2_ASAP7_75t_L g1650 ( 
.A1(n_1512),
.A2(n_79),
.A3(n_81),
.B(n_82),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1410),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1467),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_1652)
);

NAND2xp33_ASAP7_75t_SL g1653 ( 
.A(n_1432),
.B(n_84),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1467),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1470),
.B(n_146),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1401),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1429),
.B(n_88),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1429),
.B(n_88),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1536),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1458),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1417),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1407),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1482),
.B(n_91),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1474),
.B(n_93),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1470),
.A2(n_95),
.B1(n_98),
.B2(n_100),
.Y(n_1665)
);

INVx4_ASAP7_75t_L g1666 ( 
.A(n_1417),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1470),
.A2(n_95),
.B1(n_100),
.B2(n_102),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1410),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1482),
.A2(n_104),
.B1(n_105),
.B2(n_116),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_SL g1670 ( 
.A(n_1539),
.B(n_126),
.C(n_127),
.Y(n_1670)
);

CKINVDCx16_ASAP7_75t_R g1671 ( 
.A(n_1452),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1482),
.B(n_130),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1384),
.B(n_1473),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1384),
.B(n_1497),
.Y(n_1674)
);

XNOR2xp5_ASAP7_75t_L g1675 ( 
.A(n_1414),
.B(n_138),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1432),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1526),
.A2(n_145),
.B1(n_148),
.B2(n_158),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1532),
.A2(n_163),
.B1(n_169),
.B2(n_179),
.C(n_191),
.Y(n_1678)
);

AOI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1416),
.A2(n_193),
.B1(n_198),
.B2(n_199),
.C(n_202),
.Y(n_1679)
);

OAI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1452),
.A2(n_204),
.B1(n_210),
.B2(n_213),
.Y(n_1680)
);

OAI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1526),
.A2(n_217),
.B1(n_224),
.B2(n_225),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1384),
.B(n_1497),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1381),
.B(n_1394),
.Y(n_1683)
);

OAI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1386),
.A2(n_1489),
.B(n_1391),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1536),
.B(n_1458),
.Y(n_1685)
);

OAI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1433),
.A2(n_1542),
.B(n_1511),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1468),
.A2(n_1385),
.B(n_1503),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1381),
.B(n_1394),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1413),
.B(n_1426),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1451),
.A2(n_1549),
.B1(n_1472),
.B2(n_1463),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1468),
.A2(n_1385),
.B(n_1483),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_SL g1692 ( 
.A1(n_1469),
.A2(n_1549),
.B1(n_1522),
.B2(n_1457),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1413),
.B(n_1426),
.Y(n_1693)
);

OAI222xp33_ASAP7_75t_L g1694 ( 
.A1(n_1441),
.A2(n_1414),
.B1(n_1546),
.B2(n_1460),
.C1(n_1545),
.C2(n_1547),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1441),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1461),
.B(n_1478),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1512),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1523),
.A2(n_1547),
.B1(n_1545),
.B2(n_1546),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1461),
.B(n_1421),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1461),
.B(n_1421),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1523),
.A2(n_1372),
.B1(n_1468),
.B2(n_1469),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1434),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1506),
.B(n_1461),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1372),
.A2(n_1468),
.B1(n_1528),
.B2(n_1518),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1519),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1519),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1506),
.B(n_1461),
.Y(n_1707)
);

OR2x6_ASAP7_75t_L g1708 ( 
.A(n_1411),
.B(n_1440),
.Y(n_1708)
);

NAND2xp33_ASAP7_75t_SL g1709 ( 
.A(n_1406),
.B(n_1490),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1522),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1535),
.B(n_1417),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1520),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1424),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1424),
.B(n_1490),
.Y(n_1714)
);

OAI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1457),
.A2(n_1466),
.B1(n_1476),
.B2(n_1406),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1535),
.B(n_1424),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1489),
.A2(n_1391),
.B(n_1368),
.Y(n_1717)
);

AOI222xp33_ASAP7_75t_L g1718 ( 
.A1(n_1431),
.A2(n_1520),
.B1(n_1411),
.B2(n_1493),
.C1(n_1495),
.C2(n_1485),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1460),
.A2(n_1419),
.B1(n_1383),
.B2(n_1476),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1518),
.A2(n_1372),
.B1(n_1528),
.B2(n_1495),
.C(n_1492),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1517),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1434),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1485),
.Y(n_1723)
);

BUFx8_ASAP7_75t_SL g1724 ( 
.A(n_1424),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1460),
.A2(n_1419),
.B1(n_1383),
.B2(n_1476),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1535),
.B(n_1424),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1383),
.Y(n_1727)
);

NAND2x1p5_ASAP7_75t_L g1728 ( 
.A(n_1466),
.B(n_1449),
.Y(n_1728)
);

A2O1A1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1525),
.A2(n_1399),
.B(n_1529),
.C(n_1510),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1490),
.A2(n_1448),
.B1(n_1449),
.B2(n_1373),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_SL g1731 ( 
.A1(n_1448),
.A2(n_1528),
.B1(n_1445),
.B2(n_1505),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1419),
.A2(n_1430),
.B1(n_1449),
.B2(n_1543),
.Y(n_1732)
);

BUFx2_ASAP7_75t_L g1733 ( 
.A(n_1449),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1492),
.Y(n_1734)
);

AOI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1480),
.A2(n_1504),
.B(n_1493),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1448),
.B(n_1373),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1535),
.B(n_1525),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1385),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1450),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1445),
.A2(n_1440),
.B(n_1505),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1450),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1430),
.A2(n_1480),
.B1(n_1504),
.B2(n_1456),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1555),
.A2(n_1373),
.B1(n_1430),
.B2(n_1529),
.Y(n_1743)
);

OAI221xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1649),
.A2(n_1456),
.B1(n_1430),
.B2(n_1390),
.C(n_1544),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_SL g1745 ( 
.A1(n_1585),
.A2(n_1496),
.B1(n_1544),
.B2(n_1494),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1605),
.B(n_1390),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1581),
.A2(n_1439),
.B1(n_1501),
.B2(n_1462),
.Y(n_1747)
);

AOI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1613),
.A2(n_1649),
.B1(n_1652),
.B2(n_1654),
.C(n_1665),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1583),
.A2(n_1516),
.B1(n_1390),
.B2(n_1496),
.C(n_1548),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1619),
.A2(n_1393),
.B1(n_1398),
.B2(n_1370),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1652),
.A2(n_1393),
.B1(n_1398),
.B2(n_1370),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1654),
.A2(n_1390),
.B1(n_1376),
.B2(n_1516),
.C(n_1439),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1686),
.A2(n_1621),
.B1(n_1580),
.B2(n_1599),
.Y(n_1753)
);

OAI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1583),
.A2(n_1390),
.B1(n_1548),
.B2(n_1501),
.C(n_1462),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1656),
.B(n_1415),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1589),
.A2(n_1509),
.B(n_1415),
.Y(n_1756)
);

AND2x6_ASAP7_75t_SL g1757 ( 
.A(n_1605),
.B(n_1435),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1559),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1633),
.A2(n_1446),
.B1(n_1509),
.B2(n_1479),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1559),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_SL g1761 ( 
.A1(n_1580),
.A2(n_1534),
.B1(n_1550),
.B2(n_1488),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1674),
.B(n_1488),
.Y(n_1762)
);

CKINVDCx20_ASAP7_75t_R g1763 ( 
.A(n_1608),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1682),
.B(n_1534),
.Y(n_1764)
);

OAI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1662),
.A2(n_1479),
.B1(n_1550),
.B2(n_1580),
.Y(n_1765)
);

A2O1A1Ixp33_ASAP7_75t_L g1766 ( 
.A1(n_1679),
.A2(n_1678),
.B(n_1561),
.C(n_1653),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1565),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1575),
.B(n_1645),
.Y(n_1768)
);

AOI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1602),
.A2(n_1735),
.B(n_1601),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1667),
.A2(n_1625),
.B1(n_1630),
.B2(n_1634),
.Y(n_1770)
);

OAI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1667),
.A2(n_1630),
.B1(n_1625),
.B2(n_1552),
.C(n_1669),
.Y(n_1771)
);

AOI322xp5_ASAP7_75t_L g1772 ( 
.A1(n_1634),
.A2(n_1611),
.A3(n_1618),
.B1(n_1669),
.B2(n_1653),
.C1(n_1624),
.C2(n_1552),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_1608),
.Y(n_1773)
);

OAI211xp5_ASAP7_75t_SL g1774 ( 
.A1(n_1573),
.A2(n_1718),
.B(n_1569),
.C(n_1616),
.Y(n_1774)
);

OAI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1573),
.A2(n_1692),
.B1(n_1677),
.B2(n_1670),
.C(n_1597),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1646),
.A2(n_1642),
.B1(n_1615),
.B2(n_1647),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1575),
.B(n_1645),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1631),
.B(n_1657),
.Y(n_1778)
);

OAI322xp33_ASAP7_75t_L g1779 ( 
.A1(n_1604),
.A2(n_1664),
.A3(n_1560),
.B1(n_1551),
.B2(n_1707),
.C1(n_1703),
.C2(n_1680),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1578),
.B(n_1598),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1574),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1595),
.A2(n_1600),
.B1(n_1578),
.B2(n_1558),
.Y(n_1782)
);

BUFx3_ASAP7_75t_L g1783 ( 
.A(n_1724),
.Y(n_1783)
);

OAI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1600),
.A2(n_1671),
.B1(n_1576),
.B2(n_1584),
.Y(n_1784)
);

OAI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1597),
.A2(n_1590),
.B1(n_1592),
.B2(n_1593),
.C(n_1675),
.Y(n_1785)
);

OAI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1600),
.A2(n_1558),
.B1(n_1603),
.B2(n_1681),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1663),
.A2(n_1658),
.B1(n_1626),
.B2(n_1623),
.Y(n_1787)
);

OAI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1648),
.A2(n_1595),
.B1(n_1710),
.B2(n_1564),
.C(n_1591),
.Y(n_1788)
);

OAI211xp5_ASAP7_75t_L g1789 ( 
.A1(n_1701),
.A2(n_1587),
.B(n_1730),
.C(n_1696),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1676),
.Y(n_1790)
);

OAI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1603),
.A2(n_1570),
.B1(n_1566),
.B2(n_1690),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1577),
.A2(n_1687),
.B(n_1691),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1685),
.B(n_1673),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1655),
.A2(n_1567),
.B1(n_1571),
.B2(n_1557),
.Y(n_1794)
);

OAI222xp33_ASAP7_75t_L g1795 ( 
.A1(n_1655),
.A2(n_1587),
.B1(n_1588),
.B2(n_1701),
.C1(n_1562),
.C2(n_1554),
.Y(n_1795)
);

OAI211xp5_ASAP7_75t_L g1796 ( 
.A1(n_1591),
.A2(n_1737),
.B(n_1710),
.C(n_1641),
.Y(n_1796)
);

INVx5_ASAP7_75t_SL g1797 ( 
.A(n_1557),
.Y(n_1797)
);

OAI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1731),
.A2(n_1586),
.B1(n_1594),
.B2(n_1708),
.C(n_1672),
.Y(n_1798)
);

AO221x2_ASAP7_75t_L g1799 ( 
.A1(n_1694),
.A2(n_1643),
.B1(n_1715),
.B2(n_1732),
.C(n_1640),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1614),
.Y(n_1800)
);

OAI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1586),
.A2(n_1594),
.B1(n_1708),
.B2(n_1644),
.C(n_1554),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1655),
.A2(n_1567),
.B1(n_1571),
.B2(n_1563),
.Y(n_1802)
);

OAI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1554),
.A2(n_1562),
.B1(n_1660),
.B2(n_1636),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1567),
.A2(n_1563),
.B1(n_1637),
.B2(n_1607),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1724),
.Y(n_1805)
);

INVxp67_ASAP7_75t_SL g1806 ( 
.A(n_1683),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_SL g1807 ( 
.A1(n_1610),
.A2(n_1563),
.B1(n_1562),
.B2(n_1637),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_SL g1808 ( 
.A1(n_1711),
.A2(n_1716),
.B1(n_1726),
.B2(n_1559),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1644),
.A2(n_1579),
.B1(n_1568),
.B2(n_1559),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1607),
.A2(n_1628),
.B1(n_1606),
.B2(n_1695),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1607),
.A2(n_1700),
.B1(n_1699),
.B2(n_1582),
.Y(n_1811)
);

OR2x6_ASAP7_75t_L g1812 ( 
.A(n_1708),
.B(n_1740),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1729),
.A2(n_1553),
.B(n_1709),
.Y(n_1813)
);

OAI211xp5_ASAP7_75t_L g1814 ( 
.A1(n_1736),
.A2(n_1704),
.B(n_1720),
.C(n_1689),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1659),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1723),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1734),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1659),
.B(n_1721),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1714),
.B(n_1688),
.Y(n_1819)
);

AOI21xp33_ASAP7_75t_SL g1820 ( 
.A1(n_1620),
.A2(n_1639),
.B(n_1719),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1620),
.A2(n_1639),
.B1(n_1727),
.B2(n_1579),
.Y(n_1821)
);

OAI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1739),
.A2(n_1568),
.B1(n_1693),
.B2(n_1727),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_SL g1823 ( 
.A1(n_1725),
.A2(n_1727),
.B1(n_1572),
.B2(n_1635),
.Y(n_1823)
);

AOI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1704),
.A2(n_1698),
.B1(n_1742),
.B2(n_1709),
.C(n_1733),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1739),
.B(n_1705),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1698),
.A2(n_1635),
.B1(n_1638),
.B2(n_1572),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1697),
.B(n_1706),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1713),
.B(n_1627),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1582),
.A2(n_1738),
.B1(n_1553),
.B2(n_1712),
.Y(n_1829)
);

AOI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1738),
.A2(n_1729),
.B1(n_1741),
.B2(n_1638),
.C(n_1728),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1738),
.A2(n_1741),
.B1(n_1728),
.B2(n_1702),
.C(n_1722),
.Y(n_1831)
);

AOI21xp33_ASAP7_75t_L g1832 ( 
.A1(n_1622),
.A2(n_1556),
.B(n_1741),
.Y(n_1832)
);

AOI222xp33_ASAP7_75t_L g1833 ( 
.A1(n_1627),
.A2(n_1722),
.B1(n_1702),
.B2(n_1668),
.C1(n_1651),
.C2(n_1617),
.Y(n_1833)
);

OAI211xp5_ASAP7_75t_L g1834 ( 
.A1(n_1632),
.A2(n_1666),
.B(n_1650),
.C(n_1640),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1622),
.A2(n_1668),
.B1(n_1666),
.B2(n_1632),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1596),
.A2(n_1661),
.B1(n_1640),
.B2(n_1650),
.Y(n_1836)
);

AOI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1661),
.A2(n_1640),
.B1(n_1650),
.B2(n_1609),
.C(n_1717),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1661),
.A2(n_1650),
.B1(n_1609),
.B2(n_1684),
.Y(n_1838)
);

AOI221xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1609),
.A2(n_872),
.B1(n_1208),
.B2(n_1223),
.C(n_854),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1609),
.A2(n_1208),
.B1(n_1223),
.B2(n_1555),
.Y(n_1840)
);

OAI22xp33_ASAP7_75t_SL g1841 ( 
.A1(n_1612),
.A2(n_701),
.B1(n_1244),
.B2(n_1208),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1612),
.B(n_1208),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1629),
.B(n_1208),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1676),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1555),
.A2(n_1208),
.B1(n_1223),
.B2(n_1132),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1559),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1682),
.B(n_1659),
.Y(n_1847)
);

OAI21x1_ASAP7_75t_L g1848 ( 
.A1(n_1717),
.A2(n_1684),
.B(n_1436),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1555),
.A2(n_1208),
.B1(n_1223),
.B2(n_1132),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1583),
.A2(n_1132),
.B1(n_1223),
.B2(n_1208),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1585),
.A2(n_1208),
.B1(n_843),
.B2(n_1126),
.Y(n_1851)
);

OAI21xp33_ASAP7_75t_L g1852 ( 
.A1(n_1555),
.A2(n_872),
.B(n_843),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1629),
.B(n_1208),
.Y(n_1853)
);

OAI21x1_ASAP7_75t_L g1854 ( 
.A1(n_1717),
.A2(n_1684),
.B(n_1436),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_1598),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1583),
.A2(n_1132),
.B1(n_1223),
.B2(n_1208),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1676),
.Y(n_1857)
);

AOI221xp5_ASAP7_75t_L g1858 ( 
.A1(n_1613),
.A2(n_1208),
.B1(n_872),
.B2(n_1223),
.C(n_1465),
.Y(n_1858)
);

OR2x6_ASAP7_75t_L g1859 ( 
.A(n_1580),
.B(n_1708),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1555),
.A2(n_843),
.B1(n_872),
.B2(n_1132),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1555),
.A2(n_1208),
.B1(n_1223),
.B2(n_1132),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1629),
.B(n_1208),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1686),
.A2(n_872),
.B(n_1132),
.Y(n_1863)
);

AO31x2_ASAP7_75t_L g1864 ( 
.A1(n_1729),
.A2(n_1601),
.A3(n_1738),
.B(n_1742),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1629),
.B(n_1208),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_SL g1866 ( 
.A1(n_1585),
.A2(n_1208),
.B1(n_843),
.B2(n_1126),
.Y(n_1866)
);

INVx4_ASAP7_75t_L g1867 ( 
.A(n_1559),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1629),
.B(n_1208),
.Y(n_1868)
);

OAI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1662),
.A2(n_701),
.B1(n_1208),
.B2(n_846),
.Y(n_1869)
);

AOI322xp5_ASAP7_75t_L g1870 ( 
.A1(n_1625),
.A2(n_1208),
.A3(n_1223),
.B1(n_1630),
.B2(n_1654),
.C1(n_1652),
.C2(n_1649),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1676),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1656),
.B(n_1208),
.Y(n_1872)
);

CKINVDCx20_ASAP7_75t_R g1873 ( 
.A(n_1608),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1555),
.A2(n_843),
.B1(n_872),
.B2(n_1132),
.Y(n_1874)
);

AOI221x1_ASAP7_75t_SL g1875 ( 
.A1(n_1662),
.A2(n_1208),
.B1(n_1223),
.B2(n_872),
.C(n_458),
.Y(n_1875)
);

OAI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1662),
.A2(n_701),
.B1(n_1208),
.B2(n_846),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1686),
.A2(n_1589),
.B(n_1305),
.Y(n_1877)
);

INVxp67_ASAP7_75t_L g1878 ( 
.A(n_1598),
.Y(n_1878)
);

INVx5_ASAP7_75t_L g1879 ( 
.A(n_1724),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1629),
.B(n_1674),
.Y(n_1880)
);

AO221x2_ASAP7_75t_L g1881 ( 
.A1(n_1585),
.A2(n_1397),
.B1(n_1662),
.B2(n_1618),
.C(n_854),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1586),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1555),
.A2(n_1208),
.B1(n_1223),
.B2(n_1132),
.Y(n_1883)
);

OAI211xp5_ASAP7_75t_L g1884 ( 
.A1(n_1561),
.A2(n_1465),
.B(n_1555),
.C(n_1132),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_SL g1885 ( 
.A1(n_1608),
.A2(n_1395),
.B1(n_1379),
.B2(n_1132),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1555),
.A2(n_1208),
.B1(n_1223),
.B2(n_1132),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1682),
.B(n_1659),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_SL g1888 ( 
.A1(n_1608),
.A2(n_1395),
.B1(n_1379),
.B2(n_1132),
.Y(n_1888)
);

OAI221xp5_ASAP7_75t_SL g1889 ( 
.A1(n_1555),
.A2(n_846),
.B1(n_1465),
.B2(n_872),
.C(n_843),
.Y(n_1889)
);

OAI21x1_ASAP7_75t_L g1890 ( 
.A1(n_1717),
.A2(n_1684),
.B(n_1436),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1629),
.B(n_1208),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1555),
.A2(n_1208),
.B1(n_1223),
.B2(n_1132),
.Y(n_1892)
);

OAI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1583),
.A2(n_1132),
.B1(n_872),
.B2(n_843),
.C(n_840),
.Y(n_1893)
);

OAI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1662),
.A2(n_701),
.B1(n_1208),
.B2(n_846),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1555),
.A2(n_1208),
.B1(n_1223),
.B2(n_1132),
.Y(n_1895)
);

BUFx12f_ASAP7_75t_L g1896 ( 
.A(n_1563),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1555),
.A2(n_1208),
.B1(n_1223),
.B2(n_1132),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1816),
.Y(n_1898)
);

NOR2x1_ASAP7_75t_SL g1899 ( 
.A(n_1859),
.B(n_1812),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1808),
.B(n_1811),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1817),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1838),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1827),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1767),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1781),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1806),
.B(n_1746),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1800),
.Y(n_1907)
);

INVx2_ASAP7_75t_SL g1908 ( 
.A(n_1859),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1819),
.B(n_1768),
.Y(n_1909)
);

OR2x2_ASAP7_75t_SL g1910 ( 
.A(n_1777),
.B(n_1825),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1864),
.B(n_1829),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1842),
.B(n_1836),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1842),
.B(n_1836),
.Y(n_1913)
);

NAND2x1p5_ASAP7_75t_L g1914 ( 
.A(n_1877),
.B(n_1769),
.Y(n_1914)
);

AND2x4_ASAP7_75t_SL g1915 ( 
.A(n_1859),
.B(n_1812),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1848),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1755),
.B(n_1837),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1755),
.B(n_1824),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1789),
.B(n_1792),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1762),
.B(n_1813),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1790),
.Y(n_1921)
);

INVxp67_ASAP7_75t_L g1922 ( 
.A(n_1844),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1812),
.B(n_1854),
.Y(n_1923)
);

CKINVDCx20_ASAP7_75t_R g1924 ( 
.A(n_1763),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1810),
.B(n_1799),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1810),
.B(n_1799),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1890),
.B(n_1756),
.Y(n_1927)
);

BUFx3_ASAP7_75t_L g1928 ( 
.A(n_1879),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1863),
.B(n_1860),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1799),
.B(n_1830),
.Y(n_1930)
);

INVx2_ASAP7_75t_SL g1931 ( 
.A(n_1857),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1780),
.B(n_1880),
.Y(n_1932)
);

INVxp67_ASAP7_75t_SL g1933 ( 
.A(n_1871),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1743),
.B(n_1745),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1834),
.Y(n_1935)
);

OR2x6_ASAP7_75t_L g1936 ( 
.A(n_1764),
.B(n_1759),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1743),
.B(n_1831),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1852),
.B(n_1850),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1754),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1839),
.B(n_1751),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1856),
.B(n_1889),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1751),
.B(n_1832),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1814),
.B(n_1750),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1750),
.B(n_1752),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1761),
.B(n_1835),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1845),
.A2(n_1897),
.B1(n_1883),
.B2(n_1892),
.Y(n_1946)
);

INVx2_ASAP7_75t_SL g1947 ( 
.A(n_1815),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1835),
.B(n_1747),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1840),
.B(n_1872),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1749),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1757),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1840),
.B(n_1872),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_SL g1953 ( 
.A(n_1893),
.B(n_1766),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1826),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1884),
.A2(n_1874),
.B1(n_1858),
.B2(n_1897),
.Y(n_1955)
);

NOR2x1_ASAP7_75t_L g1956 ( 
.A(n_1788),
.B(n_1803),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1843),
.B(n_1853),
.Y(n_1957)
);

HB1xp67_ASAP7_75t_L g1958 ( 
.A(n_1803),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1862),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1822),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1865),
.B(n_1868),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1891),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1791),
.B(n_1822),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1791),
.B(n_1845),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1821),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1849),
.B(n_1861),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1796),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1879),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1849),
.B(n_1861),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1883),
.B(n_1886),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1793),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1833),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1886),
.A2(n_1892),
.B1(n_1895),
.B2(n_1771),
.Y(n_1973)
);

OR2x6_ASAP7_75t_L g1974 ( 
.A(n_1809),
.B(n_1766),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1847),
.Y(n_1975)
);

INVxp67_ASAP7_75t_L g1976 ( 
.A(n_1818),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1823),
.B(n_1778),
.Y(n_1977)
);

BUFx3_ASAP7_75t_L g1978 ( 
.A(n_1879),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1820),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1895),
.B(n_1776),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1744),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1879),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1765),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1887),
.Y(n_1984)
);

OAI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1953),
.A2(n_1748),
.B1(n_1894),
.B2(n_1869),
.Y(n_1985)
);

NAND4xp25_ASAP7_75t_SL g1986 ( 
.A(n_1955),
.B(n_1851),
.C(n_1866),
.D(n_1870),
.Y(n_1986)
);

NAND4xp25_ASAP7_75t_L g1987 ( 
.A(n_1941),
.B(n_1875),
.C(n_1776),
.D(n_1770),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1898),
.Y(n_1988)
);

A2O1A1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1941),
.A2(n_1772),
.B(n_1774),
.C(n_1770),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1921),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1898),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_1931),
.Y(n_1992)
);

OAI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1946),
.A2(n_1888),
.B1(n_1885),
.B2(n_1876),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1901),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1929),
.A2(n_1753),
.B(n_1775),
.Y(n_1995)
);

OAI221xp5_ASAP7_75t_SL g1996 ( 
.A1(n_1955),
.A2(n_1973),
.B1(n_1946),
.B2(n_1938),
.C(n_1894),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1906),
.B(n_1855),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1901),
.Y(n_1998)
);

NOR3xp33_ASAP7_75t_L g1999 ( 
.A(n_1929),
.B(n_1876),
.C(n_1869),
.Y(n_1999)
);

OAI221xp5_ASAP7_75t_L g2000 ( 
.A1(n_1953),
.A2(n_1785),
.B1(n_1787),
.B2(n_1798),
.C(n_1801),
.Y(n_2000)
);

AOI221xp5_ASAP7_75t_L g2001 ( 
.A1(n_1938),
.A2(n_1841),
.B1(n_1779),
.B2(n_1878),
.C(n_1784),
.Y(n_2001)
);

AOI221xp5_ASAP7_75t_L g2002 ( 
.A1(n_1918),
.A2(n_1784),
.B1(n_1782),
.B2(n_1787),
.C(n_1795),
.Y(n_2002)
);

AOI221xp5_ASAP7_75t_L g2003 ( 
.A1(n_1918),
.A2(n_1765),
.B1(n_1786),
.B2(n_1804),
.C(n_1794),
.Y(n_2003)
);

NOR3xp33_ASAP7_75t_L g2004 ( 
.A(n_1980),
.B(n_1786),
.C(n_1807),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1924),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1906),
.B(n_1804),
.Y(n_2006)
);

OR2x2_ASAP7_75t_L g2007 ( 
.A(n_1932),
.B(n_1794),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1932),
.B(n_1881),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1984),
.B(n_1975),
.Y(n_2009)
);

OAI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1973),
.A2(n_1802),
.B1(n_1783),
.B2(n_1805),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_R g2011 ( 
.A(n_1924),
.B(n_1896),
.Y(n_2011)
);

OAI221xp5_ASAP7_75t_L g2012 ( 
.A1(n_1980),
.A2(n_1802),
.B1(n_1760),
.B2(n_1846),
.C(n_1758),
.Y(n_2012)
);

AND2x2_ASAP7_75t_SL g2013 ( 
.A(n_1915),
.B(n_1867),
.Y(n_2013)
);

AOI33xp33_ASAP7_75t_L g2014 ( 
.A1(n_1917),
.A2(n_1918),
.A3(n_1930),
.B1(n_1981),
.B2(n_1926),
.B3(n_1925),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1904),
.Y(n_2015)
);

AND2x4_ASAP7_75t_L g2016 ( 
.A(n_1908),
.B(n_1783),
.Y(n_2016)
);

AOI33xp33_ASAP7_75t_L g2017 ( 
.A1(n_1917),
.A2(n_1881),
.A3(n_1828),
.B1(n_1797),
.B2(n_1773),
.B3(n_1873),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1904),
.Y(n_2018)
);

NAND4xp25_ASAP7_75t_SL g2019 ( 
.A(n_1956),
.B(n_1881),
.C(n_1797),
.D(n_1882),
.Y(n_2019)
);

INVx3_ASAP7_75t_L g2020 ( 
.A(n_1928),
.Y(n_2020)
);

OAI33xp33_ASAP7_75t_L g2021 ( 
.A1(n_1981),
.A2(n_1797),
.A3(n_1760),
.B1(n_1758),
.B2(n_1846),
.B3(n_1867),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1979),
.B(n_1951),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1905),
.Y(n_2023)
);

NAND3xp33_ASAP7_75t_L g2024 ( 
.A(n_1919),
.B(n_1943),
.C(n_1967),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1905),
.Y(n_2025)
);

AO21x2_ASAP7_75t_L g2026 ( 
.A1(n_1916),
.A2(n_1927),
.B(n_1963),
.Y(n_2026)
);

AOI211xp5_ASAP7_75t_L g2027 ( 
.A1(n_1919),
.A2(n_1930),
.B(n_1967),
.C(n_1943),
.Y(n_2027)
);

BUFx3_ASAP7_75t_L g2028 ( 
.A(n_1947),
.Y(n_2028)
);

OAI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1966),
.A2(n_1969),
.B1(n_1970),
.B2(n_1974),
.Y(n_2029)
);

OAI33xp33_ASAP7_75t_L g2030 ( 
.A1(n_1935),
.A2(n_1964),
.A3(n_1922),
.B1(n_1969),
.B2(n_1970),
.B3(n_1966),
.Y(n_2030)
);

NAND2xp33_ASAP7_75t_R g2031 ( 
.A(n_1930),
.B(n_1974),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1959),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1974),
.A2(n_1964),
.B1(n_1956),
.B2(n_1910),
.Y(n_2033)
);

OAI211xp5_ASAP7_75t_L g2034 ( 
.A1(n_1943),
.A2(n_1963),
.B(n_1919),
.C(n_1925),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_1908),
.B(n_1947),
.Y(n_2035)
);

OAI33xp33_ASAP7_75t_L g2036 ( 
.A1(n_1935),
.A2(n_1922),
.A3(n_1979),
.B1(n_1957),
.B2(n_1961),
.B3(n_1951),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1907),
.Y(n_2037)
);

BUFx10_ASAP7_75t_L g2038 ( 
.A(n_1965),
.Y(n_2038)
);

NAND4xp25_ASAP7_75t_L g2039 ( 
.A(n_1957),
.B(n_1961),
.C(n_1972),
.D(n_1952),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1959),
.B(n_1962),
.Y(n_2040)
);

NAND4xp25_ASAP7_75t_L g2041 ( 
.A(n_1957),
.B(n_1961),
.C(n_1972),
.D(n_1949),
.Y(n_2041)
);

OAI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1974),
.A2(n_1925),
.B1(n_1926),
.B2(n_1951),
.Y(n_2042)
);

OAI221xp5_ASAP7_75t_L g2043 ( 
.A1(n_1974),
.A2(n_1965),
.B1(n_1902),
.B2(n_1914),
.C(n_1960),
.Y(n_2043)
);

AOI21xp33_ASAP7_75t_SL g2044 ( 
.A1(n_1974),
.A2(n_1909),
.B(n_1977),
.Y(n_2044)
);

OA21x2_ASAP7_75t_L g2045 ( 
.A1(n_1916),
.A2(n_1983),
.B(n_1942),
.Y(n_2045)
);

NAND2xp33_ASAP7_75t_R g2046 ( 
.A(n_1974),
.B(n_1926),
.Y(n_2046)
);

NAND3xp33_ASAP7_75t_L g2047 ( 
.A(n_1944),
.B(n_1940),
.C(n_1960),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1947),
.B(n_1915),
.Y(n_2048)
);

BUFx2_ASAP7_75t_L g2049 ( 
.A(n_1928),
.Y(n_2049)
);

NAND3xp33_ASAP7_75t_SL g2050 ( 
.A(n_1949),
.B(n_1952),
.C(n_1934),
.Y(n_2050)
);

INVxp67_ASAP7_75t_L g2051 ( 
.A(n_1958),
.Y(n_2051)
);

AOI21xp33_ASAP7_75t_L g2052 ( 
.A1(n_1944),
.A2(n_1940),
.B(n_1952),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2051),
.B(n_1917),
.Y(n_2053)
);

AND2x4_ASAP7_75t_L g2054 ( 
.A(n_2026),
.B(n_1923),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2045),
.B(n_2009),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_2045),
.B(n_2026),
.Y(n_2056)
);

NAND3xp33_ASAP7_75t_L g2057 ( 
.A(n_1995),
.B(n_1902),
.C(n_1949),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2051),
.B(n_1933),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1988),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1991),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1994),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1998),
.Y(n_2062)
);

NAND4xp25_ASAP7_75t_L g2063 ( 
.A(n_1987),
.B(n_1944),
.C(n_1940),
.D(n_1934),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2015),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2018),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1990),
.B(n_1933),
.Y(n_2066)
);

INVx1_ASAP7_75t_SL g2067 ( 
.A(n_2028),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2023),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2035),
.B(n_1911),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2025),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_2049),
.Y(n_2071)
);

INVx3_ASAP7_75t_L g2072 ( 
.A(n_2020),
.Y(n_2072)
);

AND2x4_ASAP7_75t_SL g2073 ( 
.A(n_2038),
.B(n_1958),
.Y(n_2073)
);

INVxp67_ASAP7_75t_SL g2074 ( 
.A(n_1990),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_SL g2075 ( 
.A1(n_2034),
.A2(n_1934),
.B1(n_1900),
.B2(n_1937),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2037),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2035),
.B(n_1911),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2022),
.B(n_1912),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_2040),
.B(n_1920),
.Y(n_2079)
);

BUFx3_ASAP7_75t_L g2080 ( 
.A(n_2038),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2050),
.B(n_1920),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2032),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2050),
.B(n_1920),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2022),
.B(n_1912),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2008),
.B(n_1962),
.Y(n_2085)
);

INVx1_ASAP7_75t_SL g2086 ( 
.A(n_1992),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2048),
.B(n_1913),
.Y(n_2087)
);

INVx3_ASAP7_75t_L g2088 ( 
.A(n_2013),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2006),
.B(n_1913),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2007),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2047),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2013),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2052),
.B(n_1997),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2014),
.B(n_1903),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2039),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2044),
.B(n_1913),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2016),
.B(n_1948),
.Y(n_2097)
);

OR2x2_ASAP7_75t_L g2098 ( 
.A(n_2041),
.B(n_1983),
.Y(n_2098)
);

INVx1_ASAP7_75t_SL g2099 ( 
.A(n_2016),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2033),
.B(n_1948),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2024),
.Y(n_2101)
);

AOI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_1999),
.A2(n_1950),
.B1(n_1937),
.B2(n_1900),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2059),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2101),
.B(n_2027),
.Y(n_2104)
);

HB1xp67_ASAP7_75t_L g2105 ( 
.A(n_2090),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2059),
.Y(n_2106)
);

OR2x2_ASAP7_75t_L g2107 ( 
.A(n_2081),
.B(n_1910),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2060),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2060),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2061),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2061),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2090),
.B(n_1899),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2081),
.B(n_1910),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2101),
.B(n_1976),
.Y(n_2114)
);

BUFx3_ASAP7_75t_L g2115 ( 
.A(n_2080),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2062),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_2056),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2090),
.B(n_1899),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_2081),
.B(n_1939),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2064),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2089),
.B(n_1976),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2064),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2089),
.B(n_1945),
.Y(n_2123)
);

NAND2x1p5_ASAP7_75t_L g2124 ( 
.A(n_2088),
.B(n_1923),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2083),
.B(n_2079),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2089),
.B(n_2042),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_2083),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2065),
.Y(n_2128)
);

OAI21xp33_ASAP7_75t_L g2129 ( 
.A1(n_2075),
.A2(n_1995),
.B(n_1989),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2068),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2068),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_SL g2132 ( 
.A(n_2057),
.B(n_2043),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2070),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2085),
.B(n_2042),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2087),
.B(n_1945),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2087),
.B(n_1945),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2085),
.B(n_2034),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2070),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2087),
.B(n_1923),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_2083),
.B(n_1939),
.Y(n_2140)
);

INVx2_ASAP7_75t_SL g2141 ( 
.A(n_2080),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2056),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2076),
.Y(n_2143)
);

NOR2xp33_ASAP7_75t_R g2144 ( 
.A(n_2080),
.B(n_2031),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2091),
.B(n_1971),
.Y(n_2145)
);

INVx1_ASAP7_75t_SL g2146 ( 
.A(n_2067),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_2063),
.B(n_2005),
.Y(n_2147)
);

OR2x6_ASAP7_75t_L g2148 ( 
.A(n_2057),
.B(n_1914),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2069),
.B(n_1923),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_2063),
.B(n_2029),
.Y(n_2150)
);

NAND3xp33_ASAP7_75t_L g2151 ( 
.A(n_2075),
.B(n_1999),
.C(n_2001),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2069),
.B(n_1948),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2069),
.B(n_1936),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2077),
.B(n_1936),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_2079),
.B(n_1939),
.Y(n_2155)
);

NOR2x1p5_ASAP7_75t_SL g2156 ( 
.A(n_2056),
.B(n_1916),
.Y(n_2156)
);

BUFx2_ASAP7_75t_L g2157 ( 
.A(n_2088),
.Y(n_2157)
);

INVx1_ASAP7_75t_SL g2158 ( 
.A(n_2146),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2137),
.B(n_2091),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2117),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2103),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2103),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2123),
.B(n_2095),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2106),
.Y(n_2164)
);

AOI21xp33_ASAP7_75t_L g2165 ( 
.A1(n_2129),
.A2(n_1993),
.B(n_1985),
.Y(n_2165)
);

BUFx2_ASAP7_75t_L g2166 ( 
.A(n_2144),
.Y(n_2166)
);

NOR3xp33_ASAP7_75t_L g2167 ( 
.A(n_2151),
.B(n_1996),
.C(n_1986),
.Y(n_2167)
);

AND2x4_ASAP7_75t_L g2168 ( 
.A(n_2157),
.B(n_2054),
.Y(n_2168)
);

HB1xp67_ASAP7_75t_L g2169 ( 
.A(n_2135),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2106),
.Y(n_2170)
);

OAI33xp33_ASAP7_75t_L g2171 ( 
.A1(n_2104),
.A2(n_1985),
.A3(n_2053),
.B1(n_2095),
.B2(n_2094),
.B3(n_2098),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2108),
.Y(n_2172)
);

INVxp67_ASAP7_75t_L g2173 ( 
.A(n_2132),
.Y(n_2173)
);

INVx1_ASAP7_75t_SL g2174 ( 
.A(n_2119),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2123),
.B(n_2053),
.Y(n_2175)
);

BUFx3_ASAP7_75t_L g2176 ( 
.A(n_2115),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2119),
.B(n_2098),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2157),
.B(n_2054),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2124),
.B(n_2054),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2124),
.B(n_2054),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2124),
.B(n_2054),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2153),
.B(n_2055),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2153),
.B(n_2055),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2154),
.B(n_2055),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2108),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2117),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2154),
.B(n_2127),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2109),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2149),
.B(n_2096),
.Y(n_2189)
);

OAI33xp33_ASAP7_75t_L g2190 ( 
.A1(n_2140),
.A2(n_2094),
.A3(n_2098),
.B1(n_2058),
.B2(n_2066),
.B3(n_2093),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2149),
.B(n_2096),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2134),
.B(n_2078),
.Y(n_2192)
);

INVx3_ASAP7_75t_SL g2193 ( 
.A(n_2141),
.Y(n_2193)
);

CKINVDCx20_ASAP7_75t_R g2194 ( 
.A(n_2147),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2142),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2109),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2112),
.B(n_2096),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2140),
.B(n_2078),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2112),
.B(n_2077),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2126),
.B(n_2078),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2118),
.B(n_2077),
.Y(n_2201)
);

HB1xp67_ASAP7_75t_L g2202 ( 
.A(n_2135),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2110),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2136),
.B(n_2084),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2110),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2142),
.Y(n_2206)
);

INVx1_ASAP7_75t_SL g2207 ( 
.A(n_2115),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2116),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2116),
.Y(n_2209)
);

OAI31xp33_ASAP7_75t_L g2210 ( 
.A1(n_2150),
.A2(n_1996),
.A3(n_2000),
.B(n_2019),
.Y(n_2210)
);

BUFx2_ASAP7_75t_L g2211 ( 
.A(n_2141),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2120),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2120),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2161),
.Y(n_2214)
);

OAI322xp33_ASAP7_75t_L g2215 ( 
.A1(n_2173),
.A2(n_2113),
.A3(n_2107),
.B1(n_2125),
.B2(n_2155),
.C1(n_2114),
.C2(n_2093),
.Y(n_2215)
);

AOI221xp5_ASAP7_75t_L g2216 ( 
.A1(n_2167),
.A2(n_2030),
.B1(n_2102),
.B2(n_2036),
.C(n_2002),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2166),
.B(n_2136),
.Y(n_2217)
);

INVx1_ASAP7_75t_SL g2218 ( 
.A(n_2158),
.Y(n_2218)
);

NAND4xp25_ASAP7_75t_L g2219 ( 
.A(n_2167),
.B(n_2165),
.C(n_2173),
.D(n_2210),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2163),
.B(n_2107),
.Y(n_2220)
);

OAI21xp33_ASAP7_75t_L g2221 ( 
.A1(n_2159),
.A2(n_2148),
.B(n_2113),
.Y(n_2221)
);

AOI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_2171),
.A2(n_2166),
.B1(n_2194),
.B2(n_2158),
.Y(n_2222)
);

INVxp67_ASAP7_75t_L g2223 ( 
.A(n_2176),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2159),
.B(n_2152),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_L g2225 ( 
.A(n_2171),
.B(n_2121),
.Y(n_2225)
);

AOI22xp33_ASAP7_75t_SL g2226 ( 
.A1(n_2210),
.A2(n_2148),
.B1(n_2100),
.B2(n_2031),
.Y(n_2226)
);

INVx2_ASAP7_75t_SL g2227 ( 
.A(n_2176),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2161),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2187),
.B(n_2152),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2187),
.B(n_2139),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2162),
.Y(n_2231)
);

INVxp67_ASAP7_75t_L g2232 ( 
.A(n_2211),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2162),
.Y(n_2233)
);

OAI321xp33_ASAP7_75t_L g2234 ( 
.A1(n_2163),
.A2(n_2148),
.A3(n_2012),
.B1(n_2125),
.B2(n_2100),
.C(n_2003),
.Y(n_2234)
);

OAI221xp5_ASAP7_75t_L g2235 ( 
.A1(n_2165),
.A2(n_2148),
.B1(n_2155),
.B2(n_2145),
.C(n_2004),
.Y(n_2235)
);

OR2x2_ASAP7_75t_L g2236 ( 
.A(n_2200),
.B(n_2192),
.Y(n_2236)
);

OAI32xp33_ASAP7_75t_L g2237 ( 
.A1(n_2207),
.A2(n_2046),
.A3(n_2100),
.B1(n_2088),
.B2(n_2004),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2207),
.B(n_2084),
.Y(n_2238)
);

O2A1O1Ixp5_ASAP7_75t_L g2239 ( 
.A1(n_2190),
.A2(n_2030),
.B(n_2036),
.C(n_2118),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2164),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2164),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2170),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2170),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2176),
.B(n_2084),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2211),
.B(n_2088),
.Y(n_2245)
);

OAI222xp33_ASAP7_75t_L g2246 ( 
.A1(n_2174),
.A2(n_2010),
.B1(n_2105),
.B2(n_1900),
.C1(n_1977),
.C2(n_1914),
.Y(n_2246)
);

OAI221xp5_ASAP7_75t_L g2247 ( 
.A1(n_2193),
.A2(n_2088),
.B1(n_2046),
.B2(n_2092),
.C(n_2082),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2172),
.Y(n_2248)
);

AOI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2190),
.A2(n_2092),
.B1(n_1937),
.B2(n_2097),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2172),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2192),
.B(n_2097),
.Y(n_2251)
);

OAI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_2193),
.A2(n_2092),
.B1(n_2073),
.B2(n_2082),
.Y(n_2252)
);

OAI221xp5_ASAP7_75t_SL g2253 ( 
.A1(n_2177),
.A2(n_2017),
.B1(n_1939),
.B2(n_1950),
.C(n_1954),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2200),
.B(n_2097),
.Y(n_2254)
);

INVx4_ASAP7_75t_L g2255 ( 
.A(n_2193),
.Y(n_2255)
);

INVxp67_ASAP7_75t_L g2256 ( 
.A(n_2217),
.Y(n_2256)
);

INVx1_ASAP7_75t_SL g2257 ( 
.A(n_2218),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2229),
.B(n_2199),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2214),
.Y(n_2259)
);

OAI21xp33_ASAP7_75t_L g2260 ( 
.A1(n_2226),
.A2(n_2187),
.B(n_2177),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2228),
.Y(n_2261)
);

OAI21xp5_ASAP7_75t_L g2262 ( 
.A1(n_2226),
.A2(n_2174),
.B(n_2169),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2255),
.B(n_2199),
.Y(n_2263)
);

AOI22xp33_ASAP7_75t_SL g2264 ( 
.A1(n_2225),
.A2(n_2202),
.B1(n_2197),
.B2(n_2011),
.Y(n_2264)
);

XOR2x2_ASAP7_75t_L g2265 ( 
.A(n_2222),
.B(n_2011),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2255),
.B(n_2199),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2231),
.Y(n_2267)
);

BUFx2_ASAP7_75t_SL g2268 ( 
.A(n_2227),
.Y(n_2268)
);

OAI221xp5_ASAP7_75t_SL g2269 ( 
.A1(n_2219),
.A2(n_2178),
.B1(n_2175),
.B2(n_2198),
.C(n_2204),
.Y(n_2269)
);

OR2x6_ASAP7_75t_L g2270 ( 
.A(n_2223),
.B(n_2168),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2233),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2216),
.B(n_2197),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2240),
.Y(n_2273)
);

NAND4xp25_ASAP7_75t_SL g2274 ( 
.A(n_2216),
.B(n_2197),
.C(n_2175),
.D(n_2198),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2230),
.B(n_2201),
.Y(n_2275)
);

OAI21xp5_ASAP7_75t_L g2276 ( 
.A1(n_2234),
.A2(n_2213),
.B(n_2212),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2241),
.Y(n_2277)
);

AOI21xp5_ASAP7_75t_L g2278 ( 
.A1(n_2237),
.A2(n_2204),
.B(n_2212),
.Y(n_2278)
);

INVx2_ASAP7_75t_SL g2279 ( 
.A(n_2245),
.Y(n_2279)
);

AOI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_2221),
.A2(n_2168),
.B1(n_2191),
.B2(n_2189),
.Y(n_2280)
);

NOR2xp33_ASAP7_75t_L g2281 ( 
.A(n_2215),
.B(n_2201),
.Y(n_2281)
);

OAI21xp5_ASAP7_75t_L g2282 ( 
.A1(n_2239),
.A2(n_2213),
.B(n_2185),
.Y(n_2282)
);

OAI221xp5_ASAP7_75t_L g2283 ( 
.A1(n_2253),
.A2(n_2178),
.B1(n_2208),
.B2(n_2188),
.C(n_2205),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2232),
.B(n_2189),
.Y(n_2284)
);

AOI211x1_ASAP7_75t_L g2285 ( 
.A1(n_2246),
.A2(n_2179),
.B(n_2180),
.C(n_2181),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2242),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2257),
.B(n_2232),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2264),
.B(n_2244),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2268),
.Y(n_2289)
);

BUFx2_ASAP7_75t_L g2290 ( 
.A(n_2270),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2284),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2270),
.Y(n_2292)
);

OAI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_2260),
.A2(n_2239),
.B(n_2246),
.Y(n_2293)
);

INVx1_ASAP7_75t_SL g2294 ( 
.A(n_2263),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2259),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2263),
.B(n_2245),
.Y(n_2296)
);

AOI211x1_ASAP7_75t_SL g2297 ( 
.A1(n_2276),
.A2(n_2252),
.B(n_2224),
.C(n_2238),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2270),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2261),
.Y(n_2299)
);

AOI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_2265),
.A2(n_2272),
.B1(n_2274),
.B2(n_2281),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2256),
.B(n_2236),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2266),
.B(n_2201),
.Y(n_2302)
);

A2O1A1Ixp33_ASAP7_75t_L g2303 ( 
.A1(n_2281),
.A2(n_2253),
.B(n_2235),
.C(n_2249),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2267),
.Y(n_2304)
);

NAND2x1p5_ASAP7_75t_L g2305 ( 
.A(n_2266),
.B(n_2243),
.Y(n_2305)
);

BUFx2_ASAP7_75t_L g2306 ( 
.A(n_2270),
.Y(n_2306)
);

AND2x2_ASAP7_75t_SL g2307 ( 
.A(n_2265),
.B(n_2220),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2271),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2279),
.B(n_2254),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2273),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_2289),
.B(n_2262),
.Y(n_2311)
);

INVx2_ASAP7_75t_SL g2312 ( 
.A(n_2302),
.Y(n_2312)
);

AOI21xp5_ASAP7_75t_L g2313 ( 
.A1(n_2293),
.A2(n_2282),
.B(n_2278),
.Y(n_2313)
);

NOR3xp33_ASAP7_75t_L g2314 ( 
.A(n_2287),
.B(n_2269),
.C(n_2279),
.Y(n_2314)
);

AOI211xp5_ASAP7_75t_L g2315 ( 
.A1(n_2303),
.A2(n_2283),
.B(n_2247),
.C(n_2286),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2305),
.Y(n_2316)
);

O2A1O1Ixp33_ASAP7_75t_L g2317 ( 
.A1(n_2290),
.A2(n_2277),
.B(n_2248),
.C(n_2250),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2300),
.B(n_2258),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2305),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2296),
.B(n_2258),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2300),
.B(n_2280),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2305),
.Y(n_2322)
);

AOI22xp5_ASAP7_75t_L g2323 ( 
.A1(n_2307),
.A2(n_2275),
.B1(n_2251),
.B2(n_2168),
.Y(n_2323)
);

AOI22xp33_ASAP7_75t_SL g2324 ( 
.A1(n_2307),
.A2(n_2275),
.B1(n_2168),
.B2(n_2178),
.Y(n_2324)
);

AOI221xp5_ASAP7_75t_L g2325 ( 
.A1(n_2294),
.A2(n_2285),
.B1(n_2168),
.B2(n_2160),
.C(n_2206),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2320),
.B(n_2296),
.Y(n_2326)
);

A2O1A1Ixp33_ASAP7_75t_L g2327 ( 
.A1(n_2313),
.A2(n_2307),
.B(n_2297),
.C(n_2290),
.Y(n_2327)
);

OAI21xp5_ASAP7_75t_L g2328 ( 
.A1(n_2311),
.A2(n_2288),
.B(n_2306),
.Y(n_2328)
);

AOI321xp33_ASAP7_75t_L g2329 ( 
.A1(n_2321),
.A2(n_2291),
.A3(n_2301),
.B1(n_2292),
.B2(n_2298),
.C(n_2309),
.Y(n_2329)
);

AOI222xp33_ASAP7_75t_L g2330 ( 
.A1(n_2318),
.A2(n_2306),
.B1(n_2291),
.B2(n_2308),
.C1(n_2304),
.C2(n_2299),
.Y(n_2330)
);

OAI221xp5_ASAP7_75t_L g2331 ( 
.A1(n_2315),
.A2(n_2292),
.B1(n_2298),
.B2(n_2304),
.C(n_2299),
.Y(n_2331)
);

NAND5xp2_ASAP7_75t_L g2332 ( 
.A(n_2314),
.B(n_2302),
.C(n_2308),
.D(n_2310),
.E(n_2295),
.Y(n_2332)
);

OAI211xp5_ASAP7_75t_L g2333 ( 
.A1(n_2318),
.A2(n_2310),
.B(n_2295),
.C(n_2160),
.Y(n_2333)
);

OAI211xp5_ASAP7_75t_L g2334 ( 
.A1(n_2324),
.A2(n_2160),
.B(n_2195),
.C(n_2206),
.Y(n_2334)
);

OAI221xp5_ASAP7_75t_L g2335 ( 
.A1(n_2323),
.A2(n_2195),
.B1(n_2186),
.B2(n_2206),
.C(n_2181),
.Y(n_2335)
);

A2O1A1Ixp33_ASAP7_75t_L g2336 ( 
.A1(n_2325),
.A2(n_2156),
.B(n_2073),
.C(n_2179),
.Y(n_2336)
);

AOI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2317),
.A2(n_2322),
.B(n_2319),
.Y(n_2337)
);

AOI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_2312),
.A2(n_2209),
.B1(n_2185),
.B2(n_2208),
.Y(n_2338)
);

INVx1_ASAP7_75t_SL g2339 ( 
.A(n_2326),
.Y(n_2339)
);

AOI22xp5_ASAP7_75t_L g2340 ( 
.A1(n_2328),
.A2(n_2316),
.B1(n_2186),
.B2(n_2195),
.Y(n_2340)
);

NOR2x1p5_ASAP7_75t_L g2341 ( 
.A(n_2329),
.B(n_2186),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2330),
.B(n_2327),
.Y(n_2342)
);

NOR2xp67_ASAP7_75t_L g2343 ( 
.A(n_2333),
.B(n_2188),
.Y(n_2343)
);

AOI31xp33_ASAP7_75t_L g2344 ( 
.A1(n_2327),
.A2(n_2180),
.A3(n_2181),
.B(n_2179),
.Y(n_2344)
);

AOI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_2331),
.A2(n_2180),
.B1(n_2191),
.B2(n_2189),
.Y(n_2345)
);

AOI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_2335),
.A2(n_2191),
.B1(n_2205),
.B2(n_2203),
.Y(n_2346)
);

A2O1A1Ixp33_ASAP7_75t_L g2347 ( 
.A1(n_2337),
.A2(n_2156),
.B(n_2073),
.C(n_2196),
.Y(n_2347)
);

NAND3xp33_ASAP7_75t_L g2348 ( 
.A(n_2342),
.B(n_2340),
.C(n_2347),
.Y(n_2348)
);

NOR3xp33_ASAP7_75t_L g2349 ( 
.A(n_2339),
.B(n_2332),
.C(n_2344),
.Y(n_2349)
);

AOI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_2343),
.A2(n_2336),
.B(n_2334),
.Y(n_2350)
);

AND3x2_ASAP7_75t_L g2351 ( 
.A(n_2341),
.B(n_2071),
.C(n_2209),
.Y(n_2351)
);

OAI22xp33_ASAP7_75t_SL g2352 ( 
.A1(n_2345),
.A2(n_2338),
.B1(n_2203),
.B2(n_2196),
.Y(n_2352)
);

XNOR2xp5_ASAP7_75t_L g2353 ( 
.A(n_2346),
.B(n_1928),
.Y(n_2353)
);

NAND2x1p5_ASAP7_75t_L g2354 ( 
.A(n_2339),
.B(n_1928),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2339),
.B(n_2182),
.Y(n_2355)
);

NOR2x1p5_ASAP7_75t_L g2356 ( 
.A(n_2342),
.B(n_1968),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2354),
.Y(n_2357)
);

NAND4xp25_ASAP7_75t_L g2358 ( 
.A(n_2349),
.B(n_2348),
.C(n_2350),
.D(n_2355),
.Y(n_2358)
);

NOR3xp33_ASAP7_75t_SL g2359 ( 
.A(n_2353),
.B(n_2021),
.C(n_2058),
.Y(n_2359)
);

OAI211xp5_ASAP7_75t_SL g2360 ( 
.A1(n_2356),
.A2(n_2082),
.B(n_2067),
.C(n_2099),
.Y(n_2360)
);

NAND3xp33_ASAP7_75t_SL g2361 ( 
.A(n_2351),
.B(n_2184),
.C(n_2183),
.Y(n_2361)
);

AO22x2_ASAP7_75t_L g2362 ( 
.A1(n_2352),
.A2(n_2184),
.B1(n_2183),
.B2(n_2182),
.Y(n_2362)
);

NAND4xp25_ASAP7_75t_L g2363 ( 
.A(n_2358),
.B(n_2360),
.C(n_2361),
.D(n_2357),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2362),
.Y(n_2364)
);

NOR3xp33_ASAP7_75t_L g2365 ( 
.A(n_2359),
.B(n_2021),
.C(n_2183),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2357),
.B(n_2182),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2364),
.B(n_2184),
.Y(n_2367)
);

HB1xp67_ASAP7_75t_L g2368 ( 
.A(n_2367),
.Y(n_2368)
);

BUFx12f_ASAP7_75t_L g2369 ( 
.A(n_2368),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2368),
.Y(n_2370)
);

XNOR2xp5_ASAP7_75t_L g2371 ( 
.A(n_2370),
.B(n_2363),
.Y(n_2371)
);

OAI222xp33_ASAP7_75t_L g2372 ( 
.A1(n_2370),
.A2(n_2366),
.B1(n_2365),
.B2(n_2086),
.C1(n_2143),
.C2(n_2122),
.Y(n_2372)
);

AOI22xp33_ASAP7_75t_L g2373 ( 
.A1(n_2371),
.A2(n_2369),
.B1(n_2072),
.B2(n_2071),
.Y(n_2373)
);

AOI222xp33_ASAP7_75t_L g2374 ( 
.A1(n_2372),
.A2(n_2143),
.B1(n_2122),
.B2(n_2128),
.C1(n_2130),
.C2(n_2131),
.Y(n_2374)
);

AOI322xp5_ASAP7_75t_L g2375 ( 
.A1(n_2373),
.A2(n_2086),
.A3(n_2074),
.B1(n_2099),
.B2(n_2139),
.C1(n_2130),
.C2(n_2128),
.Y(n_2375)
);

OAI221xp5_ASAP7_75t_L g2376 ( 
.A1(n_2375),
.A2(n_2374),
.B1(n_2111),
.B2(n_2138),
.C(n_2133),
.Y(n_2376)
);

AOI211xp5_ASAP7_75t_L g2377 ( 
.A1(n_2376),
.A2(n_1982),
.B(n_1968),
.C(n_1978),
.Y(n_2377)
);


endmodule