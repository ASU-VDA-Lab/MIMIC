module fake_jpeg_26198_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_30),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_42),
.B(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_24),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_24),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_17),
.B1(n_32),
.B2(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_25),
.B1(n_28),
.B2(n_20),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_52),
.B(n_54),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_28),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_55),
.C(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_32),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_19),
.B1(n_22),
.B2(n_33),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_68),
.Y(n_93)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_59),
.A2(n_63),
.B1(n_69),
.B2(n_74),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_56),
.A2(n_22),
.B1(n_36),
.B2(n_18),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_62),
.B(n_70),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_36),
.B1(n_31),
.B2(n_29),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_36),
.B1(n_32),
.B2(n_16),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_67),
.B1(n_79),
.B2(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_27),
.B1(n_18),
.B2(n_29),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_26),
.B1(n_30),
.B2(n_25),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_28),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_46),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_82),
.B(n_83),
.Y(n_91)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_42),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_16),
.B1(n_20),
.B2(n_3),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_43),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_12),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_15),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_110),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_89),
.A2(n_10),
.B(n_4),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_44),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_96),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_44),
.C(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_45),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_45),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_42),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_99),
.B(n_102),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_72),
.A2(n_47),
.B1(n_54),
.B2(n_20),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_79),
.B1(n_67),
.B2(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_112),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_59),
.B1(n_74),
.B2(n_64),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_0),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_0),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_72),
.B(n_86),
.C(n_87),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_142),
.B(n_90),
.Y(n_150)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_120),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_132),
.B1(n_111),
.B2(n_114),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_128),
.B1(n_140),
.B2(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_124),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_108),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_122),
.Y(n_143)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_61),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_80),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_81),
.B1(n_82),
.B2(n_65),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_133),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_84),
.B1(n_71),
.B2(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_9),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_9),
.Y(n_138)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_101),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_9),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_141),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_153),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_154),
.B1(n_140),
.B2(n_118),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_89),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_148),
.A2(n_149),
.B(n_150),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_90),
.B(n_93),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_112),
.B(n_92),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_151),
.A2(n_161),
.B(n_169),
.Y(n_192)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_117),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_158),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_91),
.B1(n_95),
.B2(n_113),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_102),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_157),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_95),
.C(n_5),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_12),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_119),
.B(n_135),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_5),
.C(n_6),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_166),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_124),
.C(n_125),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_119),
.A2(n_0),
.B(n_7),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_7),
.C(n_13),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_13),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_172),
.A2(n_174),
.B1(n_191),
.B2(n_194),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_160),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_176),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_142),
.B1(n_122),
.B2(n_126),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_175),
.A2(n_184),
.B(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_159),
.B(n_121),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

NAND2xp67_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_139),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_188),
.B(n_169),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_146),
.Y(n_189)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_156),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_205),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_161),
.C(n_151),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_209),
.C(n_192),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_174),
.B(n_175),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_204),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

OAI22x1_ASAP7_75t_SL g207 ( 
.A1(n_188),
.A2(n_144),
.B1(n_148),
.B2(n_150),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_171),
.C(n_158),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_182),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_212),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_165),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_217),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_195),
.C(n_185),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_173),
.C(n_180),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_220),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_203),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_179),
.C(n_164),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_222),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_212),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_183),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_228),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_189),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_153),
.B(n_204),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_208),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_207),
.B(n_202),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_225),
.B(n_218),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_213),
.B1(n_178),
.B2(n_176),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_237),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_198),
.C(n_209),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_201),
.C(n_211),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_238),
.B(n_240),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_215),
.A2(n_172),
.B1(n_186),
.B2(n_184),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_239),
.A2(n_190),
.B1(n_200),
.B2(n_155),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_206),
.CI(n_181),
.CON(n_240),
.SN(n_240)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_241),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_244),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_231),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_167),
.B(n_191),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_248),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_239),
.B(n_170),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_250),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_190),
.Y(n_250)
);

NOR3xp33_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_200),
.C(n_14),
.Y(n_251)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_251),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_232),
.C(n_237),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_238),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_258),
.B(n_243),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_252),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_262),
.A3(n_251),
.B1(n_244),
.B2(n_254),
.C1(n_240),
.C2(n_123),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_230),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_254),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_258),
.B(n_257),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_263),
.A2(n_236),
.B(n_256),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_264),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_240),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_133),
.Y(n_270)
);

OAI221xp5_ASAP7_75t_SL g271 ( 
.A1(n_270),
.A2(n_268),
.B1(n_14),
.B2(n_15),
.C(n_13),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_15),
.Y(n_272)
);


endmodule