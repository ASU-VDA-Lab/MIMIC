module real_jpeg_32348_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_704;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_338;
wire n_175;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_707;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_710;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_703;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_670;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_546;
wire n_285;
wire n_172;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_699;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_708;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_675;
wire n_179;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_709;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_702;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_706;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_705;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_0),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_0),
.Y(n_217)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_0),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_0),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_2),
.A2(n_20),
.B(n_21),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_3),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_3),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_3),
.A2(n_242),
.B1(n_263),
.B2(n_266),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_3),
.A2(n_242),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_3),
.A2(n_242),
.B1(n_411),
.B2(n_413),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_4),
.A2(n_166),
.B1(n_169),
.B2(n_170),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_4),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_4),
.A2(n_169),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_4),
.A2(n_169),
.B1(n_285),
.B2(n_287),
.Y(n_284)
);

AO22x1_ASAP7_75t_L g669 ( 
.A1(n_4),
.A2(n_169),
.B1(n_643),
.B2(n_670),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_5),
.A2(n_231),
.B1(n_232),
.B2(n_235),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_5),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_5),
.A2(n_166),
.B1(n_231),
.B2(n_366),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_5),
.A2(n_231),
.B1(n_461),
.B2(n_464),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_5),
.A2(n_231),
.B1(n_537),
.B2(n_541),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_6),
.A2(n_222),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_6),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_6),
.A2(n_226),
.B1(n_308),
.B2(n_313),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_6),
.A2(n_226),
.B1(n_390),
.B2(n_392),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_6),
.A2(n_226),
.B1(n_489),
.B2(n_493),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_7),
.B(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_7),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g418 ( 
.A(n_7),
.B(n_72),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_7),
.A2(n_384),
.B1(n_522),
.B2(n_525),
.Y(n_521)
);

OAI21xp33_ASAP7_75t_L g611 ( 
.A1(n_7),
.A2(n_203),
.B(n_546),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_9),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_9),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_10),
.Y(n_116)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_10),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_11),
.A2(n_299),
.B1(n_300),
.B2(n_303),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_11),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_11),
.A2(n_299),
.B1(n_397),
.B2(n_401),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_11),
.A2(n_299),
.B1(n_513),
.B2(n_517),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_SL g594 ( 
.A1(n_11),
.A2(n_299),
.B1(n_595),
.B2(n_598),
.Y(n_594)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_12),
.Y(n_119)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_12),
.Y(n_566)
);

CKINVDCx11_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_13),
.B(n_709),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_14),
.A2(n_57),
.B1(n_95),
.B2(n_99),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_14),
.A2(n_57),
.B1(n_195),
.B2(n_198),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g647 ( 
.A1(n_14),
.A2(n_57),
.B1(n_523),
.B2(n_648),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_15),
.Y(n_127)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_15),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_16),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_16),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_16),
.A2(n_136),
.B1(n_181),
.B2(n_184),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_16),
.A2(n_136),
.B1(n_350),
.B2(n_352),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_16),
.A2(n_136),
.B1(n_637),
.B2(n_643),
.Y(n_636)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_17),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_17),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_17),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_18),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_18),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_18),
.A2(n_75),
.B1(n_124),
.B2(n_128),
.Y(n_123)
);

AO22x1_ASAP7_75t_SL g210 ( 
.A1(n_18),
.A2(n_75),
.B1(n_120),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_18),
.A2(n_75),
.B1(n_677),
.B2(n_678),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_83),
.B(n_708),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_81),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_23),
.B(n_701),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_23),
.B(n_701),
.Y(n_707)
);

CKINVDCx16_ASAP7_75t_R g710 ( 
.A(n_23),
.Y(n_710)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_55),
.B1(n_70),
.B2(n_73),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g82 ( 
.A1(n_24),
.A2(n_70),
.B(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_24),
.Y(n_635)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2x1_ASAP7_75t_L g229 ( 
.A(n_25),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_25),
.B(n_221),
.Y(n_270)
);

AO22x1_ASAP7_75t_SL g297 ( 
.A1(n_25),
.A2(n_72),
.B1(n_230),
.B2(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_25),
.B(n_382),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_35),
.B2(n_38),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_27),
.Y(n_235)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_29),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_29),
.Y(n_644)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_34),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_34),
.Y(n_346)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_38),
.Y(n_342)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_41),
.Y(n_642)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_42),
.Y(n_268)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_45),
.Y(n_135)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_45),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_46),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_54),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_56),
.A2(n_71),
.B1(n_635),
.B2(n_669),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_62),
.Y(n_234)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_62),
.Y(n_302)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_66),
.Y(n_303)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_67),
.Y(n_265)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_67),
.Y(n_672)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_70),
.Y(n_668)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g261 ( 
.A(n_71),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_71),
.A2(n_262),
.B1(n_635),
.B2(n_636),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_72),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_72),
.B(n_298),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_78),
.Y(n_228)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g331 ( 
.A1(n_80),
.A2(n_332),
.A3(n_338),
.B1(n_341),
.B2(n_343),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_82),
.B(n_710),
.Y(n_709)
);

AO21x2_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_627),
.B(n_702),
.Y(n_83)
);

NAND2x1_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_444),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_376),
.B(n_440),
.Y(n_85)
);

NOR2xp67_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_322),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_87),
.A2(n_441),
.B(n_442),
.Y(n_440)
);

NOR3xp33_ASAP7_75t_L g445 ( 
.A(n_87),
.B(n_322),
.C(n_446),
.Y(n_445)
);

AOI21x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_271),
.B(n_274),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_251),
.Y(n_88)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_89),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_89),
.A2(n_251),
.B1(n_272),
.B2(n_273),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_176),
.B1(n_177),
.B2(n_250),
.Y(n_89)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_90),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_90),
.B(n_176),
.C(n_272),
.Y(n_630)
);

NAND2x1_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_175),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_131),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_92),
.B(n_131),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_101),
.B1(n_123),
.B2(n_130),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_94),
.A2(n_102),
.B1(n_186),
.B2(n_187),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_98),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_100),
.Y(n_183)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

AO22x1_ASAP7_75t_L g387 ( 
.A1(n_101),
.A2(n_130),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_101),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_101),
.A2(n_509),
.B1(n_510),
.B2(n_511),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_101),
.B(n_577),
.Y(n_576)
);

OA21x2_ASAP7_75t_L g652 ( 
.A1(n_101),
.A2(n_123),
.B(n_130),
.Y(n_652)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_102),
.A2(n_180),
.B1(n_186),
.B2(n_187),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_102),
.A2(n_180),
.B1(n_186),
.B2(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_102),
.A2(n_512),
.B1(n_551),
.B2(n_552),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_103)
);

BUFx4f_ASAP7_75t_SL g561 ( 
.A(n_104),
.Y(n_561)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_106),
.Y(n_145)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_106),
.Y(n_474)
);

OAI22x1_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_114),
.B1(n_117),
.B2(n_120),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_108),
.Y(n_572)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_113),
.Y(n_186)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_114),
.Y(n_351)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_115),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_116),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_116),
.Y(n_286)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_121),
.Y(n_545)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_122),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_122),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_125),
.Y(n_393)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_126),
.Y(n_518)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_127),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_127),
.Y(n_485)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_129),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_130),
.B(n_389),
.Y(n_468)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_130),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_142),
.B1(n_165),
.B2(n_173),
.Y(n_131)
);

AOI22x1_ASAP7_75t_L g237 ( 
.A1(n_132),
.A2(n_142),
.B1(n_238),
.B2(n_247),
.Y(n_237)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_141),
.Y(n_337)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_141),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_142),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_142),
.A2(n_173),
.B1(n_395),
.B2(n_396),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_142),
.B(n_307),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_142),
.A2(n_165),
.B1(n_173),
.B2(n_647),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_142),
.B(n_647),
.Y(n_680)
);

OA21x2_ASAP7_75t_SL g694 ( 
.A1(n_142),
.A2(n_173),
.B(n_695),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_156),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_143),
.Y(n_247)
);

AOI22x1_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_149),
.B2(n_152),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_146),
.A2(n_157),
.B1(n_160),
.B2(n_163),
.Y(n_156)
);

INVx5_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_148),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_154),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g467 ( 
.A(n_155),
.Y(n_467)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_163),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_168),
.Y(n_400)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_168),
.Y(n_525)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_174),
.A2(n_305),
.B1(n_306),
.B2(n_317),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_174),
.A2(n_407),
.B(n_408),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_R g549 ( 
.A(n_174),
.B(n_384),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_174),
.A2(n_675),
.B(n_680),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_175),
.A2(n_633),
.B1(n_654),
.B2(n_655),
.Y(n_632)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_175),
.Y(n_654)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_218),
.B(n_248),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_178),
.B(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_193),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_179),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_186),
.Y(n_509)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2x2_ASAP7_75t_L g372 ( 
.A(n_193),
.B(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_203),
.B1(n_209),
.B2(n_213),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_194),
.A2(n_203),
.B1(n_281),
.B2(n_283),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_196),
.Y(n_558)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_197),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_197),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_197),
.Y(n_570)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_203),
.B(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_203),
.A2(n_349),
.B1(n_410),
.B2(n_415),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_203),
.A2(n_536),
.B(n_546),
.Y(n_535)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_204),
.A2(n_284),
.B1(n_348),
.B2(n_355),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_204),
.B(n_488),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_204),
.A2(n_589),
.B1(n_592),
.B2(n_593),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_207),
.Y(n_416)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_SL g548 ( 
.A(n_208),
.Y(n_548)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_211),
.Y(n_412)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx2_ASAP7_75t_R g282 ( 
.A(n_216),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_217),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_236),
.Y(n_218)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_219),
.A2(n_236),
.B1(n_237),
.B2(n_249),
.Y(n_277)
);

NAND2x1_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_229),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_220),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_238),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_247),
.B(n_307),
.Y(n_370)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_259),
.Y(n_251)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_252),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_253),
.A2(n_258),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_253),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_257),
.Y(n_591)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_260),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_269),
.Y(n_260)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_266),
.Y(n_383)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_270),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_274),
.B(n_443),
.Y(n_442)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.C(n_318),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_276),
.B(n_319),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_278),
.B(n_375),
.Y(n_374)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_297),
.C(n_304),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_R g324 ( 
.A1(n_279),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_291),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_280),
.B(n_291),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx2_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_289),
.Y(n_495)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_290),
.Y(n_540)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_292),
.Y(n_388)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_294),
.Y(n_463)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_296),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_304),
.Y(n_325)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_311),
.Y(n_483)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_312),
.Y(n_650)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_317),
.A2(n_365),
.B(n_370),
.Y(n_364)
);

OA21x2_ASAP7_75t_L g520 ( 
.A1(n_317),
.A2(n_370),
.B(n_521),
.Y(n_520)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_320),
.A2(n_657),
.B(n_658),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_374),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_323),
.B(n_374),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.C(n_371),
.Y(n_323)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_325),
.A2(n_326),
.B1(n_372),
.B2(n_439),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_327),
.B(n_329),
.Y(n_437)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

MAJx2_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_360),
.C(n_363),
.Y(n_329)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_347),
.Y(n_330)
);

XOR2x2_ASAP7_75t_L g403 ( 
.A(n_331),
.B(n_347),
.Y(n_403)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_336),
.Y(n_344)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_341),
.Y(n_385)
);

NAND2xp33_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx2_ASAP7_75t_SL g597 ( 
.A(n_354),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_355),
.B(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_360),
.A2(n_361),
.B1(n_363),
.B2(n_364),
.Y(n_429)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_365),
.Y(n_395)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_366),
.Y(n_677)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_372),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_432),
.C(n_435),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_419),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_378),
.B(n_419),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_403),
.C(n_404),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_379),
.B(n_499),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_386),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_380),
.B(n_387),
.C(n_424),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_383),
.A2(n_384),
.B(n_385),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_384),
.B(n_472),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_384),
.B(n_482),
.C(n_484),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_384),
.B(n_574),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_384),
.A2(n_573),
.B(n_578),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_384),
.B(n_551),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_384),
.B(n_614),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_394),
.Y(n_386)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_389),
.Y(n_552)
);

INVx3_ASAP7_75t_SL g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_396),
.Y(n_407)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_402),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_403),
.A2(n_404),
.B1(n_405),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_403),
.Y(n_500)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.C(n_417),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_406),
.B(n_455),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_409),
.A2(n_417),
.B1(n_418),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_409),
.Y(n_456)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_426),
.B(n_430),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_431),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_422),
.B1(n_423),
.B2(n_425),
.Y(n_420)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_421),
.Y(n_425)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_423),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_425),
.Y(n_434)
);

MAJx2_ASAP7_75t_L g432 ( 
.A(n_426),
.B(n_433),
.C(n_434),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_427),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_432),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_436),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_436),
.A2(n_447),
.B(n_448),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_449),
.Y(n_444)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_501),
.B(n_625),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_498),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_452),
.B(n_626),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_457),
.C(n_469),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_454),
.B(n_527),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_457),
.A2(n_458),
.B1(n_469),
.B2(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_459),
.A2(n_460),
.B(n_468),
.Y(n_458)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_460),
.Y(n_510)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_468),
.B(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_469),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_486),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_470),
.B(n_486),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_475),
.B(n_481),
.Y(n_470)
);

INVx4_ASAP7_75t_SL g472 ( 
.A(n_473),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_484),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_496),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_487),
.A2(n_594),
.B(n_607),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_488),
.B(n_547),
.Y(n_546)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_498),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_529),
.B(n_624),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_526),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g624 ( 
.A(n_503),
.B(n_526),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_506),
.C(n_519),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_505),
.B(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_520),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_523),
.Y(n_679)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_584),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_531),
.A2(n_553),
.B(n_583),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_534),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_532),
.B(n_534),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_549),
.C(n_550),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_535),
.A2(n_580),
.B1(n_581),
.B2(n_582),
.Y(n_579)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_535),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_536),
.Y(n_592)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_539),
.Y(n_598)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_549),
.B(n_550),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_579),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_554),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_575),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_555),
.A2(n_575),
.B1(n_600),
.B2(n_601),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_555),
.Y(n_600)
);

AO221x1_ASAP7_75t_L g620 ( 
.A1(n_555),
.A2(n_575),
.B1(n_588),
.B2(n_600),
.C(n_601),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_556),
.A2(n_559),
.B(n_567),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_562),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_568),
.A2(n_571),
.B(n_573),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_575),
.Y(n_601)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_579),
.Y(n_622)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_580),
.Y(n_581)
);

NAND3xp33_ASAP7_75t_L g584 ( 
.A(n_583),
.B(n_585),
.C(n_621),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_586),
.A2(n_602),
.B(n_620),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_599),
.Y(n_587)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_589),
.Y(n_614)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_591),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_604),
.A2(n_610),
.B(n_619),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_605),
.B(n_606),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_605),
.B(n_606),
.Y(n_619)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_611),
.B(n_612),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_613),
.B(n_615),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_616),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_622),
.B(n_623),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g627 ( 
.A(n_628),
.B(n_686),
.C(n_700),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_629),
.B(n_659),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_630),
.B(n_631),
.Y(n_629)
);

NOR2xp67_ASAP7_75t_L g705 ( 
.A(n_630),
.B(n_631),
.Y(n_705)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_632),
.B(n_656),
.Y(n_631)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_633),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_633),
.Y(n_683)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_634),
.B(n_645),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_634),
.Y(n_662)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_634),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_635),
.A2(n_636),
.B1(n_668),
.B2(n_669),
.Y(n_667)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_639),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_641),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_642),
.Y(n_641)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_646),
.A2(n_651),
.B1(n_652),
.B2(n_653),
.Y(n_645)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_646),
.Y(n_653)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_649),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_651),
.A2(n_652),
.B1(n_674),
.B2(n_681),
.Y(n_673)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_652),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_652),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g661 ( 
.A(n_653),
.B(n_662),
.C(n_663),
.Y(n_661)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_654),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_656),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_659),
.A2(n_687),
.B(n_705),
.C(n_706),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_660),
.B(n_682),
.Y(n_659)
);

NOR2xp67_ASAP7_75t_L g706 ( 
.A(n_660),
.B(n_682),
.Y(n_706)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_661),
.B(n_664),
.Y(n_660)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_661),
.Y(n_699)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_663),
.Y(n_692)
);

XNOR2xp5_ASAP7_75t_L g664 ( 
.A(n_665),
.B(n_666),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g697 ( 
.A(n_665),
.B(n_698),
.C(n_699),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_666),
.Y(n_698)
);

XNOR2xp5_ASAP7_75t_L g666 ( 
.A(n_667),
.B(n_673),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_667),
.Y(n_690)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_671),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_672),
.Y(n_671)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_674),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_674),
.Y(n_691)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_676),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_676),
.Y(n_695)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_679),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g682 ( 
.A(n_683),
.B(n_684),
.C(n_685),
.Y(n_682)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_687),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_688),
.B(n_697),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_688),
.B(n_697),
.Y(n_703)
);

XNOR2xp5_ASAP7_75t_L g688 ( 
.A(n_689),
.B(n_693),
.Y(n_688)
);

MAJIxp5_ASAP7_75t_L g701 ( 
.A(n_689),
.B(n_694),
.C(n_696),
.Y(n_701)
);

MAJIxp5_ASAP7_75t_L g689 ( 
.A(n_690),
.B(n_691),
.C(n_692),
.Y(n_689)
);

XNOR2xp5_ASAP7_75t_L g693 ( 
.A(n_694),
.B(n_696),
.Y(n_693)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_700),
.A2(n_703),
.B(n_704),
.C(n_707),
.Y(n_702)
);


endmodule