module fake_jpeg_12035_n_657 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_657);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_657;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_68),
.Y(n_210)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_21),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_76),
.Y(n_132)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_74),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_77),
.Y(n_185)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx5_ASAP7_75t_SL g148 ( 
.A(n_79),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_34),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_80),
.B(n_81),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_83),
.Y(n_193)
);

INVx11_ASAP7_75t_SL g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_85),
.Y(n_204)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_88),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_89),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_8),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_90),
.B(n_91),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_34),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_30),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_101),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_94),
.Y(n_214)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_95),
.Y(n_201)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

BUFx4f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_100),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_37),
.B(n_8),
.Y(n_101)
);

BUFx16f_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g190 ( 
.A(n_102),
.Y(n_190)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_24),
.B(n_8),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_108),
.B(n_14),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_34),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_117),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

BUFx16f_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_24),
.B(n_7),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_49),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_122),
.Y(n_173)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_121),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_49),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_32),
.Y(n_124)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_53),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_127),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_28),
.B(n_6),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_49),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_35),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_32),
.Y(n_130)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx11_ASAP7_75t_L g262 ( 
.A(n_141),
.Y(n_262)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_150),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_SL g157 ( 
.A(n_111),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_157),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_92),
.B(n_58),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_158),
.B(n_160),
.Y(n_233)
);

AND2x4_ASAP7_75t_L g160 ( 
.A(n_68),
.B(n_35),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_169),
.B(n_177),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_123),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_170),
.B(n_192),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_123),
.Y(n_174)
);

HAxp5_ASAP7_75t_SL g227 ( 
.A(n_174),
.B(n_128),
.CON(n_227),
.SN(n_227)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_81),
.B(n_43),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_78),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_195),
.Y(n_235)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_75),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_187),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_107),
.B(n_36),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_69),
.Y(n_194)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_71),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_102),
.B(n_36),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_197),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_82),
.B(n_42),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_82),
.B(n_42),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_87),
.Y(n_199)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_96),
.Y(n_202)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_104),
.A2(n_53),
.B1(n_59),
.B2(n_46),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_67),
.B1(n_105),
.B2(n_99),
.Y(n_228)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_75),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g258 ( 
.A(n_208),
.Y(n_258)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_63),
.Y(n_211)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_128),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_54),
.Y(n_249)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_64),
.Y(n_216)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_216),
.Y(n_279)
);

BUFx4f_ASAP7_75t_SL g218 ( 
.A(n_157),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_218),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_144),
.A2(n_119),
.B1(n_113),
.B2(n_110),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_219),
.Y(n_319)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_134),
.A2(n_47),
.B(n_41),
.C(n_57),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_221),
.B(n_229),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_144),
.A2(n_126),
.B1(n_47),
.B2(n_41),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_222),
.A2(n_290),
.B1(n_195),
.B2(n_142),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_145),
.Y(n_223)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_223),
.Y(n_331)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_133),
.Y(n_225)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_225),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_160),
.A2(n_130),
.B1(n_124),
.B2(n_120),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_SL g309 ( 
.A1(n_226),
.A2(n_172),
.B(n_164),
.C(n_159),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_227),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_228),
.A2(n_185),
.B1(n_207),
.B2(n_165),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_143),
.B(n_154),
.Y(n_229)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_148),
.Y(n_231)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_151),
.B(n_54),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_232),
.B(n_244),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_175),
.A2(n_89),
.B1(n_65),
.B2(n_74),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_234),
.A2(n_238),
.B1(n_294),
.B2(n_139),
.Y(n_296)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_135),
.Y(n_236)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_236),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_139),
.A2(n_112),
.B1(n_94),
.B2(n_88),
.Y(n_238)
);

CKINVDCx12_ASAP7_75t_R g239 ( 
.A(n_182),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_239),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_145),
.Y(n_241)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_241),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_242),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_166),
.B(n_57),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_158),
.B(n_0),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_252),
.C(n_283),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_203),
.A2(n_85),
.B1(n_83),
.B2(n_77),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_246),
.A2(n_164),
.B1(n_172),
.B2(n_217),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_147),
.Y(n_247)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_147),
.Y(n_248)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_256),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_135),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_250),
.B(n_255),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_132),
.B(n_45),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_251),
.B(n_253),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_160),
.B(n_0),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_149),
.B(n_45),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_161),
.Y(n_254)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_254),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_131),
.B(n_60),
.Y(n_255)
);

CKINVDCx12_ASAP7_75t_R g256 ( 
.A(n_182),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_173),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_257),
.B(n_265),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_174),
.B(n_43),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_260),
.B(n_261),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_156),
.B(n_28),
.Y(n_261)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_184),
.Y(n_263)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_263),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_156),
.B(n_60),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_264),
.B(n_275),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_176),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_184),
.Y(n_266)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_184),
.Y(n_268)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_153),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_142),
.Y(n_270)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_210),
.Y(n_271)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_136),
.B(n_0),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_281),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_189),
.B(n_59),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_176),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_276),
.B(n_278),
.Y(n_317)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_210),
.Y(n_277)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_148),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_189),
.Y(n_280)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_280),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_140),
.B(n_0),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_162),
.B(n_186),
.C(n_180),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_188),
.Y(n_284)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_161),
.Y(n_285)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_285),
.Y(n_341)
);

BUFx12f_ASAP7_75t_L g286 ( 
.A(n_205),
.Y(n_286)
);

INVx11_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_167),
.Y(n_287)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_287),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_181),
.Y(n_288)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_191),
.A2(n_46),
.B1(n_44),
.B2(n_100),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_289),
.A2(n_163),
.B(n_207),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_137),
.A2(n_200),
.B1(n_138),
.B2(n_171),
.Y(n_290)
);

INVx3_ASAP7_75t_SL g292 ( 
.A(n_217),
.Y(n_292)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_155),
.B(n_44),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_293),
.B(n_165),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_159),
.A2(n_46),
.B1(n_44),
.B2(n_61),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_296),
.B(n_309),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_300),
.A2(n_345),
.B1(n_231),
.B2(n_242),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_301),
.A2(n_305),
.B1(n_342),
.B2(n_282),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_215),
.B1(n_201),
.B2(n_142),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_233),
.B(n_190),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_312),
.B(n_318),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_233),
.A2(n_168),
.B1(n_152),
.B2(n_214),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_316),
.A2(n_330),
.B1(n_352),
.B2(n_282),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_233),
.B(n_190),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_255),
.A2(n_214),
.B1(n_213),
.B2(n_209),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_320),
.A2(n_323),
.B1(n_334),
.B2(n_338),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_272),
.B(n_168),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_322),
.B(n_226),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_229),
.A2(n_213),
.B1(n_209),
.B2(n_204),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_252),
.A2(n_185),
.B1(n_181),
.B2(n_193),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_283),
.B(n_204),
.C(n_193),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_348),
.C(n_226),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_273),
.A2(n_243),
.B1(n_289),
.B2(n_281),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_294),
.A2(n_221),
.B1(n_232),
.B2(n_244),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_346),
.B(n_350),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_245),
.B(n_207),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_227),
.B(n_61),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_225),
.Y(n_351)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_351),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_252),
.A2(n_49),
.B1(n_61),
.B2(n_2),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_224),
.Y(n_355)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_355),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_317),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_356),
.B(n_361),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_358),
.A2(n_377),
.B1(n_327),
.B2(n_335),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_359),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_360),
.B(n_364),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_314),
.Y(n_361)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_362),
.Y(n_429)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_303),
.B(n_245),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_236),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_366),
.B(n_376),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_303),
.B(n_220),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_367),
.B(n_370),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_326),
.A2(n_271),
.B1(n_277),
.B2(n_226),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_368),
.A2(n_375),
.B(n_401),
.Y(n_412)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_297),
.Y(n_369)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_369),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_322),
.B(n_237),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_371),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_383),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_309),
.A2(n_287),
.B1(n_279),
.B2(n_267),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_374),
.A2(n_389),
.B1(n_400),
.B2(n_345),
.Y(n_406)
);

AOI32xp33_ASAP7_75t_L g375 ( 
.A1(n_353),
.A2(n_240),
.A3(n_291),
.B1(n_274),
.B2(n_258),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_328),
.Y(n_376)
);

INVx13_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_378),
.Y(n_403)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_313),
.Y(n_379)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_379),
.Y(n_414)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_381),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_224),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_332),
.B(n_230),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_388),
.Y(n_418)
);

AO22x1_ASAP7_75t_SL g386 ( 
.A1(n_300),
.A2(n_230),
.B1(n_259),
.B2(n_267),
.Y(n_386)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_386),
.Y(n_426)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_299),
.Y(n_387)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_387),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_307),
.B(n_235),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_319),
.A2(n_307),
.B1(n_318),
.B2(n_312),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_298),
.B(n_280),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_390),
.B(n_391),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_348),
.B(n_347),
.Y(n_391)
);

AND2x6_ASAP7_75t_L g392 ( 
.A(n_350),
.B(n_291),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_394),
.Y(n_423)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_297),
.Y(n_393)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_393),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_325),
.B(n_259),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_319),
.A2(n_333),
.B1(n_342),
.B2(n_335),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_395),
.A2(n_397),
.B1(n_402),
.B2(n_286),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_295),
.B(n_269),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_398),
.C(n_399),
.Y(n_421)
);

BUFx12_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_344),
.B(n_286),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_310),
.B(n_284),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_312),
.A2(n_279),
.B1(n_288),
.B2(n_241),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_306),
.B(n_0),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_339),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_406),
.A2(n_408),
.B1(n_432),
.B2(n_433),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_384),
.A2(n_318),
.B(n_321),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_407),
.A2(n_440),
.B(n_362),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_360),
.A2(n_330),
.B1(n_316),
.B2(n_352),
.Y(n_408)
);

OAI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_410),
.A2(n_426),
.B1(n_416),
.B2(n_427),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_368),
.A2(n_311),
.B(n_302),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_415),
.A2(n_417),
.B(n_419),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_365),
.A2(n_329),
.B1(n_341),
.B2(n_349),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_416),
.A2(n_425),
.B1(n_427),
.B2(n_400),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_365),
.A2(n_311),
.B(n_302),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_366),
.A2(n_274),
.B(n_262),
.Y(n_419)
);

AO21x2_ASAP7_75t_L g420 ( 
.A1(n_365),
.A2(n_262),
.B(n_313),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_420),
.B(n_386),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_377),
.A2(n_372),
.B1(n_385),
.B2(n_370),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_357),
.A2(n_341),
.B1(n_349),
.B2(n_331),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_389),
.A2(n_327),
.B(n_321),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_430),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_431),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_357),
.A2(n_248),
.B1(n_223),
.B2(n_247),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_374),
.A2(n_254),
.B1(n_285),
.B2(n_324),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_382),
.A2(n_308),
.B(n_343),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_434),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_382),
.A2(n_392),
.B(n_383),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_394),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_382),
.A2(n_266),
.B(n_268),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_367),
.A2(n_340),
.B1(n_324),
.B2(n_343),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_442),
.A2(n_369),
.B1(n_393),
.B2(n_379),
.Y(n_470)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_435),
.Y(n_443)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_443),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_413),
.B(n_388),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_447),
.B(n_460),
.Y(n_500)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_435),
.Y(n_448)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_448),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_391),
.C(n_364),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_449),
.B(n_452),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_423),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_451),
.B(n_478),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_418),
.B(n_373),
.C(n_380),
.Y(n_452)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_411),
.Y(n_454)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_454),
.Y(n_487)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_411),
.Y(n_455)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_455),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_308),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_456),
.B(n_461),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_428),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_457),
.B(n_459),
.Y(n_495)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_437),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_458),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_418),
.B(n_399),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_406),
.B(n_359),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_422),
.B(n_378),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_462),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_463),
.A2(n_477),
.B1(n_408),
.B2(n_432),
.Y(n_499)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_464),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_403),
.B(n_401),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g480 ( 
.A(n_465),
.Y(n_480)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_468),
.Y(n_485)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_436),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_469),
.B(n_470),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_425),
.B(n_397),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_471),
.B(n_475),
.Y(n_511)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_434),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_472),
.B(n_441),
.Y(n_497)
);

INVx13_ASAP7_75t_L g473 ( 
.A(n_403),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_473),
.Y(n_503)
);

INVx13_ASAP7_75t_L g474 ( 
.A(n_429),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_479),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_409),
.A2(n_381),
.B1(n_363),
.B2(n_386),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_476),
.A2(n_415),
.B(n_417),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_SL g478 ( 
.A(n_419),
.B(n_397),
.C(n_282),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_424),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_466),
.A2(n_420),
.B1(n_409),
.B2(n_426),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_484),
.A2(n_489),
.B1(n_498),
.B2(n_513),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_488),
.A2(n_446),
.B(n_458),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_466),
.A2(n_420),
.B1(n_410),
.B2(n_404),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_464),
.B(n_439),
.Y(n_494)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_494),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_497),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_450),
.A2(n_420),
.B1(n_404),
.B2(n_439),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_499),
.A2(n_445),
.B1(n_470),
.B2(n_453),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_452),
.B(n_430),
.Y(n_502)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_502),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_449),
.B(n_424),
.Y(n_505)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_505),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_454),
.B(n_420),
.Y(n_507)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_507),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_460),
.A2(n_433),
.B1(n_412),
.B2(n_407),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_508),
.A2(n_510),
.B1(n_514),
.B2(n_444),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_467),
.B(n_405),
.Y(n_509)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_509),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_460),
.A2(n_412),
.B1(n_405),
.B2(n_414),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_468),
.B(n_414),
.Y(n_512)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_512),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_444),
.A2(n_476),
.B1(n_475),
.B2(n_460),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_463),
.A2(n_421),
.B1(n_340),
.B2(n_440),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_501),
.Y(n_515)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_515),
.Y(n_550)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_491),
.Y(n_517)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_517),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_500),
.B(n_447),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_SL g549 ( 
.A(n_519),
.B(n_494),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_520),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_471),
.C(n_459),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_521),
.B(n_528),
.C(n_511),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_495),
.B(n_469),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_522),
.B(n_524),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_500),
.B(n_421),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_523),
.B(n_541),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_451),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_485),
.B(n_479),
.Y(n_526)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_526),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_527),
.A2(n_543),
.B1(n_492),
.B2(n_503),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_511),
.B(n_453),
.C(n_446),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_480),
.A2(n_445),
.B1(n_448),
.B2(n_443),
.Y(n_529)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_529),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_531),
.B(n_504),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_508),
.A2(n_462),
.B1(n_473),
.B2(n_474),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_532),
.B(n_533),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_499),
.A2(n_339),
.B1(n_336),
.B2(n_270),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_501),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_534),
.B(n_535),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_490),
.A2(n_258),
.B1(n_263),
.B2(n_165),
.Y(n_535)
);

BUFx5_ASAP7_75t_L g539 ( 
.A(n_491),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g559 ( 
.A(n_539),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_485),
.B(n_1),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_540),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_512),
.B(n_2),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_493),
.B(n_258),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_509),
.B(n_3),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_544),
.B(n_481),
.Y(n_564)
);

INVxp33_ASAP7_75t_SL g545 ( 
.A(n_498),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_545),
.A2(n_490),
.B1(n_514),
.B2(n_510),
.Y(n_546)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_546),
.Y(n_575)
);

MAJx2_ASAP7_75t_L g591 ( 
.A(n_547),
.B(n_568),
.C(n_570),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_521),
.B(n_511),
.C(n_504),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_548),
.B(n_554),
.C(n_557),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_549),
.B(n_553),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_SL g553 ( 
.A(n_519),
.B(n_482),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_524),
.B(n_504),
.C(n_482),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_536),
.A2(n_493),
.B1(n_488),
.B2(n_506),
.Y(n_555)
);

INVxp33_ASAP7_75t_L g588 ( 
.A(n_555),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_556),
.A2(n_542),
.B(n_538),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_523),
.B(n_513),
.Y(n_557)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_562),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_518),
.A2(n_506),
.B1(n_503),
.B2(n_492),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_563),
.B(n_564),
.Y(n_576)
);

FAx1_ASAP7_75t_SL g565 ( 
.A(n_528),
.B(n_489),
.CI(n_484),
.CON(n_565),
.SN(n_565)
);

FAx1_ASAP7_75t_SL g572 ( 
.A(n_565),
.B(n_536),
.CI(n_531),
.CON(n_572),
.SN(n_572)
);

XNOR2xp5_ASAP7_75t_SL g568 ( 
.A(n_522),
.B(n_520),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_525),
.B(n_487),
.C(n_507),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_572),
.B(n_574),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_558),
.A2(n_537),
.B1(n_542),
.B2(n_516),
.Y(n_573)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_573),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_564),
.B(n_526),
.Y(n_577)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_577),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_556),
.A2(n_532),
.B(n_530),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_578),
.A2(n_583),
.B(n_584),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_560),
.B(n_487),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_579),
.B(n_582),
.Y(n_602)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_551),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_581),
.B(n_589),
.Y(n_606)
);

NOR2xp67_ASAP7_75t_R g582 ( 
.A(n_554),
.B(n_540),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_556),
.A2(n_535),
.B(n_544),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_558),
.A2(n_517),
.B(n_486),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_567),
.B(n_541),
.Y(n_585)
);

NOR2xp67_ASAP7_75t_L g603 ( 
.A(n_585),
.B(n_561),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_SL g587 ( 
.A1(n_566),
.A2(n_496),
.B1(n_486),
.B2(n_481),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_587),
.B(n_593),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_565),
.A2(n_496),
.B1(n_491),
.B2(n_539),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_565),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_592),
.B(n_5),
.Y(n_610)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_550),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_586),
.A2(n_547),
.B(n_548),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_594),
.A2(n_600),
.B(n_605),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_586),
.B(n_568),
.C(n_570),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_596),
.B(n_607),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_552),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_599),
.B(n_608),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_578),
.A2(n_557),
.B(n_552),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_603),
.B(n_592),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_580),
.A2(n_571),
.B(n_569),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_591),
.B(n_553),
.C(n_549),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_590),
.B(n_561),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_588),
.B(n_559),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_610),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_580),
.A2(n_218),
.B(n_12),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_611),
.A2(n_581),
.B(n_583),
.Y(n_625)
);

MAJx2_ASAP7_75t_L g612 ( 
.A(n_602),
.B(n_607),
.C(n_597),
.Y(n_612)
);

AOI31xp67_ASAP7_75t_L g630 ( 
.A1(n_612),
.A2(n_620),
.A3(n_598),
.B(n_574),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_596),
.B(n_591),
.C(n_575),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_613),
.B(n_617),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_599),
.B(n_575),
.C(n_576),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_608),
.B(n_584),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_618),
.B(n_619),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_SL g619 ( 
.A(n_600),
.B(n_590),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_604),
.B(n_593),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_597),
.A2(n_582),
.B(n_579),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_621),
.A2(n_602),
.B(n_598),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_605),
.Y(n_622)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_622),
.Y(n_627)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_623),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_625),
.B(n_576),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_606),
.B(n_572),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_626),
.B(n_577),
.Y(n_635)
);

INVxp33_ASAP7_75t_L g628 ( 
.A(n_622),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_628),
.B(n_631),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_629),
.A2(n_612),
.B(n_573),
.Y(n_639)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_630),
.Y(n_638)
);

MAJx2_ASAP7_75t_L g634 ( 
.A(n_616),
.B(n_595),
.C(n_601),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_634),
.B(n_218),
.C(n_15),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_635),
.B(n_11),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_615),
.A2(n_611),
.B1(n_585),
.B2(n_572),
.Y(n_636)
);

AOI322xp5_ASAP7_75t_L g640 ( 
.A1(n_636),
.A2(n_619),
.A3(n_618),
.B1(n_614),
.B2(n_624),
.C1(n_610),
.C2(n_61),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_639),
.A2(n_642),
.B(n_17),
.Y(n_649)
);

OAI21x1_ASAP7_75t_SL g650 ( 
.A1(n_640),
.A2(n_643),
.B(n_11),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_633),
.A2(n_614),
.B1(n_14),
.B2(n_15),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_641),
.B(n_644),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_637),
.B(n_632),
.C(n_627),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_644),
.B(n_631),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_647),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_638),
.B(n_628),
.C(n_15),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_648),
.B(n_649),
.C(n_650),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_SL g653 ( 
.A(n_652),
.B(n_639),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_653),
.B(n_645),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_654),
.A2(n_646),
.B(n_642),
.Y(n_655)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_655),
.B(n_651),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_656),
.A2(n_11),
.B(n_15),
.Y(n_657)
);


endmodule