module fake_jpeg_29041_n_381 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_381);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_381;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_1),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_54),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_29),
.Y(n_102)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_60),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_59),
.Y(n_106)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_70),
.Y(n_99)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g107 ( 
.A(n_62),
.Y(n_107)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx2_ASAP7_75t_R g103 ( 
.A(n_66),
.Y(n_103)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_43),
.B1(n_24),
.B2(n_27),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_73),
.A2(n_55),
.B1(n_41),
.B2(n_33),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_31),
.B1(n_23),
.B2(n_22),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_76),
.A2(n_38),
.B1(n_31),
.B2(n_29),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_85),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_38),
.B1(n_24),
.B2(n_27),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_38),
.B1(n_66),
.B2(n_71),
.Y(n_109)
);

INVx2_ASAP7_75t_R g94 ( 
.A(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_97),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_35),
.B(n_37),
.Y(n_97)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_22),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_105),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_102),
.B(n_21),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_71),
.B(n_21),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_109),
.A2(n_41),
.B(n_90),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_110),
.B(n_1),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_111),
.A2(n_128),
.B1(n_131),
.B2(n_134),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_80),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_112),
.Y(n_168)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_102),
.B(n_23),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_72),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_136),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_126),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_83),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_86),
.A2(n_65),
.B1(n_68),
.B2(n_24),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_67),
.C(n_51),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_130),
.C(n_106),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_79),
.A2(n_41),
.B(n_33),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_86),
.A2(n_27),
.B1(n_57),
.B2(n_44),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_44),
.B1(n_42),
.B2(n_31),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_78),
.B(n_39),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_26),
.B1(n_42),
.B2(n_44),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_140),
.B1(n_93),
.B2(n_75),
.Y(n_176)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_95),
.A2(n_49),
.B1(n_41),
.B2(n_33),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_143),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_42),
.B1(n_36),
.B2(n_28),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_142),
.A2(n_107),
.B1(n_83),
.B2(n_104),
.Y(n_155)
);

AO22x1_ASAP7_75t_L g143 ( 
.A1(n_95),
.A2(n_41),
.B1(n_59),
.B2(n_32),
.Y(n_143)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_144),
.Y(n_150)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_176),
.B1(n_143),
.B2(n_141),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_152),
.A2(n_139),
.B(n_127),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_79),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_156),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_155),
.A2(n_167),
.B1(n_124),
.B2(n_123),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_113),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_175),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_77),
.C(n_91),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_161),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_108),
.A2(n_77),
.B(n_88),
.Y(n_161)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_121),
.B(n_39),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_173),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_84),
.B1(n_88),
.B2(n_40),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_93),
.C(n_75),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_140),
.B1(n_122),
.B2(n_120),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_178),
.A2(n_150),
.B1(n_169),
.B2(n_168),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_182),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_180),
.A2(n_176),
.B1(n_150),
.B2(n_169),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_177),
.B(n_125),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_196),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_111),
.B1(n_138),
.B2(n_133),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_194),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_130),
.B1(n_134),
.B2(n_132),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_177),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_198),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_160),
.Y(n_196)
);

BUFx12_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_197),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_135),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_200),
.A2(n_131),
.B(n_147),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_126),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_201),
.B(n_193),
.Y(n_214)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_168),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_187),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_137),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_161),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_185),
.C(n_198),
.Y(n_232)
);

OAI221xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_146),
.B1(n_170),
.B2(n_156),
.C(n_151),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_207),
.B(n_215),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_151),
.B(n_171),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_208),
.A2(n_199),
.B(n_189),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_193),
.B1(n_192),
.B2(n_196),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_211),
.B1(n_218),
.B2(n_186),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_221),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_191),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_219),
.B(n_144),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_SL g221 ( 
.A(n_191),
.B(n_146),
.C(n_136),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_182),
.B(n_175),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_226),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_225),
.Y(n_257)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_159),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_229),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_159),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_149),
.Y(n_230)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_197),
.B(n_112),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_231),
.A2(n_181),
.B(n_112),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_234),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_203),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_236),
.B(n_239),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_215),
.A2(n_200),
.B1(n_180),
.B2(n_194),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_242),
.B1(n_245),
.B2(n_209),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_222),
.B(n_206),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_204),
.C(n_194),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_213),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_255),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_194),
.B1(n_178),
.B2(n_184),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_246),
.A2(n_209),
.B(n_227),
.Y(n_278)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_199),
.C(n_188),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_214),
.B(n_190),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_223),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_258),
.A2(n_259),
.B(n_231),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_181),
.B(n_202),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

AOI322xp5_ASAP7_75t_SL g261 ( 
.A1(n_233),
.A2(n_207),
.A3(n_218),
.B1(n_208),
.B2(n_211),
.C1(n_217),
.C2(n_228),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_261),
.B(n_255),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_217),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_247),
.Y(n_267)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_284),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_212),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_277),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_278),
.B(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_283),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_233),
.A2(n_212),
.B(n_219),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_246),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_230),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_259),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_241),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_232),
.C(n_234),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_266),
.C(n_271),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_292),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_294),
.B(n_275),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_240),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_256),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_299),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_271),
.A2(n_245),
.B(n_238),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_243),
.B1(n_238),
.B2(n_249),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_295),
.A2(n_302),
.B1(n_265),
.B2(n_266),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_277),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_269),
.B(n_229),
.Y(n_299)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_267),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_305),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_278),
.A2(n_260),
.B1(n_165),
.B2(n_145),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_281),
.B(n_26),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_304),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_165),
.C(n_115),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_284),
.B(n_2),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_165),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_262),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_308),
.A2(n_298),
.B(n_287),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_324),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_313),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_317),
.C(n_321),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_262),
.C(n_276),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_273),
.Y(n_318)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_318),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_273),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_319),
.B(n_322),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_300),
.A2(n_270),
.B(n_264),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_306),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_276),
.C(n_270),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_264),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_296),
.A2(n_115),
.B1(n_149),
.B2(n_116),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_116),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_298),
.A2(n_290),
.B1(n_291),
.B2(n_288),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_295),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_335),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_338),
.B(n_334),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_314),
.C(n_321),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_333),
.C(n_104),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_304),
.C(n_302),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_334),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_294),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_307),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_339),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_320),
.A2(n_303),
.B(n_145),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_3),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_343),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_336),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_341),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_333),
.A2(n_316),
.B1(n_311),
.B2(n_145),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_316),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_345),
.B(n_349),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_332),
.B(n_3),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_347),
.B(n_348),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_329),
.B(n_3),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_329),
.B(n_4),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_351),
.B(n_4),
.Y(n_355)
);

NAND2x1_ASAP7_75t_SL g354 ( 
.A(n_344),
.B(n_331),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_355),
.B(n_356),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_330),
.Y(n_356)
);

AO21x1_ASAP7_75t_L g357 ( 
.A1(n_342),
.A2(n_325),
.B(n_6),
.Y(n_357)
);

AOI31xp67_ASAP7_75t_L g366 ( 
.A1(n_357),
.A2(n_9),
.A3(n_10),
.B(n_11),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_346),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_358),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_346),
.A2(n_343),
.B(n_345),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_360),
.B(n_5),
.C(n_7),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_364),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_353),
.A2(n_5),
.B(n_7),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_357),
.A2(n_40),
.B1(n_36),
.B2(n_30),
.Y(n_365)
);

OAI321xp33_ASAP7_75t_L g373 ( 
.A1(n_365),
.A2(n_366),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_373)
);

AOI31xp67_ASAP7_75t_L g367 ( 
.A1(n_354),
.A2(n_9),
.A3(n_10),
.B(n_11),
.Y(n_367)
);

NOR3xp33_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_9),
.C(n_10),
.Y(n_372)
);

NAND3xp33_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_352),
.C(n_361),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_371),
.B(n_372),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_373),
.A2(n_374),
.B1(n_30),
.B2(n_36),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_369),
.A2(n_361),
.B(n_359),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_370),
.B(n_368),
.C(n_359),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_377),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_375),
.A2(n_30),
.B1(n_40),
.B2(n_19),
.Y(n_378)
);

AOI321xp33_ASAP7_75t_L g380 ( 
.A1(n_378),
.A2(n_15),
.A3(n_18),
.B1(n_19),
.B2(n_32),
.C(n_379),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_18),
.Y(n_381)
);


endmodule