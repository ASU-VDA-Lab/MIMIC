module fake_jpeg_21202_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx2_ASAP7_75t_SL g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_31),
.B1(n_27),
.B2(n_17),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_31),
.B1(n_19),
.B2(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_23),
.B1(n_18),
.B2(n_25),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_17),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_31),
.B1(n_27),
.B2(n_25),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_17),
.B1(n_15),
.B2(n_28),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_46),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_55),
.B(n_23),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_60),
.B(n_69),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_76),
.B1(n_81),
.B2(n_82),
.Y(n_91)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_72),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_33),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_18),
.B1(n_23),
.B2(n_15),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_83),
.Y(n_100)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_80),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_21),
.Y(n_81)
);

AOI22x1_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_43),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_110),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_92),
.B(n_108),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_32),
.C(n_30),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_81),
.C(n_30),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_22),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_65),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_112),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_74),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_120),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_117),
.B(n_22),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_77),
.B1(n_85),
.B2(n_62),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_73),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_82),
.B1(n_81),
.B2(n_51),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_126),
.B1(n_136),
.B2(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_82),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_127),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_51),
.B1(n_78),
.B2(n_67),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_90),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_89),
.B(n_28),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_107),
.A3(n_24),
.B1(n_20),
.B2(n_29),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_58),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_135),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_58),
.B1(n_75),
.B2(n_28),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_85),
.B1(n_95),
.B2(n_86),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_30),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_19),
.B1(n_29),
.B2(n_24),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_19),
.B1(n_29),
.B2(n_24),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_30),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_30),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_30),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_68),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_155),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_147),
.A2(n_159),
.B1(n_163),
.B2(n_26),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_127),
.B(n_10),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_8),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_117),
.A2(n_95),
.B1(n_96),
.B2(n_94),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_106),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_152),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_199)
);

HAxp5_ASAP7_75t_SL g153 ( 
.A(n_141),
.B(n_106),
.CON(n_153),
.SN(n_153)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_153),
.B(n_8),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_86),
.B1(n_109),
.B2(n_94),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_129),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_120),
.A2(n_109),
.B1(n_96),
.B2(n_93),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_115),
.B1(n_136),
.B2(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_93),
.B1(n_88),
.B2(n_20),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_88),
.B(n_71),
.C(n_70),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_173),
.B(n_122),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_21),
.C(n_22),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_22),
.C(n_121),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_116),
.A2(n_123),
.B1(n_119),
.B2(n_140),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_165),
.B(n_170),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_119),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_169),
.Y(n_179)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_116),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_135),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_0),
.B(n_1),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_115),
.B1(n_134),
.B2(n_132),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_187),
.B1(n_201),
.B2(n_164),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_175),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_167),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_180),
.B(n_182),
.C(n_205),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_121),
.C(n_137),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_184),
.B(n_204),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_128),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_191),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_142),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_186),
.A2(n_147),
.B1(n_145),
.B2(n_144),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_0),
.B(n_2),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_190),
.B(n_192),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_9),
.B(n_14),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_26),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_9),
.B(n_14),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_12),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_154),
.B1(n_161),
.B2(n_156),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_142),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_2),
.B(n_3),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_10),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_26),
.C(n_10),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_207),
.B(n_211),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_216),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_183),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_212),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_181),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_214),
.B(n_220),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_218),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_185),
.B(n_191),
.Y(n_219)
);

A2O1A1O1Ixp25_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_200),
.B(n_223),
.C(n_216),
.D(n_220),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_168),
.Y(n_227)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_229),
.B(n_186),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_230),
.B(n_189),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_231),
.B(n_225),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_176),
.C(n_182),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_243),
.C(n_246),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_200),
.B(n_175),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_240),
.B(n_245),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_146),
.Y(n_241)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_242),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_188),
.C(n_143),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_208),
.A2(n_190),
.B(n_192),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_244),
.A2(n_210),
.B1(n_224),
.B2(n_215),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_195),
.C(n_205),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_146),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_248),
.Y(n_256)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_246),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_253),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_219),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_206),
.C(n_222),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_247),
.C(n_237),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_245),
.B(n_213),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_258),
.B(n_249),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_224),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_264),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_234),
.A2(n_218),
.B1(n_210),
.B2(n_206),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_263),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_177),
.B1(n_215),
.B2(n_202),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_262),
.A2(n_244),
.B1(n_236),
.B2(n_235),
.Y(n_274)
);

XOR2x1_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_152),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_230),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_274),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_256),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_277),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_242),
.C(n_235),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_275),
.C(n_272),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_232),
.C(n_236),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_263),
.A2(n_232),
.B1(n_145),
.B2(n_5),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_3),
.B(n_4),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_7),
.C(n_11),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_278),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_270),
.C(n_268),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_282),
.A2(n_265),
.B1(n_6),
.B2(n_3),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_264),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_288),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_254),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_287),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_262),
.B(n_11),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_288),
.B1(n_289),
.B2(n_283),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_297),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_266),
.B(n_13),
.Y(n_295)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_6),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_280),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_281),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_301),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_290),
.A2(n_298),
.B(n_294),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_302),
.A2(n_292),
.B(n_293),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_307),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_301),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_306),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_303),
.C(n_304),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_296),
.Y(n_313)
);


endmodule