module fake_jpeg_30514_n_277 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_42),
.Y(n_92)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_50),
.Y(n_66)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_19),
.A2(n_1),
.B(n_3),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_33),
.B(n_24),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_53),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_32),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_27),
.B1(n_28),
.B2(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_60),
.B1(n_69),
.B2(n_79),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_27),
.B1(n_28),
.B2(n_26),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_29),
.B1(n_31),
.B2(n_28),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_61),
.A2(n_63),
.B1(n_75),
.B2(n_88),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_18),
.B1(n_24),
.B2(n_36),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_62),
.A2(n_89),
.B1(n_8),
.B2(n_9),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_31),
.B1(n_37),
.B2(n_35),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_32),
.CON(n_67),
.SN(n_67)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_72),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_38),
.B1(n_31),
.B2(n_34),
.Y(n_69)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_25),
.B1(n_37),
.B2(n_30),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_31),
.B1(n_38),
.B2(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_90),
.Y(n_98)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_38),
.B1(n_18),
.B2(n_36),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_85),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_36),
.B1(n_34),
.B2(n_33),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_84),
.B1(n_94),
.B2(n_5),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_34),
.B1(n_33),
.B2(n_18),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_87),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_30),
.B1(n_21),
.B2(n_24),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_21),
.B1(n_22),
.B2(n_19),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_1),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_49),
.A2(n_22),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_22),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_104),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_22),
.B1(n_4),
.B2(n_5),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_22),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_3),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_107),
.B(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_3),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_11),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_120),
.B1(n_90),
.B2(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_7),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_10),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_70),
.B(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_7),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_116),
.B(n_128),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_63),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_92),
.B1(n_81),
.B2(n_61),
.Y(n_142)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_82),
.B(n_9),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_66),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_149),
.C(n_109),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_142),
.B1(n_147),
.B2(n_152),
.Y(n_160)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_143),
.B(n_13),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_88),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_146),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_99),
.B(n_91),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_97),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_75),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_68),
.B1(n_71),
.B2(n_74),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_74),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_120),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_68),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_68),
.B1(n_78),
.B2(n_64),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_101),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_96),
.B(n_80),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_108),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_176),
.C(n_154),
.Y(n_200)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_106),
.B(n_108),
.Y(n_161)
);

AO22x1_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_145),
.B1(n_134),
.B2(n_139),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_166),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_112),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_169),
.B(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_115),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_179),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_125),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_164),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_133),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_144),
.A2(n_107),
.B1(n_127),
.B2(n_103),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_142),
.B1(n_149),
.B2(n_145),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_123),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_178),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_118),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_126),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_102),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_181),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_124),
.B1(n_113),
.B2(n_78),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_156),
.B1(n_141),
.B2(n_132),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_153),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_185),
.A2(n_132),
.B(n_141),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_193),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_194),
.B1(n_204),
.B2(n_173),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_197),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_139),
.B1(n_143),
.B2(n_134),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_154),
.B1(n_130),
.B2(n_150),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_200),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_160),
.A2(n_150),
.B1(n_130),
.B2(n_113),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_218),
.B1(n_225),
.B2(n_192),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_176),
.C(n_159),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_216),
.C(n_219),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_165),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_217),
.B1(n_220),
.B2(n_222),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_161),
.B(n_163),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_212),
.B(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_172),
.C(n_179),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_163),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_171),
.C(n_175),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_162),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_161),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_158),
.C(n_168),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_189),
.C(n_201),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_184),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_188),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_177),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_230),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_187),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_234),
.C(n_235),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_204),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_209),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_216),
.B(n_182),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_236),
.A2(n_219),
.B1(n_218),
.B2(n_220),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_191),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_237),
.B(n_235),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_239),
.B(n_248),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_187),
.B1(n_193),
.B2(n_202),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_244),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_212),
.B(n_234),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_249),
.B(n_233),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_240),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_224),
.C(n_213),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_213),
.C(n_203),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_232),
.B1(n_202),
.B2(n_237),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_251),
.B(n_248),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_255),
.C(n_247),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_249),
.A2(n_203),
.B1(n_198),
.B2(n_174),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_198),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_246),
.C(n_228),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_258),
.B(n_228),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_262),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_263),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_246),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_257),
.B1(n_256),
.B2(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_266),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_181),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_263),
.B1(n_183),
.B2(n_101),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_269),
.B(n_265),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_273),
.B1(n_269),
.B2(n_271),
.Y(n_274)
);

AOI332xp33_ASAP7_75t_L g273 ( 
.A1(n_270),
.A2(n_267),
.A3(n_140),
.B1(n_13),
.B2(n_14),
.B3(n_78),
.C1(n_87),
.C2(n_64),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_95),
.C(n_14),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_14),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_87),
.Y(n_277)
);


endmodule