module fake_jpeg_11456_n_208 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_8),
.B(n_12),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_50),
.Y(n_80)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_58),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_13),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_13),
.B(n_0),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_60),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_64),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_21),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_63),
.Y(n_96)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_22),
.B(n_1),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_66),
.Y(n_104)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_70),
.Y(n_87)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_75)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_25),
.B(n_2),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_23),
.B1(n_21),
.B2(n_28),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_40),
.A2(n_34),
.B1(n_23),
.B2(n_5),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_97),
.B1(n_77),
.B2(n_85),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_2),
.B1(n_4),
.B2(n_9),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_53),
.A2(n_10),
.B1(n_54),
.B2(n_47),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_55),
.B1(n_57),
.B2(n_70),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_62),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_50),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_108),
.B(n_118),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_121),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_130),
.C(n_131),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_88),
.C(n_106),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_119),
.C(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_126),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_97),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_93),
.B1(n_75),
.B2(n_85),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_124),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_89),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_75),
.B(n_94),
.C(n_105),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_89),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_99),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_132),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_100),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_73),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_101),
.B1(n_74),
.B2(n_73),
.Y(n_132)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_73),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_146),
.Y(n_157)
);

AOI32xp33_ASAP7_75t_L g146 ( 
.A1(n_112),
.A2(n_109),
.A3(n_107),
.B1(n_110),
.B2(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_127),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_122),
.CI(n_125),
.CON(n_150),
.SN(n_150)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_153),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_159),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_138),
.A2(n_124),
.B1(n_122),
.B2(n_132),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_155),
.A2(n_164),
.B(n_135),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_140),
.A2(n_122),
.B1(n_120),
.B2(n_129),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_158),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_123),
.B1(n_119),
.B2(n_114),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_148),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_133),
.B(n_139),
.Y(n_166)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_167),
.B(n_134),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_144),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_169),
.B(n_171),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_135),
.B(n_134),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_170),
.A2(n_155),
.B(n_157),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_151),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_156),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_177),
.A2(n_179),
.B(n_180),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_178),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_146),
.C(n_145),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_175),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_185),
.C(n_167),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_170),
.A2(n_153),
.B1(n_165),
.B2(n_150),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_184),
.A2(n_172),
.B1(n_137),
.B2(n_150),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_136),
.C(n_149),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_177),
.B(n_184),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_172),
.C(n_173),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_189),
.B(n_141),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_179),
.B1(n_137),
.B2(n_183),
.Y(n_194)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_190),
.A2(n_168),
.B(n_135),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_R g200 ( 
.A(n_195),
.B(n_187),
.C(n_141),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_196),
.A2(n_188),
.B1(n_186),
.B2(n_189),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_163),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_196),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_201),
.A2(n_203),
.B(n_200),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_198),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_199),
.A2(n_160),
.B(n_163),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_206),
.A2(n_197),
.B1(n_130),
.B2(n_111),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_119),
.Y(n_208)
);


endmodule