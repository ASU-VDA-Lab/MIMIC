module fake_jpeg_55_n_197 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_197);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_3),
.B(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_13),
.B(n_9),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_20),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_R g70 ( 
.A(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_0),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_76),
.Y(n_92)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_2),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_77),
.B(n_70),
.Y(n_82)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_61),
.B1(n_63),
.B2(n_68),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_81),
.B1(n_78),
.B2(n_65),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_54),
.B(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_74),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_57),
.B1(n_58),
.B2(n_50),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_89),
.B1(n_91),
.B2(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_57),
.B1(n_58),
.B2(n_50),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_63),
.B1(n_61),
.B2(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_94),
.B(n_97),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_95),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_92),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_107),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_106),
.Y(n_123)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_56),
.A3(n_55),
.B1(n_49),
.B2(n_78),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_6),
.Y(n_125)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_104),
.Y(n_127)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_55),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_65),
.B1(n_87),
.B2(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_108),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_48),
.B(n_41),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_52),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_116),
.C(n_126),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_122),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_90),
.Y(n_116)
);

AO22x2_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_69),
.B1(n_60),
.B2(n_51),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_3),
.B(n_5),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_119),
.A2(n_7),
.B(n_10),
.Y(n_135)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_105),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_11),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_24),
.C(n_47),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_129),
.A2(n_100),
.B1(n_8),
.B2(n_10),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_100),
.B1(n_26),
.B2(n_27),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_135),
.B(n_149),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_25),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_144),
.C(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_28),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_142),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_148),
.B1(n_150),
.B2(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

NOR2xp67_ASAP7_75t_R g162 ( 
.A(n_141),
.B(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_12),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_32),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_127),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_147),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_31),
.B1(n_44),
.B2(n_43),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_126),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_121),
.B(n_118),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_118),
.B(n_111),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_153),
.B(n_155),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_118),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_166),
.C(n_169),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_111),
.B1(n_15),
.B2(n_16),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_18),
.B(n_19),
.Y(n_164)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_34),
.C(n_35),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_167)
);

OAI321xp33_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_150),
.A3(n_134),
.B1(n_146),
.B2(n_144),
.C(n_21),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_37),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_132),
.C(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_177),
.Y(n_180)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_170),
.B(n_40),
.CI(n_159),
.CON(n_179),
.SN(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_169),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_174),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_181),
.B(n_173),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_161),
.B(n_158),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_184),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_178),
.A2(n_161),
.B(n_162),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_183),
.A2(n_185),
.B(n_186),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_153),
.B(n_176),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_166),
.B(n_165),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_190),
.B(n_185),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_180),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_172),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_193),
.Y(n_194)
);

OAI31xp33_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_179),
.A3(n_164),
.B(n_168),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_156),
.C(n_179),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_194),
.Y(n_197)
);


endmodule