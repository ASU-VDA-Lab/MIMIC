module fake_jpeg_8897_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_8),
.B(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_15),
.B(n_11),
.C(n_16),
.Y(n_24)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_10),
.B1(n_21),
.B2(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_15),
.Y(n_31)
);

NOR2x1_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_14),
.Y(n_35)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_23),
.B1(n_27),
.B2(n_18),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_35),
.B(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_25),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_37),
.B1(n_42),
.B2(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_33),
.B1(n_30),
.B2(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_47),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_35),
.C(n_29),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_49),
.C(n_50),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_34),
.C(n_29),
.Y(n_50)
);

AOI322xp5_ASAP7_75t_SL g51 ( 
.A1(n_50),
.A2(n_37),
.A3(n_36),
.B1(n_11),
.B2(n_16),
.C1(n_9),
.C2(n_5),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_5),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_40),
.C(n_16),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_56),
.C(n_9),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_16),
.C(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_57),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_62),
.C(n_51),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_49),
.B(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx24_ASAP7_75t_SL g66 ( 
.A(n_63),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_68),
.B(n_70),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_66),
.A3(n_69),
.B1(n_19),
.B2(n_17),
.C1(n_9),
.C2(n_4),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_74),
.C(n_2),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_17),
.A3(n_19),
.B1(n_3),
.B2(n_4),
.C1(n_0),
.C2(n_2),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_3),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_3),
.Y(n_77)
);


endmodule