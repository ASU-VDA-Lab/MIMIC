module real_jpeg_29357_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_0),
.A2(n_43),
.B1(n_44),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_0),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_1),
.A2(n_41),
.B(n_45),
.Y(n_40)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_3),
.B(n_24),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_3),
.A2(n_24),
.B(n_71),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_3),
.A2(n_11),
.B(n_43),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_3),
.B(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_160),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_6),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_64),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_64),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_49),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_67),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_10),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_152)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_12),
.A2(n_26),
.B1(n_91),
.B2(n_92),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_12),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_12),
.A2(n_26),
.B1(n_43),
.B2(n_44),
.Y(n_160)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_113),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_111),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_79),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_19),
.B(n_79),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_57),
.C(n_69),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_20),
.A2(n_21),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_38),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_22),
.B(n_39),
.C(n_51),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_31),
.B2(n_36),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_23),
.A2(n_27),
.B1(n_31),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_24),
.A2(n_25),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_55),
.Y(n_89)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI32xp33_ASAP7_75t_L g70 ( 
.A1(n_25),
.A2(n_32),
.A3(n_35),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_25),
.A2(n_89),
.B1(n_90),
.B2(n_93),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_27),
.A2(n_31),
.B1(n_36),
.B2(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g72 ( 
.A(n_29),
.B(n_33),
.Y(n_72)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_31),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_33),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_33),
.A2(n_52),
.B(n_61),
.C(n_136),
.Y(n_135)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_50),
.B2(n_51),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_47),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_44),
.B1(n_60),
.B2(n_61),
.Y(n_62)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_44),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_46),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_46),
.A2(n_87),
.B1(n_152),
.B2(n_160),
.Y(n_159)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_47),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_47),
.B(n_52),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_77),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

HAxp5_ASAP7_75t_SL g90 ( 
.A(n_52),
.B(n_91),
.CON(n_90),
.SN(n_90)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_52),
.B(n_62),
.Y(n_158)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_54),
.A2(n_90),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_54),
.A2(n_55),
.B(n_91),
.C(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_91),
.Y(n_93)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_57),
.B(n_69),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_63),
.B(n_65),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_58),
.A2(n_62),
.B1(n_63),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_62),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_58),
.A2(n_62),
.B1(n_123),
.B2(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_73),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_74),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_75),
.A2(n_147),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_96),
.B1(n_97),
.B2(n_110),
.Y(n_79)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_94),
.B2(n_95),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_127),
.B(n_174),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_124),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_115),
.B(n_124),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.C(n_121),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_116),
.A2(n_117),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_168),
.B(n_173),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_148),
.B(n_167),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_135),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_143),
.C(n_144),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_156),
.B(n_166),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_154),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_161),
.B(n_165),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_158),
.B(n_159),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_169),
.B(n_170),
.Y(n_173)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);


endmodule