module real_aes_8412_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g256 ( .A1(n_0), .A2(n_257), .B(n_258), .C(n_261), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_1), .B(n_198), .Y(n_262) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
NAND3xp33_ASAP7_75t_SL g730 ( .A(n_2), .B(n_704), .C(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_3), .B(n_168), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_4), .A2(n_138), .B(n_141), .C(n_446), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_5), .A2(n_158), .B(n_486), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_6), .A2(n_158), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_7), .B(n_198), .Y(n_492) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_8), .A2(n_125), .B(n_178), .Y(n_177) );
AND2x6_ASAP7_75t_L g138 ( .A(n_9), .B(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_10), .A2(n_138), .B(n_141), .C(n_144), .Y(n_140) );
INVx1_ASAP7_75t_L g462 ( .A(n_11), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_12), .B(n_39), .Y(n_113) );
INVx1_ASAP7_75t_L g728 ( .A(n_12), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_13), .B(n_148), .Y(n_448) );
INVx1_ASAP7_75t_L g130 ( .A(n_14), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_15), .B(n_168), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_16), .A2(n_146), .B(n_470), .C(n_472), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_17), .B(n_198), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_18), .B(n_222), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_19), .A2(n_141), .B(n_185), .C(n_218), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_20), .A2(n_150), .B(n_260), .C(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_21), .B(n_148), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_22), .B(n_148), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_23), .Y(n_520) );
INVx1_ASAP7_75t_L g512 ( .A(n_24), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_25), .A2(n_141), .B(n_181), .C(n_185), .Y(n_180) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_26), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_27), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_28), .Y(n_444) );
INVx1_ASAP7_75t_L g503 ( .A(n_29), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_30), .A2(n_158), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g136 ( .A(n_31), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_32), .A2(n_160), .B(n_171), .C(n_206), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_33), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_34), .A2(n_260), .B(n_489), .C(n_491), .Y(n_488) );
INVxp67_ASAP7_75t_L g504 ( .A(n_35), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_36), .B(n_183), .Y(n_182) );
CKINVDCx14_ASAP7_75t_R g487 ( .A(n_37), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_38), .A2(n_141), .B(n_185), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_39), .B(n_728), .Y(n_727) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_40), .A2(n_261), .B(n_460), .C(n_461), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_41), .B(n_216), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_42), .Y(n_153) );
AOI222xp33_ASAP7_75t_L g114 ( .A1(n_43), .A2(n_69), .B1(n_115), .B2(n_705), .C1(n_710), .C2(n_711), .Y(n_114) );
INVx1_ASAP7_75t_L g710 ( .A(n_43), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_44), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_45), .B(n_158), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_46), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_47), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g159 ( .A1(n_48), .A2(n_160), .B(n_162), .C(n_171), .Y(n_159) );
INVx1_ASAP7_75t_L g259 ( .A(n_49), .Y(n_259) );
INVx1_ASAP7_75t_L g163 ( .A(n_50), .Y(n_163) );
INVx1_ASAP7_75t_L g477 ( .A(n_51), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_52), .B(n_158), .Y(n_157) );
AOI22xp33_ASAP7_75t_SL g99 ( .A1(n_53), .A2(n_100), .B1(n_723), .B2(n_734), .Y(n_99) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_54), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_54), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_55), .Y(n_225) );
CKINVDCx14_ASAP7_75t_R g458 ( .A(n_56), .Y(n_458) );
INVx1_ASAP7_75t_L g139 ( .A(n_57), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_58), .B(n_158), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_59), .B(n_198), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_60), .A2(n_192), .B(n_194), .C(n_196), .Y(n_191) );
INVx1_ASAP7_75t_L g129 ( .A(n_61), .Y(n_129) );
INVx1_ASAP7_75t_SL g490 ( .A(n_62), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_63), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_64), .B(n_168), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_65), .B(n_198), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_66), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g523 ( .A(n_67), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_68), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_70), .B(n_165), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_71), .A2(n_141), .B(n_171), .C(n_232), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_72), .Y(n_190) );
INVx1_ASAP7_75t_L g733 ( .A(n_73), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_74), .A2(n_158), .B(n_457), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_75), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_76), .A2(n_158), .B(n_467), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_77), .A2(n_216), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g468 ( .A(n_78), .Y(n_468) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_79), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_80), .B(n_164), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_81), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_82), .A2(n_158), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g471 ( .A(n_83), .Y(n_471) );
INVx2_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
INVx1_ASAP7_75t_L g447 ( .A(n_85), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_86), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_87), .B(n_148), .Y(n_147) );
OR2x2_ASAP7_75t_L g109 ( .A(n_88), .B(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g434 ( .A(n_88), .B(n_111), .Y(n_434) );
INVx2_ASAP7_75t_L g704 ( .A(n_88), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_89), .A2(n_141), .B(n_171), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_90), .B(n_158), .Y(n_204) );
INVx1_ASAP7_75t_L g207 ( .A(n_91), .Y(n_207) );
INVxp67_ASAP7_75t_L g195 ( .A(n_92), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_93), .B(n_125), .Y(n_463) );
INVx1_ASAP7_75t_L g132 ( .A(n_94), .Y(n_132) );
INVx1_ASAP7_75t_L g233 ( .A(n_95), .Y(n_233) );
INVx2_ASAP7_75t_L g480 ( .A(n_96), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_97), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g174 ( .A(n_98), .B(n_173), .Y(n_174) );
AOI22xp5_ASAP7_75t_SL g100 ( .A1(n_101), .A2(n_114), .B1(n_714), .B2(n_715), .Y(n_100) );
NOR2xp33_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g714 ( .A(n_103), .Y(n_714) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_105), .A2(n_716), .B(n_720), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_109), .Y(n_722) );
NOR2x2_ASAP7_75t_L g713 ( .A(n_110), .B(n_704), .Y(n_713) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g703 ( .A(n_111), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
OAI22xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_432), .B1(n_435), .B2(n_701), .Y(n_115) );
INVx2_ASAP7_75t_L g707 ( .A(n_116), .Y(n_707) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_116), .Y(n_718) );
OR3x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_330), .C(n_395), .Y(n_116) );
NAND4xp25_ASAP7_75t_SL g117 ( .A(n_118), .B(n_271), .C(n_297), .D(n_320), .Y(n_117) );
AOI221xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_199), .B1(n_240), .B2(n_247), .C(n_263), .Y(n_118) );
CKINVDCx14_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_120), .A2(n_264), .B1(n_288), .B2(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_175), .Y(n_120) );
INVx1_ASAP7_75t_SL g324 ( .A(n_121), .Y(n_324) );
OR2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_155), .Y(n_121) );
OR2x2_ASAP7_75t_L g245 ( .A(n_122), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g266 ( .A(n_122), .B(n_176), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_122), .B(n_186), .Y(n_279) );
AND2x2_ASAP7_75t_L g296 ( .A(n_122), .B(n_155), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_122), .B(n_243), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_122), .B(n_295), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_122), .B(n_175), .Y(n_417) );
AOI211xp5_ASAP7_75t_SL g428 ( .A1(n_122), .A2(n_334), .B(n_429), .C(n_430), .Y(n_428) );
INVx5_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_123), .B(n_176), .Y(n_300) );
AND2x2_ASAP7_75t_L g303 ( .A(n_123), .B(n_177), .Y(n_303) );
OR2x2_ASAP7_75t_L g348 ( .A(n_123), .B(n_176), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_123), .B(n_186), .Y(n_357) );
AO21x2_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_131), .B(n_152), .Y(n_123) );
INVx3_ASAP7_75t_L g198 ( .A(n_124), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_124), .B(n_210), .Y(n_209) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_124), .A2(n_230), .B(n_238), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_124), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_124), .B(n_451), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_124), .B(n_515), .Y(n_514) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_124), .A2(n_519), .B(n_525), .Y(n_518) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_125), .A2(n_179), .B(n_180), .Y(n_178) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_127), .B(n_128), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
OAI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_140), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g443 ( .A1(n_133), .A2(n_444), .B(n_445), .Y(n_443) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_133), .A2(n_173), .B(n_509), .C(n_510), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_133), .A2(n_520), .B(n_521), .Y(n_519) );
NAND2x1p5_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
AND2x4_ASAP7_75t_L g158 ( .A(n_134), .B(n_138), .Y(n_158) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g196 ( .A(n_135), .Y(n_196) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx1_ASAP7_75t_L g151 ( .A(n_136), .Y(n_151) );
INVx1_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
INVx3_ASAP7_75t_L g146 ( .A(n_137), .Y(n_146) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_137), .Y(n_148) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_137), .Y(n_166) );
INVx1_ASAP7_75t_L g183 ( .A(n_137), .Y(n_183) );
INVx4_ASAP7_75t_SL g172 ( .A(n_138), .Y(n_172) );
BUFx3_ASAP7_75t_L g185 ( .A(n_138), .Y(n_185) );
INVx5_ASAP7_75t_L g161 ( .A(n_141), .Y(n_161) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx3_ASAP7_75t_L g170 ( .A(n_142), .Y(n_170) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_142), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_147), .B(n_149), .Y(n_144) );
INVx5_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_146), .B(n_462), .Y(n_461) );
INVx4_ASAP7_75t_L g260 ( .A(n_148), .Y(n_260) );
INVx2_ASAP7_75t_L g460 ( .A(n_148), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_149), .A2(n_182), .B(n_184), .Y(n_181) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
INVx2_ASAP7_75t_L g497 ( .A(n_154), .Y(n_497) );
INVx5_ASAP7_75t_SL g246 ( .A(n_155), .Y(n_246) );
AND2x2_ASAP7_75t_L g265 ( .A(n_155), .B(n_266), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_155), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g351 ( .A(n_155), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g383 ( .A(n_155), .B(n_186), .Y(n_383) );
OR2x2_ASAP7_75t_L g389 ( .A(n_155), .B(n_279), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_155), .B(n_339), .Y(n_398) );
OR2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_174), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_173), .Y(n_156) );
BUFx2_ASAP7_75t_L g216 ( .A(n_158), .Y(n_216) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_161), .A2(n_172), .B(n_190), .C(n_191), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_SL g254 ( .A1(n_161), .A2(n_172), .B(n_255), .C(n_256), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g457 ( .A1(n_161), .A2(n_172), .B(n_458), .C(n_459), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_SL g467 ( .A1(n_161), .A2(n_172), .B(n_468), .C(n_469), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_SL g476 ( .A1(n_161), .A2(n_172), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_161), .A2(n_172), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_SL g499 ( .A1(n_161), .A2(n_172), .B(n_500), .C(n_501), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_167), .C(n_169), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_164), .A2(n_169), .B(n_207), .C(n_208), .Y(n_206) );
O2A1O1Ixp5_ASAP7_75t_L g446 ( .A1(n_164), .A2(n_447), .B(n_448), .C(n_449), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_164), .A2(n_449), .B(n_523), .C(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx4_ASAP7_75t_L g193 ( .A(n_166), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_168), .B(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g257 ( .A(n_168), .Y(n_257) );
OAI22xp33_ASAP7_75t_L g502 ( .A1(n_168), .A2(n_193), .B1(n_503), .B2(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_168), .A2(n_221), .B(n_512), .C(n_513), .Y(n_511) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g261 ( .A(n_170), .Y(n_261) );
INVx1_ASAP7_75t_L g472 ( .A(n_170), .Y(n_472) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_173), .A2(n_204), .B(n_205), .Y(n_203) );
INVx2_ASAP7_75t_L g223 ( .A(n_173), .Y(n_223) );
INVx1_ASAP7_75t_L g226 ( .A(n_173), .Y(n_226) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_173), .A2(n_456), .B(n_463), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_186), .Y(n_175) );
AND2x2_ASAP7_75t_L g280 ( .A(n_176), .B(n_246), .Y(n_280) );
INVx1_ASAP7_75t_SL g293 ( .A(n_176), .Y(n_293) );
OR2x2_ASAP7_75t_L g328 ( .A(n_176), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g334 ( .A(n_176), .B(n_186), .Y(n_334) );
AND2x2_ASAP7_75t_L g392 ( .A(n_176), .B(n_243), .Y(n_392) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_177), .B(n_246), .Y(n_319) );
INVx3_ASAP7_75t_L g243 ( .A(n_186), .Y(n_243) );
OR2x2_ASAP7_75t_L g285 ( .A(n_186), .B(n_246), .Y(n_285) );
AND2x2_ASAP7_75t_L g295 ( .A(n_186), .B(n_293), .Y(n_295) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_186), .Y(n_343) );
AND2x2_ASAP7_75t_L g352 ( .A(n_186), .B(n_266), .Y(n_352) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_197), .Y(n_186) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_187), .A2(n_466), .B(n_473), .Y(n_465) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_187), .A2(n_475), .B(n_481), .Y(n_474) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_187), .A2(n_485), .B(n_492), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_192), .A2(n_233), .B(n_234), .C(n_235), .Y(n_232) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_193), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_193), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g221 ( .A(n_196), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_196), .B(n_502), .Y(n_501) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_198), .A2(n_253), .B(n_262), .Y(n_252) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_199), .A2(n_369), .B1(n_371), .B2(n_373), .C(n_376), .Y(n_368) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
AND2x2_ASAP7_75t_L g342 ( .A(n_201), .B(n_323), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_201), .B(n_401), .Y(n_405) );
OR2x2_ASAP7_75t_L g426 ( .A(n_201), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_201), .B(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx5_ASAP7_75t_L g273 ( .A(n_202), .Y(n_273) );
AND2x2_ASAP7_75t_L g350 ( .A(n_202), .B(n_213), .Y(n_350) );
AND2x2_ASAP7_75t_L g411 ( .A(n_202), .B(n_290), .Y(n_411) );
AND2x2_ASAP7_75t_L g424 ( .A(n_202), .B(n_243), .Y(n_424) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_209), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_227), .Y(n_211) );
AND2x4_ASAP7_75t_L g250 ( .A(n_212), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g269 ( .A(n_212), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g276 ( .A(n_212), .Y(n_276) );
AND2x2_ASAP7_75t_L g345 ( .A(n_212), .B(n_323), .Y(n_345) );
AND2x2_ASAP7_75t_L g355 ( .A(n_212), .B(n_273), .Y(n_355) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_212), .Y(n_363) );
AND2x2_ASAP7_75t_L g375 ( .A(n_212), .B(n_252), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_212), .B(n_307), .Y(n_379) );
AND2x2_ASAP7_75t_L g416 ( .A(n_212), .B(n_411), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_212), .B(n_290), .Y(n_427) );
OR2x2_ASAP7_75t_L g429 ( .A(n_212), .B(n_365), .Y(n_429) );
INVx5_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g315 ( .A(n_213), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g325 ( .A(n_213), .B(n_270), .Y(n_325) );
AND2x2_ASAP7_75t_L g337 ( .A(n_213), .B(n_252), .Y(n_337) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_213), .Y(n_367) );
AND2x4_ASAP7_75t_L g401 ( .A(n_213), .B(n_251), .Y(n_401) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
AOI21xp5_ASAP7_75t_SL g214 ( .A1(n_215), .A2(n_217), .B(n_222), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_218) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_223), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
AO21x2_ASAP7_75t_L g442 ( .A1(n_226), .A2(n_443), .B(n_450), .Y(n_442) );
BUFx2_ASAP7_75t_L g249 ( .A(n_227), .Y(n_249) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g290 ( .A(n_228), .Y(n_290) );
AND2x2_ASAP7_75t_L g323 ( .A(n_228), .B(n_252), .Y(n_323) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g270 ( .A(n_229), .B(n_252), .Y(n_270) );
BUFx2_ASAP7_75t_L g316 ( .A(n_229), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_237), .Y(n_230) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g491 ( .A(n_236), .Y(n_491) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_242), .B(n_324), .Y(n_403) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_243), .B(n_266), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_243), .B(n_246), .Y(n_305) );
AND2x2_ASAP7_75t_L g360 ( .A(n_243), .B(n_296), .Y(n_360) );
AOI221xp5_ASAP7_75t_SL g297 ( .A1(n_244), .A2(n_298), .B1(n_306), .B2(n_308), .C(n_312), .Y(n_297) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g292 ( .A(n_245), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g333 ( .A(n_245), .B(n_334), .Y(n_333) );
OAI321xp33_ASAP7_75t_L g340 ( .A1(n_245), .A2(n_299), .A3(n_341), .B1(n_343), .B2(n_344), .C(n_346), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_246), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_249), .B(n_401), .Y(n_419) );
AND2x2_ASAP7_75t_L g306 ( .A(n_250), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_250), .B(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_251), .Y(n_282) );
AND2x2_ASAP7_75t_L g289 ( .A(n_251), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_251), .B(n_364), .Y(n_394) );
INVx1_ASAP7_75t_L g431 ( .A(n_251), .Y(n_431) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_260), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g449 ( .A(n_261), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_267), .B(n_268), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g423 ( .A1(n_265), .A2(n_375), .B(n_424), .C(n_425), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_266), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_266), .B(n_304), .Y(n_370) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g313 ( .A(n_270), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_270), .B(n_273), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_270), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_270), .B(n_355), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_274), .B1(n_286), .B2(n_291), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g287 ( .A(n_273), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g310 ( .A(n_273), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g322 ( .A(n_273), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_273), .B(n_316), .Y(n_358) );
OR2x2_ASAP7_75t_L g365 ( .A(n_273), .B(n_290), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_273), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g415 ( .A(n_273), .B(n_401), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_277), .B1(n_281), .B2(n_283), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g321 ( .A(n_276), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
OAI22xp33_ASAP7_75t_L g361 ( .A1(n_279), .A2(n_294), .B1(n_362), .B2(n_366), .Y(n_361) );
INVx1_ASAP7_75t_L g409 ( .A(n_280), .Y(n_409) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_284), .A2(n_321), .B1(n_324), .B2(n_325), .C(n_326), .Y(n_320) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g299 ( .A(n_285), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_289), .B(n_355), .Y(n_387) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_290), .Y(n_307) );
INVx1_ASAP7_75t_L g311 ( .A(n_290), .Y(n_311) );
NAND2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g329 ( .A(n_296), .Y(n_329) );
AND2x2_ASAP7_75t_L g338 ( .A(n_296), .B(n_339), .Y(n_338) );
NAND2xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x2_ASAP7_75t_L g382 ( .A(n_303), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g331 ( .A1(n_306), .A2(n_332), .B1(n_335), .B2(n_338), .C(n_340), .Y(n_331) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_310), .B(n_367), .Y(n_366) );
AOI21xp33_ASAP7_75t_SL g312 ( .A1(n_313), .A2(n_314), .B(n_317), .Y(n_312) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
CKINVDCx16_ASAP7_75t_R g414 ( .A(n_317), .Y(n_414) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
OR2x2_ASAP7_75t_L g356 ( .A(n_319), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g377 ( .A(n_322), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_322), .B(n_382), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_325), .B(n_347), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NAND4xp25_ASAP7_75t_L g330 ( .A(n_331), .B(n_349), .C(n_368), .D(n_381), .Y(n_330) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g339 ( .A(n_334), .Y(n_339) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g372 ( .A(n_343), .B(n_348), .Y(n_372) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI211xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B(n_353), .C(n_361), .Y(n_349) );
AOI211xp5_ASAP7_75t_L g420 ( .A1(n_351), .A2(n_393), .B(n_421), .C(n_428), .Y(n_420) );
INVx1_ASAP7_75t_SL g380 ( .A(n_352), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_356), .B1(n_358), .B2(n_359), .Y(n_353) );
INVx1_ASAP7_75t_L g384 ( .A(n_358), .Y(n_384) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_364), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_364), .B(n_375), .Y(n_408) );
INVx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g385 ( .A(n_375), .Y(n_385) );
AOI21xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B(n_380), .Y(n_376) );
INVxp33_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI322xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .A3(n_385), .B1(n_386), .B2(n_388), .C1(n_390), .C2(n_393), .Y(n_381) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND3xp33_ASAP7_75t_SL g395 ( .A(n_396), .B(n_413), .C(n_420), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B1(n_402), .B2(n_404), .C(n_406), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g412 ( .A(n_401), .Y(n_412) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_409), .B2(n_410), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B1(n_416), .B2(n_417), .C(n_418), .Y(n_413) );
NAND2xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g706 ( .A(n_433), .Y(n_706) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g708 ( .A(n_435), .Y(n_708) );
OR2x2_ASAP7_75t_SL g435 ( .A(n_436), .B(n_656), .Y(n_435) );
NAND5xp2_ASAP7_75t_L g436 ( .A(n_437), .B(n_568), .C(n_606), .D(n_627), .E(n_644), .Y(n_436) );
NOR3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_540), .C(n_561), .Y(n_437) );
OAI221xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_482), .B1(n_506), .B2(n_527), .C(n_531), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_452), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_441), .B(n_529), .Y(n_548) );
OR2x2_ASAP7_75t_L g575 ( .A(n_441), .B(n_465), .Y(n_575) );
AND2x2_ASAP7_75t_L g589 ( .A(n_441), .B(n_465), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_441), .B(n_455), .Y(n_603) );
AND2x2_ASAP7_75t_L g641 ( .A(n_441), .B(n_605), .Y(n_641) );
AND2x2_ASAP7_75t_L g670 ( .A(n_441), .B(n_580), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_441), .B(n_552), .Y(n_687) );
INVx4_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g567 ( .A(n_442), .B(n_464), .Y(n_567) );
BUFx3_ASAP7_75t_L g592 ( .A(n_442), .Y(n_592) );
AND2x2_ASAP7_75t_L g621 ( .A(n_442), .B(n_465), .Y(n_621) );
AND3x2_ASAP7_75t_L g634 ( .A(n_442), .B(n_635), .C(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g557 ( .A(n_452), .Y(n_557) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_464), .Y(n_452) );
AOI32xp33_ASAP7_75t_L g612 ( .A1(n_453), .A2(n_564), .A3(n_613), .B1(n_616), .B2(n_617), .Y(n_612) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g539 ( .A(n_454), .B(n_464), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_454), .B(n_567), .Y(n_610) );
AND2x2_ASAP7_75t_L g617 ( .A(n_454), .B(n_589), .Y(n_617) );
OR2x2_ASAP7_75t_L g623 ( .A(n_454), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_454), .B(n_578), .Y(n_648) );
OR2x2_ASAP7_75t_L g666 ( .A(n_454), .B(n_494), .Y(n_666) );
BUFx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g530 ( .A(n_455), .B(n_474), .Y(n_530) );
INVx2_ASAP7_75t_L g552 ( .A(n_455), .Y(n_552) );
OR2x2_ASAP7_75t_L g574 ( .A(n_455), .B(n_474), .Y(n_574) );
AND2x2_ASAP7_75t_L g579 ( .A(n_455), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_455), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g635 ( .A(n_455), .B(n_529), .Y(n_635) );
INVx1_ASAP7_75t_SL g686 ( .A(n_464), .Y(n_686) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_474), .Y(n_464) );
INVx1_ASAP7_75t_SL g529 ( .A(n_465), .Y(n_529) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_465), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_465), .B(n_615), .Y(n_614) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_465), .B(n_552), .C(n_670), .Y(n_681) );
INVx2_ASAP7_75t_L g580 ( .A(n_474), .Y(n_580) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_474), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_493), .Y(n_482) );
INVx1_ASAP7_75t_L g616 ( .A(n_483), .Y(n_616) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g534 ( .A(n_484), .B(n_517), .Y(n_534) );
INVx2_ASAP7_75t_L g551 ( .A(n_484), .Y(n_551) );
AND2x2_ASAP7_75t_L g556 ( .A(n_484), .B(n_518), .Y(n_556) );
AND2x2_ASAP7_75t_L g571 ( .A(n_484), .B(n_507), .Y(n_571) );
AND2x2_ASAP7_75t_L g583 ( .A(n_484), .B(n_555), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_493), .B(n_599), .Y(n_598) );
NAND2x1p5_ASAP7_75t_L g655 ( .A(n_493), .B(n_556), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_493), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_493), .B(n_550), .Y(n_678) );
BUFx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OR2x2_ASAP7_75t_L g516 ( .A(n_494), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_494), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g560 ( .A(n_494), .B(n_507), .Y(n_560) );
AND2x2_ASAP7_75t_L g586 ( .A(n_494), .B(n_517), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_494), .B(n_626), .Y(n_625) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .B(n_505), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_496), .A2(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g545 ( .A(n_498), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_505), .Y(n_546) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_507), .B(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g550 ( .A(n_507), .B(n_551), .Y(n_550) );
INVx3_ASAP7_75t_SL g555 ( .A(n_507), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_507), .B(n_542), .Y(n_608) );
OR2x2_ASAP7_75t_L g618 ( .A(n_507), .B(n_544), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_507), .B(n_586), .Y(n_646) );
OR2x2_ASAP7_75t_L g676 ( .A(n_507), .B(n_517), .Y(n_676) );
AND2x2_ASAP7_75t_L g680 ( .A(n_507), .B(n_518), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_507), .B(n_556), .Y(n_693) );
AND2x2_ASAP7_75t_L g700 ( .A(n_507), .B(n_582), .Y(n_700) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .Y(n_507) );
INVx1_ASAP7_75t_SL g643 ( .A(n_516), .Y(n_643) );
AND2x2_ASAP7_75t_L g582 ( .A(n_517), .B(n_544), .Y(n_582) );
AND2x2_ASAP7_75t_L g596 ( .A(n_517), .B(n_551), .Y(n_596) );
AND2x2_ASAP7_75t_L g599 ( .A(n_517), .B(n_555), .Y(n_599) );
INVx1_ASAP7_75t_L g626 ( .A(n_517), .Y(n_626) );
INVx2_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g538 ( .A(n_518), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g697 ( .A1(n_528), .A2(n_574), .B(n_698), .C(n_699), .Y(n_697) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g604 ( .A(n_529), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_530), .B(n_547), .Y(n_562) );
AND2x2_ASAP7_75t_L g588 ( .A(n_530), .B(n_589), .Y(n_588) );
OAI21xp5_ASAP7_75t_SL g531 ( .A1(n_532), .A2(n_535), .B(n_539), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_533), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g559 ( .A(n_534), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_534), .B(n_555), .Y(n_600) );
AND2x2_ASAP7_75t_L g691 ( .A(n_534), .B(n_542), .Y(n_691) );
INVxp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g564 ( .A(n_538), .B(n_551), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_538), .B(n_549), .Y(n_565) );
OAI322xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_548), .A3(n_549), .B1(n_552), .B2(n_553), .C1(n_557), .C2(n_558), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_547), .Y(n_541) );
AND2x2_ASAP7_75t_L g652 ( .A(n_542), .B(n_564), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_542), .B(n_616), .Y(n_698) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g595 ( .A(n_544), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g661 ( .A(n_548), .B(n_574), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_549), .B(n_643), .Y(n_642) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_550), .B(n_582), .Y(n_639) );
AND2x2_ASAP7_75t_L g585 ( .A(n_551), .B(n_555), .Y(n_585) );
AND2x2_ASAP7_75t_L g593 ( .A(n_552), .B(n_594), .Y(n_593) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_552), .A2(n_631), .B(n_691), .C(n_692), .Y(n_690) );
AOI21xp33_ASAP7_75t_L g663 ( .A1(n_553), .A2(n_566), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_555), .B(n_582), .Y(n_622) );
AND2x2_ASAP7_75t_L g628 ( .A(n_555), .B(n_596), .Y(n_628) );
AND2x2_ASAP7_75t_L g662 ( .A(n_555), .B(n_564), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_556), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_SL g672 ( .A(n_556), .Y(n_672) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_560), .A2(n_588), .B1(n_590), .B2(n_595), .Y(n_587) );
OAI22xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_563), .B1(n_565), .B2(n_566), .Y(n_561) );
OAI22xp33_ASAP7_75t_L g597 ( .A1(n_562), .A2(n_598), .B1(n_600), .B2(n_601), .Y(n_597) );
INVxp67_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_567), .A2(n_669), .B1(n_671), .B2(n_673), .C(n_677), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_572), .B(n_576), .C(n_597), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
OR2x2_ASAP7_75t_L g638 ( .A(n_574), .B(n_591), .Y(n_638) );
INVx1_ASAP7_75t_L g689 ( .A(n_574), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g576 ( .A1(n_575), .A2(n_577), .B1(n_581), .B2(n_584), .C(n_587), .Y(n_576) );
INVx2_ASAP7_75t_SL g631 ( .A(n_575), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g696 ( .A(n_578), .Y(n_696) );
AND2x2_ASAP7_75t_L g620 ( .A(n_579), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g605 ( .A(n_580), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g667 ( .A(n_583), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_591), .B(n_693), .Y(n_692) );
CKINVDCx16_ASAP7_75t_R g591 ( .A(n_592), .Y(n_591) );
INVxp67_ASAP7_75t_L g636 ( .A(n_594), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g606 ( .A1(n_595), .A2(n_607), .B(n_609), .C(n_611), .Y(n_606) );
INVx1_ASAP7_75t_L g684 ( .A(n_598), .Y(n_684) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_602), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx2_ASAP7_75t_L g615 ( .A(n_605), .Y(n_615) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI222xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_618), .B1(n_619), .B2(n_622), .C1(n_623), .C2(n_625), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g651 ( .A(n_615), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_618), .B(n_672), .Y(n_671) );
NAND2xp33_ASAP7_75t_SL g649 ( .A(n_619), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g624 ( .A(n_621), .Y(n_624) );
AND2x2_ASAP7_75t_L g688 ( .A(n_621), .B(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g654 ( .A(n_624), .B(n_651), .Y(n_654) );
INVx1_ASAP7_75t_L g683 ( .A(n_625), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B(n_632), .C(n_637), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_631), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
AOI322xp5_ASAP7_75t_L g682 ( .A1(n_634), .A2(n_662), .A3(n_667), .B1(n_683), .B2(n_684), .C1(n_685), .C2(n_688), .Y(n_682) );
AND2x2_ASAP7_75t_L g669 ( .A(n_635), .B(n_670), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B1(n_640), .B2(n_642), .Y(n_637) );
INVxp33_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B1(n_649), .B2(n_652), .C(n_653), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NAND5xp2_ASAP7_75t_L g656 ( .A(n_657), .B(n_668), .C(n_682), .D(n_690), .E(n_694), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_662), .B(n_663), .Y(n_657) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVxp33_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_670), .A2(n_695), .B(n_696), .C(n_697), .Y(n_694) );
AOI31xp33_ASAP7_75t_L g677 ( .A1(n_672), .A2(n_678), .A3(n_679), .B(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g695 ( .A(n_693), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g709 ( .A(n_702), .Y(n_709) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI22x1_ASAP7_75t_SL g705 ( .A1(n_706), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_705) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g719 ( .A(n_718), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g734 ( .A(n_725), .Y(n_734) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_729), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
endmodule