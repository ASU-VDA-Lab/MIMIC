module fake_aes_7076_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
OR2x6_ASAP7_75t_L g3 ( .A(n_0), .B(n_1), .Y(n_3) );
BUFx6f_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_1), .B(n_2), .Y(n_6) );
BUFx2_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_5), .B(n_3), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
AOI21xp5_ASAP7_75t_SL g10 ( .A1(n_9), .A2(n_8), .B(n_7), .Y(n_10) );
NAND4xp25_ASAP7_75t_L g11 ( .A(n_9), .B(n_3), .C(n_2), .D(n_4), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
AOI22xp33_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_3), .B1(n_10), .B2(n_6), .Y(n_13) );
endmodule