module fake_jpeg_11662_n_453 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_453);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_453;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

NOR2xp67_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_58),
.Y(n_104)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_53),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_55),
.Y(n_148)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_57),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_64),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_19),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_61),
.B(n_84),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_19),
.B(n_0),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_70),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_1),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_79),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_75),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_37),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_88),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_3),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_37),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_17),
.Y(n_100)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_28),
.B(n_5),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_92),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_40),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g91 ( 
.A(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_6),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_40),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_100),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_72),
.B(n_42),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_113),
.C(n_32),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_51),
.A2(n_71),
.B1(n_65),
.B2(n_89),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_107),
.A2(n_112),
.B1(n_115),
.B2(n_125),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_34),
.B1(n_36),
.B2(n_28),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_42),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_62),
.A2(n_93),
.B1(n_85),
.B2(n_66),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_114),
.A2(n_135),
.B1(n_43),
.B2(n_45),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_68),
.A2(n_32),
.B1(n_43),
.B2(n_45),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_55),
.A2(n_32),
.B1(n_39),
.B2(n_38),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_82),
.A2(n_32),
.B1(n_38),
.B2(n_34),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_126),
.A2(n_47),
.B1(n_54),
.B2(n_77),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_74),
.A2(n_45),
.B1(n_43),
.B2(n_38),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_90),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_50),
.B(n_33),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_140),
.B(n_25),
.Y(n_182)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_49),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_142),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_59),
.B(n_25),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_149),
.B(n_137),
.C(n_117),
.Y(n_204)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_163),
.Y(n_199)
);

INVx6_ASAP7_75t_SL g153 ( 
.A(n_120),
.Y(n_153)
);

BUFx24_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_87),
.B1(n_63),
.B2(n_69),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_154),
.A2(n_162),
.B1(n_174),
.B2(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_98),
.B(n_41),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_159),
.Y(n_197)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_41),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

AND2x4_ASAP7_75t_SL g161 ( 
.A(n_101),
.B(n_81),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_178),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_129),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

AO22x1_ASAP7_75t_SL g169 ( 
.A1(n_101),
.A2(n_47),
.B1(n_80),
.B2(n_53),
.Y(n_169)
);

AO22x1_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_56),
.B1(n_57),
.B2(n_90),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_172),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_29),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_176),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_104),
.B(n_109),
.C(n_145),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_175),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_113),
.B(n_30),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_115),
.A2(n_76),
.B1(n_48),
.B2(n_45),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_130),
.B1(n_146),
.B2(n_96),
.Y(n_208)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_107),
.A2(n_43),
.B1(n_33),
.B2(n_36),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_91),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_180),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_139),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_185),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_182),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_91),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_188),
.B(n_191),
.Y(n_222)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_122),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_184),
.Y(n_227)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_190),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_100),
.A2(n_54),
.B1(n_42),
.B2(n_17),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_24),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_99),
.B(n_56),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_120),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_102),
.Y(n_217)
);

NAND2xp33_ASAP7_75t_SL g193 ( 
.A(n_169),
.B(n_105),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_194),
.B(n_202),
.Y(n_229)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_169),
.B(n_105),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_126),
.B1(n_125),
.B2(n_127),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_196),
.A2(n_213),
.B1(n_203),
.B2(n_211),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_208),
.B1(n_212),
.B2(n_215),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_191),
.A2(n_116),
.B(n_108),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_188),
.C(n_167),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_177),
.A2(n_146),
.B1(n_96),
.B2(n_131),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_149),
.A2(n_131),
.B1(n_127),
.B2(n_103),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_103),
.B1(n_128),
.B2(n_23),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_217),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_183),
.A2(n_108),
.B(n_120),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_194),
.B(n_193),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_197),
.A2(n_173),
.B1(n_176),
.B2(n_161),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_230),
.A2(n_241),
.B1(n_210),
.B2(n_221),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_231),
.B(n_237),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_201),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_232),
.Y(n_277)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_201),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_238),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_156),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_250),
.Y(n_261)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_203),
.A2(n_161),
.B1(n_152),
.B2(n_159),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_243),
.B(n_244),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_171),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_201),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_196),
.A2(n_152),
.B1(n_181),
.B2(n_161),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_246),
.A2(n_247),
.B(n_226),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_200),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_205),
.B(n_198),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_216),
.B(n_163),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_251),
.Y(n_273)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_205),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_255),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_164),
.C(n_158),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_178),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_217),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_198),
.B(n_155),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_258),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_257),
.A2(n_200),
.B1(n_211),
.B2(n_213),
.Y(n_264)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_259),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_229),
.A2(n_220),
.B(n_211),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_260),
.A2(n_278),
.B(n_236),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_271),
.B1(n_279),
.B2(n_232),
.Y(n_292)
);

AOI32xp33_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_246),
.A3(n_257),
.B1(n_248),
.B2(n_250),
.Y(n_267)
);

A2O1A1O1Ixp25_ASAP7_75t_L g301 ( 
.A1(n_267),
.A2(n_289),
.B(n_260),
.C(n_263),
.D(n_264),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_282),
.C(n_288),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_257),
.A2(n_210),
.B1(n_200),
.B2(n_179),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_233),
.A2(n_209),
.B1(n_195),
.B2(n_170),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_283),
.B1(n_232),
.B2(n_234),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_276),
.B(n_251),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_229),
.A2(n_247),
.B(n_246),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_233),
.A2(n_195),
.B1(n_170),
.B2(n_226),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_288),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_168),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_253),
.A2(n_151),
.B1(n_224),
.B2(n_227),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_235),
.A2(n_153),
.B(n_172),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_289),
.B(n_192),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_223),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_248),
.B1(n_241),
.B2(n_256),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_290),
.A2(n_295),
.B1(n_310),
.B2(n_315),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_292),
.A2(n_317),
.B1(n_242),
.B2(n_206),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_239),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_294),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_278),
.A2(n_263),
.B1(n_285),
.B2(n_267),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_245),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_259),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_308),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_286),
.Y(n_324)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_300),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_301),
.A2(n_304),
.B(n_305),
.Y(n_322)
);

AOI22x1_ASAP7_75t_L g302 ( 
.A1(n_271),
.A2(n_242),
.B1(n_230),
.B2(n_258),
.Y(n_302)
);

AOI22x1_ASAP7_75t_L g336 ( 
.A1(n_302),
.A2(n_184),
.B1(n_166),
.B2(n_207),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_303),
.B(n_318),
.Y(n_344)
);

OA21x2_ASAP7_75t_L g304 ( 
.A1(n_266),
.A2(n_242),
.B(n_252),
.Y(n_304)
);

OA21x2_ASAP7_75t_L g305 ( 
.A1(n_277),
.A2(n_242),
.B(n_249),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_306),
.Y(n_337)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_265),
.Y(n_307)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_309),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_285),
.A2(n_269),
.B1(n_272),
.B2(n_270),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_284),
.A2(n_240),
.B(n_238),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_311),
.B(n_314),
.Y(n_345)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_244),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_280),
.C(n_268),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_279),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_262),
.A2(n_242),
.B1(n_234),
.B2(n_206),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_287),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_316),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_224),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_292),
.A2(n_287),
.B1(n_286),
.B2(n_280),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_323),
.A2(n_330),
.B1(n_332),
.B2(n_305),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_329),
.C(n_346),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_325),
.B(n_160),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_326),
.A2(n_315),
.B1(n_305),
.B2(n_317),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_223),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_341),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_227),
.C(n_187),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_302),
.A2(n_219),
.B1(n_150),
.B2(n_128),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_SL g331 ( 
.A(n_316),
.B(n_165),
.C(n_44),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_219),
.C(n_30),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_306),
.A2(n_219),
.B1(n_228),
.B2(n_207),
.Y(n_332)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_336),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_299),
.B(n_185),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_308),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_343),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_290),
.B(n_165),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_347),
.A2(n_349),
.B1(n_354),
.B2(n_359),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_332),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_348),
.B(n_160),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_337),
.A2(n_301),
.B(n_322),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_350),
.A2(n_141),
.B(n_123),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_324),
.B(n_295),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_351),
.B(n_352),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_341),
.B(n_310),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_354),
.A2(n_359),
.B1(n_363),
.B2(n_160),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_344),
.B(n_313),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_352),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_334),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_358),
.B(n_362),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_323),
.A2(n_340),
.B1(n_304),
.B2(n_330),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_333),
.A2(n_311),
.B1(n_304),
.B2(n_300),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_361),
.A2(n_365),
.B1(n_339),
.B2(n_331),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_320),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_345),
.A2(n_337),
.B1(n_335),
.B2(n_333),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_228),
.Y(n_364)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_364),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_325),
.A2(n_228),
.B1(n_189),
.B2(n_157),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_367),
.B(n_329),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_336),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_368),
.B(n_369),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_319),
.Y(n_369)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_321),
.B(n_7),
.C(n_8),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_328),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_377),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_388),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_383),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_375),
.B(n_386),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_346),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_327),
.C(n_336),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_380),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_338),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_339),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_384),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_382),
.A2(n_387),
.B1(n_364),
.B2(n_348),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_353),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_366),
.Y(n_384)
);

AO22x1_ASAP7_75t_L g398 ( 
.A1(n_385),
.A2(n_355),
.B1(n_389),
.B2(n_360),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_347),
.A2(n_27),
.B1(n_24),
.B2(n_29),
.Y(n_386)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_390),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_353),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_374),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_360),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_396),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_351),
.C(n_350),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_398),
.B(n_372),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_378),
.A2(n_361),
.B(n_27),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_141),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_389),
.A2(n_97),
.B(n_123),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_401),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_23),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_118),
.C(n_44),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_404),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_118),
.C(n_148),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_406),
.B(n_410),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_408),
.A2(n_405),
.B(n_400),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_388),
.C(n_385),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_387),
.Y(n_412)
);

INVxp33_ASAP7_75t_L g431 ( 
.A(n_412),
.Y(n_431)
);

OAI321xp33_ASAP7_75t_L g413 ( 
.A1(n_402),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_413),
.A2(n_419),
.B1(n_403),
.B2(n_404),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_148),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_414),
.B(n_415),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_7),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_391),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_416),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_398),
.B(n_148),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_412),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_422),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_418),
.A2(n_405),
.B1(n_390),
.B2(n_391),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_421),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_97),
.C(n_57),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_423),
.B(n_428),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_17),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_42),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_409),
.B(n_42),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_429),
.A2(n_430),
.B(n_13),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_417),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_431),
.A2(n_86),
.B(n_11),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_432),
.A2(n_434),
.B(n_438),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_10),
.Y(n_433)
);

AOI21x1_ASAP7_75t_L g444 ( 
.A1(n_433),
.A2(n_435),
.B(n_425),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_431),
.A2(n_10),
.B(n_11),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_436),
.Y(n_445)
);

O2A1O1Ixp33_ASAP7_75t_SL g438 ( 
.A1(n_422),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_13),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_441),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_439),
.B(n_427),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_443),
.B(n_444),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_442),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_447),
.A2(n_437),
.B(n_426),
.Y(n_449)
);

O2A1O1Ixp33_ASAP7_75t_SL g451 ( 
.A1(n_449),
.A2(n_450),
.B(n_446),
.C(n_13),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_448),
.A2(n_445),
.B(n_423),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_13),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_452),
.A2(n_14),
.B(n_375),
.Y(n_453)
);


endmodule