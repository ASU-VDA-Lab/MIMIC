module fake_jpeg_1644_n_46 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_46);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_32;

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_2),
.B(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_5),
.B(n_16),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_SL g27 ( 
.A1(n_4),
.A2(n_9),
.B(n_10),
.Y(n_27)
);

HAxp5_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_1),
.CON(n_28),
.SN(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_7),
.A2(n_11),
.B(n_2),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_12),
.B1(n_13),
.B2(n_18),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_39)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_36),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_32),
.B1(n_22),
.B2(n_23),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_40),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_36),
.B(n_24),
.C(n_39),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_21),
.B(n_28),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_23),
.Y(n_46)
);


endmodule