module fake_jpeg_14838_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_40),
.Y(n_68)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_27),
.B1(n_18),
.B2(n_32),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_61),
.B1(n_63),
.B2(n_29),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_43),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_27),
.B1(n_18),
.B2(n_17),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_53),
.B1(n_56),
.B2(n_67),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_17),
.B1(n_33),
.B2(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_16),
.B1(n_33),
.B2(n_21),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_26),
.B(n_30),
.Y(n_62)
);

OR2x4_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_24),
.B1(n_21),
.B2(n_16),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_24),
.B1(n_21),
.B2(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_22),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_47),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_70),
.A2(n_73),
.B(n_74),
.Y(n_115)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_28),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_41),
.B1(n_28),
.B2(n_43),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_77),
.A2(n_87),
.B1(n_89),
.B2(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_90),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_39),
.B1(n_44),
.B2(n_40),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_82),
.B1(n_92),
.B2(n_51),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_96),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_22),
.B1(n_30),
.B2(n_26),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_43),
.B1(n_12),
.B2(n_15),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_83),
.A2(n_84),
.B1(n_86),
.B2(n_46),
.Y(n_117)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_45),
.B1(n_34),
.B2(n_29),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_45),
.B1(n_34),
.B2(n_29),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_42),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_45),
.B1(n_42),
.B2(n_34),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_11),
.B(n_15),
.Y(n_107)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_53),
.B(n_19),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_42),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_102),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_45),
.B1(n_29),
.B2(n_34),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_66),
.B(n_13),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_42),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_50),
.Y(n_134)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_107),
.A2(n_113),
.B1(n_117),
.B2(n_92),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_42),
.C(n_20),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_128),
.C(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_51),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_119),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_46),
.A3(n_20),
.B1(n_23),
.B2(n_31),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_70),
.B(n_23),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_20),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_133),
.Y(n_137)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_94),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_31),
.C(n_19),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_80),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVxp33_ASAP7_75t_SL g131 ( 
.A(n_77),
.Y(n_131)
);

AO21x2_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_92),
.B(n_89),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_0),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_125),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_139),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_102),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_143),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_142),
.B(n_148),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_88),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_72),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_147),
.C(n_165),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_72),
.B1(n_71),
.B2(n_84),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_158),
.B1(n_113),
.B2(n_128),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_90),
.C(n_88),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_149),
.B(n_151),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_161),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_111),
.B(n_91),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_104),
.B1(n_95),
.B2(n_75),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_160),
.B1(n_126),
.B2(n_121),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_80),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_76),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_98),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_167),
.B1(n_164),
.B2(n_124),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_92),
.B1(n_103),
.B2(n_14),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_111),
.B1(n_124),
.B2(n_121),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_122),
.A2(n_14),
.B1(n_11),
.B2(n_10),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_132),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_19),
.C(n_31),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_0),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_137),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_0),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_133),
.B(n_107),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_166),
.B(n_137),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_171),
.A2(n_5),
.B(n_6),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_172),
.A2(n_178),
.B1(n_196),
.B2(n_157),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_177),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_179),
.C(n_190),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_163),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_110),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_147),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_185),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_138),
.C(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_193),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_132),
.C(n_127),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_199),
.Y(n_202)
);

OAI21x1_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_10),
.B(n_9),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_195),
.B(n_1),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_196),
.B(n_198),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_197),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_130),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_136),
.B(n_127),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_172),
.A2(n_154),
.B1(n_157),
.B2(n_167),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_213),
.B1(n_218),
.B2(n_228),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_220),
.B(n_223),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_146),
.Y(n_216)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_SL g217 ( 
.A1(n_201),
.A2(n_165),
.B(n_157),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_225),
.C(n_168),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_157),
.B1(n_130),
.B2(n_3),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_191),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_186),
.A2(n_1),
.B(n_2),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_199),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_2),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_173),
.A2(n_3),
.B(n_4),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_226),
.B(n_227),
.Y(n_237)
);

XNOR2x1_ASAP7_75t_L g225 ( 
.A(n_179),
.B(n_3),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_173),
.A2(n_3),
.B(n_4),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_171),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_8),
.Y(n_229)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_250),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_176),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_241),
.C(n_243),
.Y(n_261)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_236),
.B(n_239),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_SL g262 ( 
.A(n_238),
.B(n_246),
.C(n_225),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_214),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_194),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_170),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_245),
.C(n_248),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_210),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_181),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_188),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_249),
.B(n_253),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_192),
.C(n_189),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_224),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_180),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_270),
.C(n_252),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_228),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_257),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_248),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_260),
.Y(n_278)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_226),
.C(n_244),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_174),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_222),
.B1(n_213),
.B2(n_218),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_227),
.B(n_203),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_266),
.A2(n_268),
.B(n_237),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_203),
.B(n_217),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_209),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_235),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_250),
.B(n_229),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_273),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_254),
.Y(n_298)
);

OA21x2_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_238),
.B(n_171),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_245),
.Y(n_293)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_282),
.C(n_262),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_241),
.C(n_232),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_261),
.C(n_270),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_283),
.A2(n_240),
.B1(n_204),
.B2(n_169),
.Y(n_299)
);

AO22x1_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_207),
.B1(n_171),
.B2(n_215),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_288),
.Y(n_302)
);

AO221x1_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_193),
.B1(n_211),
.B2(n_197),
.C(n_169),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_255),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_207),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_287),
.A2(n_265),
.B1(n_255),
.B2(n_267),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_292),
.B1(n_301),
.B2(n_303),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_294),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_296),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_276),
.A2(n_258),
.B(n_264),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_264),
.B(n_267),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_282),
.A2(n_220),
.B(n_221),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_285),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_269),
.B(n_223),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_283),
.B(n_285),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_280),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_311),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_290),
.B(n_280),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_308),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_278),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_312),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_288),
.B1(n_274),
.B2(n_275),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_289),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_296),
.B(n_303),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_320),
.B(n_275),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_311),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_316),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_297),
.C(n_298),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_292),
.C(n_309),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_289),
.B(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_323),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_320),
.A2(n_211),
.B(n_279),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_319),
.C(n_318),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_321),
.B(n_281),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_326),
.B(n_204),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

AOI322xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_219),
.C1(n_223),
.C2(n_328),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_223),
.Y(n_331)
);


endmodule