module real_aes_90_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_788, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_788;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g176 ( .A(n_0), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_1), .B(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_2), .B(n_182), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_3), .B(n_179), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_4), .A2(n_45), .B1(n_772), .B2(n_773), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_4), .Y(n_772) );
INVx1_ASAP7_75t_L g142 ( .A(n_5), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_6), .B(n_182), .Y(n_204) );
NAND2xp33_ASAP7_75t_SL g162 ( .A(n_7), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g133 ( .A(n_8), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_9), .Y(n_784) );
CKINVDCx16_ASAP7_75t_R g781 ( .A(n_10), .Y(n_781) );
AND2x2_ASAP7_75t_L g202 ( .A(n_11), .B(n_185), .Y(n_202) );
AND2x2_ASAP7_75t_L g472 ( .A(n_12), .B(n_158), .Y(n_472) );
AND2x2_ASAP7_75t_L g523 ( .A(n_13), .B(n_213), .Y(n_523) );
INVx2_ASAP7_75t_L g136 ( .A(n_14), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_15), .B(n_179), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_16), .Y(n_111) );
NOR3xp33_ASAP7_75t_L g779 ( .A(n_16), .B(n_780), .C(n_782), .Y(n_779) );
AOI221x1_ASAP7_75t_L g154 ( .A1(n_17), .A2(n_155), .B1(n_157), .B2(n_158), .C(n_161), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_18), .B(n_182), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_19), .B(n_182), .Y(n_528) );
INVx1_ASAP7_75t_L g115 ( .A(n_20), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_21), .A2(n_91), .B1(n_137), .B2(n_182), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_22), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_23), .A2(n_157), .B(n_206), .Y(n_205) );
AOI221xp5_ASAP7_75t_SL g249 ( .A1(n_24), .A2(n_37), .B1(n_157), .B2(n_182), .C(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_25), .B(n_177), .Y(n_207) );
OR2x2_ASAP7_75t_L g135 ( .A(n_26), .B(n_90), .Y(n_135) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_26), .A2(n_90), .B(n_136), .Y(n_160) );
INVxp67_ASAP7_75t_L g153 ( .A(n_27), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_28), .B(n_179), .Y(n_244) );
AND2x2_ASAP7_75t_L g196 ( .A(n_29), .B(n_184), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_30), .A2(n_157), .B(n_175), .Y(n_174) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_31), .A2(n_158), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_32), .B(n_179), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_33), .A2(n_157), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_34), .B(n_179), .Y(n_504) );
AND2x2_ASAP7_75t_L g144 ( .A(n_35), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g148 ( .A(n_35), .Y(n_148) );
AND2x2_ASAP7_75t_L g163 ( .A(n_35), .B(n_142), .Y(n_163) );
OR2x6_ASAP7_75t_L g113 ( .A(n_36), .B(n_114), .Y(n_113) );
INVxp67_ASAP7_75t_L g782 ( .A(n_36), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_38), .B(n_182), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_39), .A2(n_83), .B1(n_146), .B2(n_157), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_40), .B(n_179), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_41), .A2(n_50), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_41), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_42), .B(n_182), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_43), .B(n_177), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_44), .A2(n_157), .B(n_468), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_45), .Y(n_773) );
AND2x2_ASAP7_75t_L g183 ( .A(n_46), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_47), .B(n_177), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_48), .B(n_184), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_49), .B(n_182), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_50), .Y(n_750) );
INVx1_ASAP7_75t_L g140 ( .A(n_51), .Y(n_140) );
INVx1_ASAP7_75t_L g167 ( .A(n_51), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_52), .B(n_179), .Y(n_470) );
AND2x2_ASAP7_75t_L g482 ( .A(n_53), .B(n_184), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_54), .B(n_182), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_55), .B(n_177), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_56), .B(n_177), .Y(n_503) );
AND2x2_ASAP7_75t_L g225 ( .A(n_57), .B(n_184), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_58), .B(n_182), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_59), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_60), .B(n_182), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_61), .A2(n_157), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_62), .B(n_177), .Y(n_223) );
AND2x2_ASAP7_75t_SL g245 ( .A(n_63), .B(n_185), .Y(n_245) );
XNOR2xp5_ASAP7_75t_L g748 ( .A(n_64), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g534 ( .A(n_65), .B(n_185), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_66), .A2(n_157), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_67), .B(n_179), .Y(n_208) );
AND2x2_ASAP7_75t_SL g217 ( .A(n_68), .B(n_213), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_69), .B(n_177), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_70), .B(n_177), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_71), .A2(n_93), .B1(n_146), .B2(n_157), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_72), .B(n_179), .Y(n_531) );
INVx1_ASAP7_75t_L g145 ( .A(n_73), .Y(n_145) );
INVx1_ASAP7_75t_L g169 ( .A(n_73), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_74), .B(n_177), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_75), .A2(n_157), .B(n_486), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_76), .A2(n_157), .B(n_460), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_77), .A2(n_157), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g506 ( .A(n_78), .B(n_185), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_79), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_80), .B(n_184), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_81), .A2(n_85), .B1(n_137), .B2(n_182), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_82), .B(n_182), .Y(n_224) );
INVx1_ASAP7_75t_L g116 ( .A(n_84), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_84), .B(n_115), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_86), .B(n_177), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_87), .B(n_177), .Y(n_252) );
AND2x2_ASAP7_75t_L g463 ( .A(n_88), .B(n_213), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_89), .A2(n_157), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_92), .B(n_179), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_94), .A2(n_157), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_95), .B(n_179), .Y(n_461) );
OAI22x1_ASAP7_75t_R g769 ( .A1(n_96), .A2(n_770), .B1(n_771), .B2(n_774), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_96), .Y(n_774) );
INVxp67_ASAP7_75t_L g156 ( .A(n_97), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_98), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_99), .B(n_179), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_100), .A2(n_157), .B(n_242), .Y(n_241) );
BUFx2_ASAP7_75t_L g533 ( .A(n_101), .Y(n_533) );
BUFx2_ASAP7_75t_L g120 ( .A(n_102), .Y(n_120) );
AOI21xp33_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_775), .B(n_783), .Y(n_103) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_121), .B(n_761), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g105 ( .A(n_106), .B(n_118), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_SL g763 ( .A1(n_107), .A2(n_764), .B(n_767), .Y(n_763) );
NOR2xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_117), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_R g766 ( .A(n_110), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x6_ASAP7_75t_SL g449 ( .A(n_111), .B(n_113), .Y(n_449) );
OR2x6_ASAP7_75t_SL g747 ( .A(n_111), .B(n_112), .Y(n_747) );
OR2x2_ASAP7_75t_L g760 ( .A(n_111), .B(n_113), .Y(n_760) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_120), .Y(n_762) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_748), .B(n_752), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22x1_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_448), .B1(n_450), .B2(n_745), .Y(n_123) );
OAI22x1_ASAP7_75t_L g767 ( .A1(n_124), .A2(n_125), .B1(n_768), .B2(n_769), .Y(n_767) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OA22x2_ASAP7_75t_L g754 ( .A1(n_125), .A2(n_448), .B1(n_451), .B2(n_755), .Y(n_754) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_325), .Y(n_125) );
NOR4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_268), .C(n_307), .D(n_314), .Y(n_126) );
OAI221xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_186), .B1(n_226), .B2(n_235), .C(n_254), .Y(n_127) );
OR2x2_ASAP7_75t_L g398 ( .A(n_128), .B(n_260), .Y(n_398) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g313 ( .A(n_129), .B(n_238), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_129), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_SL g378 ( .A(n_129), .B(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_170), .Y(n_129) );
AND2x4_ASAP7_75t_SL g237 ( .A(n_130), .B(n_238), .Y(n_237) );
INVx3_ASAP7_75t_L g259 ( .A(n_130), .Y(n_259) );
AND2x2_ASAP7_75t_L g294 ( .A(n_130), .B(n_267), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_130), .B(n_171), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_130), .B(n_261), .Y(n_346) );
OR2x2_ASAP7_75t_L g424 ( .A(n_130), .B(n_238), .Y(n_424) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_154), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_137), .B1(n_146), .B2(n_152), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_134), .B(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_134), .B(n_156), .Y(n_155) );
NOR3xp33_ASAP7_75t_L g161 ( .A(n_134), .B(n_162), .C(n_164), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_134), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_134), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_134), .A2(n_493), .B(n_494), .Y(n_492) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_135), .B(n_136), .Y(n_185) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_143), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g151 ( .A(n_140), .B(n_142), .Y(n_151) );
AND2x4_ASAP7_75t_L g179 ( .A(n_140), .B(n_168), .Y(n_179) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x6_ASAP7_75t_L g157 ( .A(n_144), .B(n_151), .Y(n_157) );
INVx2_ASAP7_75t_L g150 ( .A(n_145), .Y(n_150) );
AND2x6_ASAP7_75t_L g177 ( .A(n_145), .B(n_166), .Y(n_177) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
NOR2x1p5_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g499 ( .A(n_158), .Y(n_499) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21x1_ASAP7_75t_L g172 ( .A1(n_159), .A2(n_173), .B(n_183), .Y(n_172) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_159), .A2(n_466), .B(n_472), .Y(n_465) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx4f_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
INVx5_ASAP7_75t_L g180 ( .A(n_163), .Y(n_180) );
AND2x4_ASAP7_75t_L g182 ( .A(n_163), .B(n_165), .Y(n_182) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_166), .B(n_168), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g246 ( .A(n_171), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_171), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g272 ( .A(n_171), .Y(n_272) );
OR2x2_ASAP7_75t_L g277 ( .A(n_171), .B(n_261), .Y(n_277) );
AND2x2_ASAP7_75t_L g290 ( .A(n_171), .B(n_248), .Y(n_290) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_171), .Y(n_293) );
INVx1_ASAP7_75t_L g305 ( .A(n_171), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_171), .B(n_259), .Y(n_370) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_181), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_178), .B(n_180), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_177), .B(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_180), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_180), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_180), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_180), .A2(n_243), .B(n_244), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_180), .A2(n_251), .B(n_252), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_180), .A2(n_461), .B(n_462), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_180), .A2(n_469), .B(n_470), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_180), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_180), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_180), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_180), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_180), .A2(n_531), .B(n_532), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_184), .Y(n_195) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_184), .A2(n_249), .B(n_253), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_184), .A2(n_458), .B(n_459), .Y(n_457) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_184), .A2(n_476), .B(n_477), .Y(n_475) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_187), .B(n_197), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g234 ( .A(n_188), .B(n_218), .Y(n_234) );
AND2x4_ASAP7_75t_L g264 ( .A(n_188), .B(n_201), .Y(n_264) );
INVx2_ASAP7_75t_L g298 ( .A(n_188), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_188), .B(n_218), .Y(n_356) );
AND2x2_ASAP7_75t_L g403 ( .A(n_188), .B(n_232), .Y(n_403) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_195), .B(n_196), .Y(n_188) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_189), .A2(n_195), .B(n_196), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_194), .Y(n_189) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_195), .A2(n_219), .B(n_225), .Y(n_218) );
AOI21x1_ASAP7_75t_L g516 ( .A1(n_195), .A2(n_517), .B(n_523), .Y(n_516) );
AOI222xp33_ASAP7_75t_L g391 ( .A1(n_197), .A2(n_263), .B1(n_306), .B2(n_366), .C1(n_392), .C2(n_394), .Y(n_391) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_209), .Y(n_198) );
AND2x2_ASAP7_75t_L g310 ( .A(n_199), .B(n_230), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_199), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g439 ( .A(n_199), .B(n_279), .Y(n_439) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_200), .A2(n_270), .B(n_274), .Y(n_269) );
AND2x2_ASAP7_75t_L g350 ( .A(n_200), .B(n_233), .Y(n_350) );
OR2x2_ASAP7_75t_L g375 ( .A(n_200), .B(n_234), .Y(n_375) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx5_ASAP7_75t_L g229 ( .A(n_201), .Y(n_229) );
AND2x2_ASAP7_75t_L g316 ( .A(n_201), .B(n_298), .Y(n_316) );
AND2x2_ASAP7_75t_L g342 ( .A(n_201), .B(n_218), .Y(n_342) );
OR2x2_ASAP7_75t_L g345 ( .A(n_201), .B(n_232), .Y(n_345) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_201), .Y(n_363) );
AND2x4_ASAP7_75t_SL g420 ( .A(n_201), .B(n_297), .Y(n_420) );
OR2x2_ASAP7_75t_L g429 ( .A(n_201), .B(n_256), .Y(n_429) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
INVx1_ASAP7_75t_L g262 ( .A(n_209), .Y(n_262) );
AOI221xp5_ASAP7_75t_SL g380 ( .A1(n_209), .A2(n_264), .B1(n_381), .B2(n_383), .C(n_384), .Y(n_380) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_218), .Y(n_209) );
OR2x2_ASAP7_75t_L g319 ( .A(n_210), .B(n_289), .Y(n_319) );
OR2x2_ASAP7_75t_L g329 ( .A(n_210), .B(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g355 ( .A(n_210), .B(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_L g361 ( .A(n_210), .B(n_280), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_210), .B(n_344), .Y(n_373) );
INVx2_ASAP7_75t_L g386 ( .A(n_210), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_210), .B(n_264), .Y(n_407) );
AND2x2_ASAP7_75t_L g411 ( .A(n_210), .B(n_233), .Y(n_411) );
AND2x2_ASAP7_75t_L g419 ( .A(n_210), .B(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g232 ( .A(n_211), .Y(n_232) );
AOI21x1_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_214), .B(n_217), .Y(n_211) );
INVx2_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_213), .A2(n_240), .B(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_213), .A2(n_528), .B(n_529), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_218), .B(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g263 ( .A(n_218), .B(n_232), .Y(n_263) );
INVx2_ASAP7_75t_L g280 ( .A(n_218), .Y(n_280) );
AND2x4_ASAP7_75t_L g297 ( .A(n_218), .B(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_218), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_230), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g409 ( .A(n_228), .B(n_231), .Y(n_409) );
AND2x4_ASAP7_75t_L g255 ( .A(n_229), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g296 ( .A(n_229), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g323 ( .A(n_229), .B(n_263), .Y(n_323) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
AND2x2_ASAP7_75t_L g427 ( .A(n_231), .B(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g279 ( .A(n_232), .B(n_280), .Y(n_279) );
OAI21xp5_ASAP7_75t_SL g299 ( .A1(n_233), .A2(n_300), .B(n_306), .Y(n_299) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_246), .Y(n_236) );
INVx1_ASAP7_75t_SL g353 ( .A(n_237), .Y(n_353) );
AND2x2_ASAP7_75t_L g383 ( .A(n_237), .B(n_293), .Y(n_383) );
AND2x4_ASAP7_75t_L g394 ( .A(n_237), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g260 ( .A(n_238), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g267 ( .A(n_238), .Y(n_267) );
AND2x4_ASAP7_75t_L g273 ( .A(n_238), .B(n_259), .Y(n_273) );
INVx2_ASAP7_75t_L g284 ( .A(n_238), .Y(n_284) );
INVx1_ASAP7_75t_L g333 ( .A(n_238), .Y(n_333) );
OR2x2_ASAP7_75t_L g354 ( .A(n_238), .B(n_338), .Y(n_354) );
OR2x2_ASAP7_75t_L g368 ( .A(n_238), .B(n_248), .Y(n_368) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_238), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_238), .B(n_290), .Y(n_440) );
OR2x6_ASAP7_75t_L g238 ( .A(n_239), .B(n_245), .Y(n_238) );
INVx1_ASAP7_75t_L g285 ( .A(n_246), .Y(n_285) );
AND2x2_ASAP7_75t_L g418 ( .A(n_246), .B(n_284), .Y(n_418) );
AND2x2_ASAP7_75t_L g443 ( .A(n_246), .B(n_273), .Y(n_443) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g261 ( .A(n_248), .Y(n_261) );
BUFx3_ASAP7_75t_L g303 ( .A(n_248), .Y(n_303) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_248), .Y(n_330) );
INVx1_ASAP7_75t_L g339 ( .A(n_248), .Y(n_339) );
AOI33xp33_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_257), .A3(n_262), .B1(n_263), .B2(n_264), .B3(n_265), .Y(n_254) );
AOI21x1_ASAP7_75t_SL g357 ( .A1(n_255), .A2(n_279), .B(n_341), .Y(n_357) );
INVx2_ASAP7_75t_L g387 ( .A(n_255), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_255), .B(n_386), .Y(n_393) );
AND2x2_ASAP7_75t_L g341 ( .A(n_256), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_L g304 ( .A(n_259), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g405 ( .A(n_260), .Y(n_405) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_261), .Y(n_395) );
OAI32xp33_ASAP7_75t_L g444 ( .A1(n_262), .A2(n_264), .A3(n_440), .B1(n_445), .B2(n_447), .Y(n_444) );
AND2x2_ASAP7_75t_L g362 ( .A(n_263), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_SL g352 ( .A(n_264), .Y(n_352) );
AND2x2_ASAP7_75t_L g417 ( .A(n_264), .B(n_361), .Y(n_417) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI221xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_278), .B1(n_281), .B2(n_295), .C(n_299), .Y(n_268) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_272), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_273), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_273), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_273), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g322 ( .A(n_277), .Y(n_322) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NOR3xp33_ASAP7_75t_L g281 ( .A(n_282), .B(n_286), .C(n_291), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_283), .A2(n_345), .B1(n_385), .B2(n_388), .Y(n_384) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g288 ( .A(n_284), .Y(n_288) );
NOR2x1p5_ASAP7_75t_L g302 ( .A(n_284), .B(n_303), .Y(n_302) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OAI322xp33_ASAP7_75t_L g351 ( .A1(n_287), .A2(n_329), .A3(n_352), .B1(n_353), .B2(n_354), .C1(n_355), .C2(n_357), .Y(n_351) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g307 ( .A1(n_289), .A2(n_308), .B(n_309), .C(n_311), .Y(n_307) );
OR2x2_ASAP7_75t_L g399 ( .A(n_289), .B(n_353), .Y(n_399) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g306 ( .A(n_290), .B(n_294), .Y(n_306) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g312 ( .A(n_296), .B(n_313), .Y(n_312) );
INVx3_ASAP7_75t_SL g344 ( .A(n_297), .Y(n_344) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_301), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_SL g348 ( .A(n_304), .Y(n_348) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_305), .Y(n_390) );
OR2x6_ASAP7_75t_SL g445 ( .A(n_308), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AOI211xp5_ASAP7_75t_L g435 ( .A1(n_313), .A2(n_436), .B(n_437), .C(n_444), .Y(n_435) );
O2A1O1Ixp33_ASAP7_75t_SL g314 ( .A1(n_315), .A2(n_317), .B(n_320), .C(n_324), .Y(n_314) );
OAI211xp5_ASAP7_75t_SL g326 ( .A1(n_315), .A2(n_327), .B(n_334), .C(n_358), .Y(n_326) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
NOR3xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_371), .C(n_415), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_330), .Y(n_422) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g377 ( .A(n_333), .Y(n_377) );
NOR3xp33_ASAP7_75t_SL g334 ( .A(n_335), .B(n_347), .C(n_351), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_340), .B1(n_343), .B2(n_346), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g379 ( .A(n_339), .Y(n_379) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_339), .Y(n_446) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_SL g432 ( .A(n_345), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
OR2x2_ASAP7_75t_L g382 ( .A(n_348), .B(n_368), .Y(n_382) );
OR2x2_ASAP7_75t_L g433 ( .A(n_348), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g431 ( .A(n_356), .Y(n_431) );
OR2x2_ASAP7_75t_L g447 ( .A(n_356), .B(n_386), .Y(n_447) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B(n_364), .Y(n_358) );
OAI31xp33_ASAP7_75t_L g372 ( .A1(n_359), .A2(n_373), .A3(n_374), .B(n_376), .Y(n_372) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g404 ( .A(n_369), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND4xp25_ASAP7_75t_SL g371 ( .A(n_372), .B(n_380), .C(n_391), .D(n_396), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .B1(n_404), .B2(n_406), .C(n_408), .Y(n_396) );
NAND2xp33_ASAP7_75t_SL g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g441 ( .A(n_400), .Y(n_441) );
AND2x2_ASAP7_75t_SL g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B(n_412), .Y(n_408) );
INVx1_ASAP7_75t_L g436 ( .A(n_410), .Y(n_436) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_416), .B(n_435), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_419), .B2(n_421), .C(n_425), .Y(n_416) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
AOI21xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_430), .B(n_433), .Y(n_425) );
INVxp33_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B1(n_441), .B2(n_442), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
CKINVDCx11_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
INVx3_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
AND2x4_ASAP7_75t_SL g451 ( .A(n_452), .B(n_641), .Y(n_451) );
NOR3xp33_ASAP7_75t_SL g452 ( .A(n_453), .B(n_550), .C(n_582), .Y(n_452) );
OAI221xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_478), .B1(n_507), .B2(n_524), .C(n_535), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_464), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g513 ( .A(n_456), .B(n_465), .Y(n_513) );
INVx4_ASAP7_75t_L g541 ( .A(n_456), .Y(n_541) );
AND2x4_ASAP7_75t_SL g581 ( .A(n_456), .B(n_515), .Y(n_581) );
BUFx2_ASAP7_75t_L g591 ( .A(n_456), .Y(n_591) );
NOR2x1_ASAP7_75t_L g657 ( .A(n_456), .B(n_596), .Y(n_657) );
AND2x2_ASAP7_75t_L g666 ( .A(n_456), .B(n_594), .Y(n_666) );
OR2x2_ASAP7_75t_L g674 ( .A(n_456), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g700 ( .A(n_456), .B(n_539), .Y(n_700) );
AND2x4_ASAP7_75t_L g719 ( .A(n_456), .B(n_720), .Y(n_719) );
OR2x6_ASAP7_75t_L g456 ( .A(n_457), .B(n_463), .Y(n_456) );
INVx2_ASAP7_75t_SL g632 ( .A(n_464), .Y(n_632) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_473), .Y(n_464) );
AND2x2_ASAP7_75t_L g539 ( .A(n_465), .B(n_516), .Y(n_539) );
INVx2_ASAP7_75t_L g566 ( .A(n_465), .Y(n_566) );
INVx2_ASAP7_75t_L g596 ( .A(n_465), .Y(n_596) );
AND2x2_ASAP7_75t_L g610 ( .A(n_465), .B(n_515), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .Y(n_466) );
AND2x2_ASAP7_75t_L g540 ( .A(n_473), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g563 ( .A(n_473), .Y(n_563) );
BUFx3_ASAP7_75t_L g577 ( .A(n_473), .Y(n_577) );
AND2x2_ASAP7_75t_L g606 ( .A(n_473), .B(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
AND2x4_ASAP7_75t_L g511 ( .A(n_474), .B(n_475), .Y(n_511) );
INVx1_ASAP7_75t_L g612 ( .A(n_478), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_489), .Y(n_478) );
OR2x2_ASAP7_75t_L g723 ( .A(n_479), .B(n_524), .Y(n_723) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g579 ( .A(n_480), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_480), .B(n_489), .Y(n_640) );
OR2x2_ASAP7_75t_L g738 ( .A(n_480), .B(n_660), .Y(n_738) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g549 ( .A(n_481), .B(n_525), .Y(n_549) );
OR2x2_ASAP7_75t_SL g559 ( .A(n_481), .B(n_560), .Y(n_559) );
INVx4_ASAP7_75t_L g570 ( .A(n_481), .Y(n_570) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_481), .Y(n_621) );
NAND2x1_ASAP7_75t_L g627 ( .A(n_481), .B(n_526), .Y(n_627) );
AND2x2_ASAP7_75t_L g652 ( .A(n_481), .B(n_491), .Y(n_652) );
OR2x2_ASAP7_75t_L g673 ( .A(n_481), .B(n_556), .Y(n_673) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g568 ( .A(n_489), .Y(n_568) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_489), .A2(n_662), .B(n_665), .C(n_667), .Y(n_661) );
AND2x2_ASAP7_75t_L g734 ( .A(n_489), .B(n_510), .Y(n_734) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_498), .Y(n_489) );
INVx1_ASAP7_75t_L g601 ( .A(n_490), .Y(n_601) );
AND2x2_ASAP7_75t_L g671 ( .A(n_490), .B(n_526), .Y(n_671) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g545 ( .A(n_491), .Y(n_545) );
OR2x2_ASAP7_75t_L g560 ( .A(n_491), .B(n_526), .Y(n_560) );
INVx1_ASAP7_75t_L g576 ( .A(n_491), .Y(n_576) );
AND2x2_ASAP7_75t_L g588 ( .A(n_491), .B(n_498), .Y(n_588) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_491), .Y(n_694) );
NOR2x1_ASAP7_75t_SL g525 ( .A(n_498), .B(n_526), .Y(n_525) );
AO21x1_ASAP7_75t_SL g498 ( .A1(n_499), .A2(n_500), .B(n_506), .Y(n_498) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_499), .A2(n_500), .B(n_506), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_505), .Y(n_500) );
INVxp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_512), .Y(n_508) );
OR2x2_ASAP7_75t_L g658 ( .A(n_509), .B(n_593), .Y(n_658) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_510), .B(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g740 ( .A(n_510), .B(n_637), .Y(n_740) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g585 ( .A(n_511), .B(n_566), .Y(n_585) );
AND2x2_ASAP7_75t_L g681 ( .A(n_511), .B(n_594), .Y(n_681) );
INVx1_ASAP7_75t_L g598 ( .A(n_512), .Y(n_598) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g648 ( .A(n_513), .Y(n_648) );
INVx2_ASAP7_75t_L g615 ( .A(n_514), .Y(n_615) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g565 ( .A(n_515), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g595 ( .A(n_515), .Y(n_595) );
INVx1_ASAP7_75t_L g720 ( .A(n_515), .Y(n_720) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_516), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_522), .Y(n_517) );
OR2x2_ASAP7_75t_L g691 ( .A(n_524), .B(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_SL g546 ( .A(n_526), .Y(n_546) );
OR2x2_ASAP7_75t_L g569 ( .A(n_526), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g580 ( .A(n_526), .B(n_556), .Y(n_580) );
AND2x2_ASAP7_75t_L g654 ( .A(n_526), .B(n_570), .Y(n_654) );
BUFx2_ASAP7_75t_L g737 ( .A(n_526), .Y(n_737) );
OR2x6_ASAP7_75t_L g526 ( .A(n_527), .B(n_534), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_542), .B(n_547), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
AND2x2_ASAP7_75t_L g689 ( .A(n_538), .B(n_611), .Y(n_689) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g548 ( .A(n_539), .B(n_541), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_540), .B(n_610), .Y(n_711) );
INVx1_ASAP7_75t_L g741 ( .A(n_540), .Y(n_741) );
NAND2x1p5_ASAP7_75t_L g637 ( .A(n_541), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_541), .B(n_677), .Y(n_714) );
INVxp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
AND2x4_ASAP7_75t_SL g578 ( .A(n_544), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_544), .B(n_572), .Y(n_725) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_545), .B(n_627), .Y(n_683) );
AND2x2_ASAP7_75t_L g701 ( .A(n_545), .B(n_654), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_546), .B(n_588), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_546), .A2(n_592), .B(n_634), .C(n_639), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_546), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_548), .A2(n_621), .B1(n_729), .B2(n_735), .C(n_739), .Y(n_728) );
INVx1_ASAP7_75t_SL g716 ( .A(n_549), .Y(n_716) );
OAI221xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_561), .B1(n_567), .B2(n_571), .C(n_788), .Y(n_550) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_553), .B(n_558), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g626 ( .A(n_555), .Y(n_626) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g600 ( .A(n_556), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g631 ( .A(n_556), .B(n_576), .Y(n_631) );
INVx2_ASAP7_75t_L g664 ( .A(n_556), .Y(n_664) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI32xp33_ASAP7_75t_L g715 ( .A1(n_559), .A2(n_606), .A3(n_637), .B1(n_716), .B2(n_717), .Y(n_715) );
OR2x2_ASAP7_75t_L g686 ( .A(n_560), .B(n_673), .Y(n_686) );
INVx1_ASAP7_75t_L g696 ( .A(n_561), .Y(n_696) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx2_ASAP7_75t_L g611 ( .A(n_562), .Y(n_611) );
AND2x2_ASAP7_75t_L g682 ( .A(n_562), .B(n_657), .Y(n_682) );
OR2x2_ASAP7_75t_L g713 ( .A(n_562), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_563), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g607 ( .A(n_566), .Y(n_607) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx2_ASAP7_75t_SL g572 ( .A(n_569), .Y(n_572) );
OR2x2_ASAP7_75t_L g659 ( .A(n_569), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_570), .B(n_588), .Y(n_587) );
NOR2xp67_ASAP7_75t_L g693 ( .A(n_570), .B(n_694), .Y(n_693) );
BUFx2_ASAP7_75t_L g706 ( .A(n_570), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B(n_578), .C(n_581), .Y(n_571) );
AND2x2_ASAP7_75t_L g721 ( .A(n_573), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g647 ( .A(n_577), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_577), .B(n_581), .Y(n_668) );
AND2x2_ASAP7_75t_L g699 ( .A(n_577), .B(n_700), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g709 ( .A1(n_579), .A2(n_710), .B(n_712), .C(n_715), .Y(n_709) );
AOI222xp33_ASAP7_75t_L g583 ( .A1(n_580), .A2(n_584), .B1(n_586), .B2(n_589), .C1(n_597), .C2(n_599), .Y(n_583) );
AND2x2_ASAP7_75t_L g651 ( .A(n_580), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g584 ( .A(n_581), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_SL g605 ( .A(n_581), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g582 ( .A(n_583), .B(n_602), .C(n_623), .D(n_633), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_585), .B(n_591), .Y(n_645) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g653 ( .A(n_588), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_SL g660 ( .A(n_588), .Y(n_660) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_590), .A2(n_624), .B(n_628), .C(n_632), .Y(n_623) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_591), .B(n_606), .Y(n_727) );
OR2x2_ASAP7_75t_L g731 ( .A(n_591), .B(n_617), .Y(n_731) );
INVx1_ASAP7_75t_L g704 ( .A(n_592), .Y(n_704) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_SL g638 ( .A(n_595), .Y(n_638) );
INVx1_ASAP7_75t_L g618 ( .A(n_596), .Y(n_618) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_598), .B(n_635), .Y(n_634) );
BUFx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g622 ( .A(n_600), .Y(n_622) );
AOI322xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_605), .A3(n_606), .B1(n_608), .B2(n_612), .C1(n_613), .C2(n_619), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_SL g684 ( .A1(n_605), .A2(n_685), .B(n_686), .C(n_687), .Y(n_684) );
INVx1_ASAP7_75t_L g707 ( .A(n_606), .Y(n_707) );
NOR2xp67_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g665 ( .A(n_611), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_617), .Y(n_687) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx3_ASAP7_75t_L g630 ( .A(n_627), .Y(n_630) );
OR2x2_ASAP7_75t_L g698 ( .A(n_627), .B(n_660), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_627), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_SL g730 ( .A(n_631), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_632), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND3xp33_ASAP7_75t_SL g735 ( .A(n_640), .B(n_736), .C(n_738), .Y(n_735) );
NOR3xp33_ASAP7_75t_SL g641 ( .A(n_642), .B(n_679), .C(n_708), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_643), .B(n_661), .Y(n_642) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B(n_649), .C(n_655), .Y(n_643) );
OAI31xp33_ASAP7_75t_L g688 ( .A1(n_644), .A2(n_666), .A3(n_689), .B(n_690), .Y(n_688) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx2_ASAP7_75t_L g703 ( .A(n_651), .Y(n_703) );
INVx1_ASAP7_75t_L g678 ( .A(n_653), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .B(n_659), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g705 ( .A(n_663), .B(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_L g744 ( .A(n_664), .Y(n_744) );
OAI22xp33_ASAP7_75t_SL g667 ( .A1(n_668), .A2(n_669), .B1(n_674), .B2(n_678), .Y(n_667) );
INVx3_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x4_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_673), .Y(n_685) );
OR2x2_ASAP7_75t_L g736 ( .A(n_673), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND3xp33_ASAP7_75t_SL g679 ( .A(n_680), .B(n_688), .C(n_695), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B(n_683), .C(n_684), .Y(n_680) );
INVx2_ASAP7_75t_L g717 ( .A(n_681), .Y(n_717) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_699), .B2(n_701), .C(n_702), .Y(n_695) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_705), .B2(n_707), .Y(n_702) );
NAND3xp33_ASAP7_75t_SL g708 ( .A(n_709), .B(n_718), .C(n_728), .Y(n_708) );
INVxp33_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B1(n_724), .B2(n_726), .Y(n_718) );
INVx2_ASAP7_75t_L g732 ( .A(n_719), .Y(n_732) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_729) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI22xp33_ASAP7_75t_SL g739 ( .A1(n_738), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
BUFx4f_ASAP7_75t_SL g755 ( .A(n_745), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
CKINVDCx11_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_748), .A2(n_753), .B(n_756), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVxp33_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx3_ASAP7_75t_SL g786 ( .A(n_777), .Y(n_786) );
AND2x2_ASAP7_75t_SL g777 ( .A(n_778), .B(n_779), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
INVx1_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
endmodule