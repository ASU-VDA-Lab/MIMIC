module fake_jpeg_16577_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_33),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_42),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_21),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_56),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_24),
.B1(n_28),
.B2(n_27),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_61),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_24),
.B1(n_28),
.B2(n_27),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_28),
.B1(n_24),
.B2(n_27),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_27),
.B1(n_29),
.B2(n_16),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_51),
.B1(n_54),
.B2(n_63),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_17),
.B1(n_29),
.B2(n_20),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_18),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_17),
.B1(n_29),
.B2(n_20),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_34),
.A2(n_23),
.B1(n_19),
.B2(n_15),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_36),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_31),
.B1(n_17),
.B2(n_20),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_59),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_31),
.B1(n_23),
.B2(n_19),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_67),
.A2(n_26),
.B1(n_49),
.B2(n_57),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_71),
.Y(n_92)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_81),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_43),
.B(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_25),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_54),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_103),
.B(n_104),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_64),
.C(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_61),
.B(n_19),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_59),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_74),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_109),
.B(n_87),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_26),
.B(n_52),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_118),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_65),
.B1(n_81),
.B2(n_66),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_116),
.B1(n_125),
.B2(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_65),
.B1(n_75),
.B2(n_70),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_129),
.B1(n_102),
.B2(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_72),
.B1(n_75),
.B2(n_45),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_131),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_18),
.B(n_46),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_132),
.B(n_101),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_68),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_124),
.B(n_126),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_77),
.B1(n_84),
.B2(n_80),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_80),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_128),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_18),
.B(n_44),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_130),
.B1(n_117),
.B2(n_113),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_142),
.B1(n_145),
.B2(n_136),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_104),
.B(n_101),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_138),
.B(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_141),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_106),
.C(n_105),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_147),
.C(n_145),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_117),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_105),
.B1(n_92),
.B2(n_91),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_22),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_92),
.B1(n_88),
.B2(n_57),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_109),
.B(n_78),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_149),
.A2(n_121),
.B1(n_122),
.B2(n_90),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_90),
.B(n_95),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_125),
.Y(n_158)
);

BUFx4f_ASAP7_75t_SL g151 ( 
.A(n_119),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_78),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_142),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_132),
.B(n_122),
.C(n_112),
.D(n_116),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_157),
.A2(n_158),
.B(n_165),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_57),
.B1(n_48),
.B2(n_76),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_163),
.A2(n_164),
.B1(n_139),
.B2(n_153),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_107),
.B1(n_30),
.B2(n_15),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_74),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_139),
.B1(n_135),
.B2(n_30),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_169),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_78),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_170),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_22),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_174),
.C(n_137),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_190),
.Y(n_192)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_144),
.C(n_133),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_184),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_133),
.C(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_191),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_150),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_188),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_154),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_189),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_135),
.C(n_22),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_30),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_166),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_196),
.Y(n_209)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_166),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_SL g198 ( 
.A1(n_188),
.A2(n_160),
.A3(n_163),
.B1(n_157),
.B2(n_170),
.C1(n_164),
.C2(n_158),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_191),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_170),
.B(n_173),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_199),
.B(n_204),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_189),
.Y(n_204)
);

XOR2x1_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_155),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_187),
.B1(n_190),
.B2(n_178),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_177),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_215),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_155),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_210),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_208),
.B(n_212),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_184),
.C(n_179),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_216),
.B(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_187),
.C(n_161),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_181),
.B1(n_0),
.B2(n_2),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_213),
.A2(n_203),
.B1(n_202),
.B2(n_195),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_8),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_8),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_200),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_9),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_217),
.A2(n_205),
.B(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_223),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_209),
.A2(n_214),
.B(n_194),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_224),
.A2(n_30),
.B1(n_4),
.B2(n_5),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_207),
.A2(n_192),
.B(n_1),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_9),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_212),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_228),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_210),
.B(n_1),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_12),
.B1(n_6),
.B2(n_7),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_10),
.B(n_5),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_218),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_231),
.A2(n_227),
.B(n_229),
.Y(n_234)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_12),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_241),
.B(n_6),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_8),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_0),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_218),
.B(n_221),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_245),
.B(n_242),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_10),
.C(n_13),
.Y(n_247)
);


endmodule