module fake_jpeg_12170_n_541 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_541);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_2),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_5),
.Y(n_112)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_60),
.B(n_65),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_78),
.Y(n_123)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_0),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_68),
.B(n_77),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_69),
.B(n_52),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_3),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

AND2x4_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_4),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_80),
.B(n_50),
.C(n_22),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_40),
.B(n_4),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_83),
.B(n_97),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_39),
.B(n_4),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_84),
.B(n_94),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_91),
.Y(n_108)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g143 ( 
.A(n_93),
.Y(n_143)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_47),
.B(n_5),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_19),
.B(n_5),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_57),
.A2(n_47),
.B1(n_42),
.B2(n_51),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_109),
.A2(n_125),
.B(n_141),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_112),
.B(n_118),
.C(n_39),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_54),
.A2(n_52),
.B1(n_45),
.B2(n_24),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_117),
.A2(n_139),
.B1(n_142),
.B2(n_36),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_46),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_70),
.A2(n_47),
.B1(n_51),
.B2(n_24),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_76),
.A2(n_44),
.B1(n_52),
.B2(n_24),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_127),
.A2(n_133),
.B1(n_38),
.B2(n_31),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_80),
.B(n_69),
.C(n_22),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_63),
.A2(n_44),
.B1(n_36),
.B2(n_38),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_67),
.A2(n_44),
.B1(n_31),
.B2(n_36),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_70),
.A2(n_34),
.B1(n_32),
.B2(n_38),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_75),
.A2(n_44),
.B1(n_31),
.B2(n_36),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_89),
.A2(n_100),
.B1(n_53),
.B2(n_32),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_144),
.A2(n_125),
.B(n_141),
.Y(n_222)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_93),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_148),
.B(n_162),
.Y(n_212)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_80),
.Y(n_185)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_93),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_171),
.B(n_202),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_106),
.A2(n_49),
.B1(n_48),
.B2(n_22),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_173),
.A2(n_222),
.B(n_117),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_174),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_41),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_175),
.B(n_192),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx4_ASAP7_75t_SL g284 ( 
.A(n_177),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_178),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g252 ( 
.A(n_180),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_181),
.A2(n_184),
.B1(n_209),
.B2(n_153),
.Y(n_273)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_183),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_130),
.A2(n_105),
.B1(n_102),
.B2(n_101),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_185),
.B(n_32),
.Y(n_265)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_186),
.Y(n_247)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_187),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_111),
.B(n_103),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_188),
.Y(n_267)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_190),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_191),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_41),
.Y(n_192)
);

BUFx6f_ASAP7_75t_SL g193 ( 
.A(n_108),
.Y(n_193)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_193),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_139),
.A2(n_86),
.B1(n_87),
.B2(n_98),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_194),
.A2(n_215),
.B1(n_135),
.B2(n_145),
.Y(n_248)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_41),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_196),
.B(n_200),
.Y(n_255)
);

AOI32xp33_ASAP7_75t_L g198 ( 
.A1(n_137),
.A2(n_150),
.A3(n_81),
.B1(n_88),
.B2(n_99),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_198),
.A2(n_227),
.B(n_9),
.C(n_10),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_126),
.Y(n_199)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_108),
.B(n_41),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_114),
.B(n_48),
.C(n_49),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_201),
.B(n_37),
.C(n_119),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_129),
.B(n_73),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_146),
.Y(n_203)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_204),
.Y(n_282)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_205),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_143),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_210),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_146),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_142),
.A2(n_90),
.B1(n_96),
.B2(n_46),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_134),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_143),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_218),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_140),
.A2(n_104),
.B1(n_38),
.B2(n_71),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_106),
.A2(n_33),
.B1(n_50),
.B2(n_85),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_216),
.A2(n_223),
.B1(n_154),
.B2(n_120),
.Y(n_245)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_132),
.B(n_138),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_220),
.Y(n_271)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_145),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_224),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_115),
.A2(n_50),
.B1(n_33),
.B2(n_32),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_113),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_228),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_109),
.A2(n_33),
.B(n_37),
.C(n_19),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_144),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_232),
.Y(n_250)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_116),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_115),
.B(n_81),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_231),
.B(n_6),
.Y(n_275)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_120),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_173),
.B(n_154),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_233),
.B(n_259),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_193),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_236),
.B(n_266),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g330 ( 
.A(n_238),
.B(n_270),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_185),
.A2(n_161),
.B(n_160),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_241),
.A2(n_190),
.B(n_177),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_248),
.A2(n_236),
.B1(n_260),
.B2(n_274),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_119),
.B1(n_128),
.B2(n_170),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_254),
.A2(n_283),
.B1(n_211),
.B2(n_178),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_128),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_264),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_265),
.B(n_270),
.C(n_260),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_188),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_212),
.B(n_32),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_268),
.B(n_277),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_185),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_279),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_214),
.A2(n_153),
.B1(n_7),
.B2(n_8),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_272),
.A2(n_276),
.B1(n_180),
.B2(n_174),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_188),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_275),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_227),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_201),
.B(n_197),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_202),
.B(n_9),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_215),
.A2(n_222),
.B1(n_179),
.B2(n_205),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_176),
.B(n_9),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_285),
.B(n_14),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_286),
.A2(n_14),
.B(n_239),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_288),
.B(n_300),
.Y(n_347)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_289),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_233),
.A2(n_179),
.B(n_225),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_290),
.A2(n_324),
.B(n_326),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_246),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_291),
.B(n_294),
.Y(n_338)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_293),
.A2(n_295),
.B1(n_332),
.B2(n_274),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_264),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_213),
.C(n_206),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_296),
.B(n_313),
.C(n_260),
.Y(n_348)
);

INVx11_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_297),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_251),
.A2(n_221),
.B1(n_220),
.B2(n_195),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_299),
.A2(n_302),
.B1(n_321),
.B2(n_252),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_251),
.A2(n_189),
.B1(n_204),
.B2(n_208),
.Y(n_302)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_306),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_307),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_264),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_308),
.B(n_311),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_SL g309 ( 
.A(n_267),
.B(n_230),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_309),
.B(n_333),
.Y(n_367)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_253),
.Y(n_310)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_310),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_259),
.B(n_187),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_240),
.A2(n_254),
.B1(n_248),
.B2(n_267),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_312),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_182),
.C(n_217),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_250),
.A2(n_219),
.B(n_199),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_314),
.A2(n_235),
.B(n_234),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_224),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_316),
.B(n_323),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_255),
.B(n_203),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_317),
.B(n_325),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_273),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_320),
.B1(n_252),
.B2(n_242),
.Y(n_340)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_253),
.Y(n_319)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_238),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_251),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_287),
.Y(n_322)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_322),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_266),
.B(n_11),
.Y(n_323)
);

AO22x1_ASAP7_75t_L g326 ( 
.A1(n_240),
.A2(n_14),
.B1(n_286),
.B2(n_241),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_287),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_327),
.A2(n_334),
.B1(n_335),
.B2(n_252),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_255),
.B(n_275),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_329),
.A2(n_330),
.B(n_265),
.Y(n_344)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_263),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_263),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_337),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_340),
.B(n_361),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_341),
.A2(n_342),
.B1(n_345),
.B2(n_350),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_290),
.A2(n_303),
.B1(n_315),
.B2(n_288),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_315),
.A2(n_237),
.B1(n_256),
.B2(n_235),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_343),
.A2(n_353),
.B1(n_362),
.B2(n_322),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_344),
.B(n_348),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_303),
.A2(n_256),
.B1(n_257),
.B2(n_237),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_297),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_346),
.B(n_351),
.Y(n_381)
);

XOR2x2_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_262),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_313),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_330),
.A2(n_257),
.B1(n_278),
.B2(n_249),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_301),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_352),
.A2(n_363),
.B(n_314),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_328),
.A2(n_234),
.B1(n_261),
.B2(n_280),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_295),
.A2(n_330),
.B1(n_320),
.B2(n_318),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_372),
.B1(n_302),
.B2(n_308),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_304),
.A2(n_262),
.B1(n_282),
.B2(n_244),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_328),
.A2(n_280),
.B1(n_261),
.B2(n_282),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_304),
.B(n_284),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_366),
.C(n_300),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_298),
.B(n_244),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_311),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_370),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_334),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_310),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_335),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_295),
.A2(n_247),
.B1(n_281),
.B2(n_293),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_291),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_378),
.B(n_384),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_379),
.B(n_393),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_380),
.A2(n_407),
.B(n_403),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_354),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_360),
.A2(n_326),
.B(n_309),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_385),
.A2(n_394),
.B(n_403),
.Y(n_422)
);

OAI32xp33_ASAP7_75t_L g386 ( 
.A1(n_374),
.A2(n_316),
.A3(n_326),
.B1(n_323),
.B2(n_296),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_386),
.B(n_387),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_345),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_389),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_390),
.A2(n_392),
.B1(n_400),
.B2(n_341),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_373),
.B(n_329),
.Y(n_391)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_391),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_369),
.A2(n_299),
.B1(n_321),
.B2(n_331),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_360),
.A2(n_324),
.B(n_331),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_396),
.A2(n_376),
.B1(n_372),
.B2(n_336),
.Y(n_421)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_355),
.Y(n_397)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_397),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_349),
.B(n_306),
.C(n_292),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_398),
.B(n_408),
.C(n_411),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_338),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_406),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_359),
.A2(n_305),
.B1(n_289),
.B2(n_327),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_319),
.Y(n_401)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_401),
.Y(n_419)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_347),
.A2(n_247),
.B(n_281),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_339),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_405),
.B(n_409),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_361),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_347),
.A2(n_356),
.B(n_352),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_344),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_371),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_410),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_370),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_367),
.B(n_348),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_407),
.A2(n_347),
.B(n_342),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_412),
.A2(n_438),
.B(n_422),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_364),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_416),
.B(n_435),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_393),
.B(n_350),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_417),
.B(n_420),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_418),
.A2(n_420),
.B1(n_441),
.B2(n_383),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_390),
.A2(n_356),
.B1(n_366),
.B2(n_354),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_421),
.A2(n_377),
.B1(n_429),
.B2(n_432),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_381),
.Y(n_424)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_424),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_358),
.C(n_365),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_431),
.C(n_381),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_382),
.A2(n_340),
.B1(n_357),
.B2(n_365),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_429),
.A2(n_395),
.B1(n_399),
.B2(n_382),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_406),
.A2(n_376),
.B1(n_336),
.B2(n_357),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_430),
.A2(n_440),
.B(n_410),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_408),
.C(n_398),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_384),
.A2(n_368),
.B1(n_375),
.B2(n_336),
.Y(n_433)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_433),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_379),
.B(n_368),
.Y(n_435)
);

NAND2x1p5_ASAP7_75t_L g438 ( 
.A(n_385),
.B(n_375),
.Y(n_438)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_439),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_387),
.A2(n_400),
.B1(n_395),
.B2(n_392),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_391),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_449),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_443),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_444),
.A2(n_458),
.B1(n_451),
.B2(n_466),
.Y(n_471)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_415),
.Y(n_445)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_445),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_425),
.C(n_426),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_401),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_416),
.B(n_386),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_441),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_452),
.B(n_461),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_440),
.A2(n_383),
.B(n_405),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_453),
.B(n_454),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_422),
.A2(n_380),
.B(n_394),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_434),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_456),
.B(n_419),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_426),
.B(n_389),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_457),
.B(n_436),
.Y(n_475)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_428),
.Y(n_458)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_458),
.Y(n_476)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_459),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_428),
.A2(n_388),
.B1(n_397),
.B2(n_402),
.Y(n_460)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_460),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_412),
.A2(n_438),
.B(n_423),
.Y(n_461)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_414),
.Y(n_463)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_463),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_464),
.B(n_417),
.Y(n_473)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_465),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_419),
.B(n_430),
.Y(n_466)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_466),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_444),
.A2(n_423),
.B1(n_431),
.B2(n_425),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_469),
.A2(n_471),
.B1(n_461),
.B2(n_462),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_485),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_464),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_479),
.Y(n_496)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_477),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_447),
.B(n_438),
.C(n_418),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_460),
.Y(n_486)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_486),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_470),
.A2(n_455),
.B1(n_445),
.B2(n_459),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_488),
.A2(n_484),
.B1(n_476),
.B2(n_478),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_487),
.A2(n_453),
.B(n_452),
.Y(n_490)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_490),
.Y(n_516)
);

MAJx2_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_494),
.C(n_502),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_448),
.C(n_442),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_495),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_482),
.B(n_446),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_467),
.B(n_448),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_499),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_467),
.B(n_449),
.C(n_457),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_501),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_479),
.Y(n_499)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_483),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_481),
.A2(n_454),
.B(n_443),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_471),
.B(n_475),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_504),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_472),
.B(n_450),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_493),
.B(n_474),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_508),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_468),
.C(n_480),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_494),
.B(n_474),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_481),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_492),
.B(n_468),
.C(n_480),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_512),
.A2(n_515),
.B(n_502),
.Y(n_519)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_500),
.Y(n_513)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_513),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_478),
.C(n_486),
.Y(n_515)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_517),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_519),
.A2(n_510),
.B(n_507),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_505),
.B(n_503),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_522),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_514),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_512),
.B(n_508),
.C(n_515),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_516),
.A2(n_490),
.B1(n_498),
.B2(n_473),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_524),
.B(n_496),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_504),
.C(n_499),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_526),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_530),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_529),
.A2(n_524),
.B(n_518),
.Y(n_533)
);

AOI21xp33_ASAP7_75t_L g536 ( 
.A1(n_533),
.A2(n_525),
.B(n_510),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_522),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_527),
.Y(n_535)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_535),
.B(n_536),
.C(n_532),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_526),
.C(n_523),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_521),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_539),
.A2(n_509),
.B1(n_511),
.B2(n_496),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_540),
.A2(n_491),
.B1(n_413),
.B2(n_437),
.Y(n_541)
);


endmodule