module fake_jpeg_26160_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_29),
.B1(n_22),
.B2(n_31),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_39),
.B1(n_24),
.B2(n_17),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_51),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_29),
.B1(n_22),
.B2(n_23),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_67),
.B1(n_77),
.B2(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_37),
.B1(n_39),
.B2(n_22),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_70),
.Y(n_98)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_80),
.B1(n_46),
.B2(n_44),
.Y(n_108)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_75),
.A2(n_46),
.B1(n_80),
.B2(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_22),
.B1(n_30),
.B2(n_27),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_39),
.B1(n_17),
.B2(n_33),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_33),
.B1(n_26),
.B2(n_16),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_81),
.B1(n_88),
.B2(n_91),
.Y(n_96)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_17),
.B1(n_33),
.B2(n_24),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_25),
.B(n_27),
.C(n_32),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_20),
.A3(n_21),
.B1(n_36),
.B2(n_34),
.Y(n_111)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_25),
.B1(n_32),
.B2(n_27),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_33),
.B1(n_24),
.B2(n_25),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_32),
.B1(n_16),
.B2(n_28),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_28),
.B1(n_26),
.B2(n_16),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_26),
.B1(n_28),
.B2(n_60),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_56),
.B(n_52),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_34),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_102),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_50),
.B1(n_57),
.B2(n_60),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_105),
.B1(n_116),
.B2(n_106),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_0),
.B(n_1),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_117),
.B1(n_90),
.B2(n_21),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_70),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_34),
.B(n_88),
.C(n_36),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_38),
.C(n_40),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_38),
.C(n_40),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_118),
.B1(n_89),
.B2(n_74),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_44),
.B1(n_41),
.B2(n_34),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_73),
.B1(n_85),
.B2(n_75),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_0),
.B(n_1),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_20),
.B1(n_19),
.B2(n_44),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_122),
.A2(n_119),
.B1(n_120),
.B2(n_100),
.Y(n_177)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_125),
.B(n_130),
.Y(n_171)
);

AOI22x1_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_68),
.B1(n_82),
.B2(n_78),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g166 ( 
.A1(n_128),
.A2(n_34),
.B(n_40),
.C(n_44),
.Y(n_166)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_65),
.B1(n_68),
.B2(n_81),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_136),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_65),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_131),
.B(n_144),
.Y(n_182)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_84),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_134),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_92),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_138),
.B(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_139),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_142),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_105),
.B1(n_93),
.B2(n_107),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_104),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_103),
.B(n_14),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_103),
.B(n_61),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_146),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_149),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_20),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_19),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_96),
.C(n_38),
.Y(n_157)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_161),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_181),
.B(n_184),
.Y(n_196)
);

OAI22x1_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_102),
.B1(n_117),
.B2(n_96),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g214 ( 
.A1(n_156),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_151),
.C(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_162),
.Y(n_213)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_163),
.A2(n_174),
.B1(n_125),
.B2(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_172),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_121),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_183),
.B(n_133),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_36),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_178),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_139),
.A2(n_120),
.B1(n_119),
.B2(n_100),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_141),
.B1(n_137),
.B2(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_126),
.A2(n_21),
.B(n_19),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_124),
.B(n_134),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_11),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_186),
.B(n_200),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_199),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_185),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_194),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_154),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_193),
.Y(n_230)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_202),
.B1(n_206),
.B2(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_212),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_129),
.C(n_119),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_62),
.B1(n_44),
.B2(n_41),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_42),
.C(n_21),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_211),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_180),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_190),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_164),
.A2(n_62),
.B1(n_21),
.B2(n_19),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_168),
.A2(n_0),
.B(n_1),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_181),
.B(n_208),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_153),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_209),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_176),
.B(n_9),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_161),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_214),
.A2(n_166),
.B(n_4),
.C(n_5),
.Y(n_236)
);

NOR2x1_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_156),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_221),
.A2(n_223),
.B1(n_228),
.B2(n_232),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_226),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_170),
.B1(n_183),
.B2(n_174),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_176),
.B(n_180),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_225),
.B(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_183),
.B1(n_157),
.B2(n_184),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_233),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_166),
.B1(n_177),
.B2(n_155),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_158),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_207),
.B(n_205),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_152),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_235),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_206),
.B1(n_193),
.B2(n_187),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_221),
.B(n_232),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_240),
.A2(n_241),
.B(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_224),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_189),
.C(n_199),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_244),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_203),
.C(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_224),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_247),
.A2(n_250),
.B1(n_236),
.B2(n_229),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_228),
.C(n_227),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_248),
.B(n_249),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_201),
.C(n_210),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_219),
.A2(n_196),
.B1(n_205),
.B2(n_211),
.Y(n_250)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_210),
.C(n_196),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_254),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_213),
.C(n_166),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_188),
.C(n_202),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_188),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_257),
.B(n_234),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_254),
.B(n_243),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_244),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_217),
.B1(n_226),
.B2(n_220),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_265),
.B1(n_272),
.B2(n_247),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_217),
.B1(n_220),
.B2(n_230),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_269),
.Y(n_284)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_255),
.A2(n_233),
.B1(n_236),
.B2(n_235),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_236),
.B1(n_249),
.B2(n_182),
.Y(n_280)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_245),
.B(n_250),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_276),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_248),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_279),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_264),
.A2(n_253),
.B(n_242),
.Y(n_278)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_260),
.B1(n_8),
.B2(n_11),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_10),
.C(n_14),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_283),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_268),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_9),
.C(n_13),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_286),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_10),
.B(n_13),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_287),
.A2(n_259),
.B1(n_273),
.B2(n_263),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_296),
.Y(n_299)
);

NOR2x1_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_272),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_297),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_286),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_277),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_300),
.B(n_303),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_298),
.A2(n_282),
.B(n_276),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_302),
.B(n_305),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_293),
.A2(n_274),
.B(n_283),
.Y(n_302)
);

NAND4xp25_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_285),
.C(n_281),
.D(n_11),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_279),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_8),
.C(n_12),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_291),
.B(n_12),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_310),
.B(n_303),
.C(n_8),
.Y(n_314)
);

NAND4xp25_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_293),
.C(n_294),
.D(n_292),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_295),
.B1(n_289),
.B2(n_288),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_311),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_309),
.B(n_299),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_314),
.C(n_307),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_312),
.A3(n_15),
.B1(n_6),
.B2(n_7),
.C1(n_5),
.C2(n_2),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_6),
.B(n_7),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_7),
.Y(n_318)
);


endmodule