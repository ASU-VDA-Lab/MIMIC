module fake_jpeg_4282_n_301 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_180;
wire n_51;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_2),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_38),
.B1(n_40),
.B2(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_36),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_28),
.B1(n_17),
.B2(n_22),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_48),
.B1(n_55),
.B2(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_15),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_28),
.B1(n_22),
.B2(n_21),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_54),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_28),
.B1(n_22),
.B2(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_47),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_22),
.B1(n_24),
.B2(n_21),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_63),
.B1(n_24),
.B2(n_17),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_17),
.B1(n_21),
.B2(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_37),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_76),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_32),
.B(n_23),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_69),
.B(n_71),
.C(n_16),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_39),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_R g71 ( 
.A(n_49),
.B(n_40),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_32),
.C(n_39),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_73),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_36),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_24),
.B1(n_38),
.B2(n_30),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_45),
.B1(n_38),
.B2(n_46),
.Y(n_101)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_30),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_15),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_53),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_100),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_55),
.B1(n_48),
.B2(n_42),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_81),
.B1(n_38),
.B2(n_65),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_82),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_20),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_99),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_33),
.B1(n_45),
.B2(n_38),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_75),
.B1(n_76),
.B2(n_44),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_18),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_20),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_54),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_25),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_111),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_72),
.C(n_64),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_129),
.C(n_107),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_66),
.B1(n_78),
.B2(n_72),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_115),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_101),
.B(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_73),
.Y(n_121)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_78),
.B1(n_76),
.B2(n_33),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_94),
.B1(n_102),
.B2(n_98),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_84),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_64),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_141),
.B1(n_144),
.B2(n_122),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_137),
.C(n_115),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_97),
.B(n_87),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_135),
.A2(n_148),
.B(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_87),
.C(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_87),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_145),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_94),
.B1(n_101),
.B2(n_91),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_111),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_143),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_105),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_109),
.B(n_105),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_154),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_98),
.B(n_106),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_98),
.B(n_92),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_112),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_152),
.B(n_156),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_106),
.B(n_88),
.Y(n_153)
);

FAx1_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_148),
.CI(n_144),
.CON(n_181),
.SN(n_181)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_109),
.B(n_96),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_110),
.Y(n_157)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_135),
.C(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_164),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_120),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_173),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_126),
.B(n_127),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_162),
.B(n_135),
.Y(n_192)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_122),
.B1(n_127),
.B2(n_125),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_181),
.B(n_163),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_168),
.A2(n_170),
.B1(n_179),
.B2(n_74),
.Y(n_206)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_171),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_117),
.B1(n_74),
.B2(n_57),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_120),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_155),
.B(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_119),
.Y(n_176)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_114),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_177),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_130),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_142),
.B1(n_152),
.B2(n_143),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_114),
.B1(n_67),
.B2(n_68),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_73),
.B1(n_63),
.B2(n_60),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_141),
.B1(n_151),
.B2(n_150),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_184),
.A2(n_186),
.B1(n_187),
.B2(n_205),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_150),
.B1(n_133),
.B2(n_134),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_133),
.B1(n_134),
.B2(n_149),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_149),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_190),
.C(n_193),
.Y(n_209)
);

AOI221xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_206),
.B1(n_19),
.B2(n_41),
.C(n_37),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_203),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_136),
.C(n_153),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_136),
.C(n_153),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_197),
.C(n_203),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_148),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_169),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_133),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_132),
.B(n_154),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_204),
.A2(n_166),
.B(n_171),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_142),
.B1(n_110),
.B2(n_104),
.Y(n_205)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_175),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_215),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_213),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_168),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_166),
.B(n_181),
.C(n_176),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_224),
.B1(n_191),
.B2(n_200),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_164),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_226),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_218),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_202),
.B(n_79),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_79),
.Y(n_219)
);

NOR2xp67_ASAP7_75t_SL g244 ( 
.A(n_219),
.B(n_221),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_159),
.C(n_179),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_223),
.C(n_227),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_159),
.C(n_165),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_80),
.B1(n_19),
.B2(n_26),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_185),
.B1(n_16),
.B2(n_25),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_193),
.C(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_80),
.B1(n_19),
.B2(n_26),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_52),
.C(n_62),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_187),
.C(n_186),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_242),
.C(n_246),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_243),
.B(n_16),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_184),
.B1(n_204),
.B2(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_192),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_37),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_80),
.B1(n_25),
.B2(n_26),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_238),
.B(n_225),
.Y(n_248)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_209),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_62),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_222),
.Y(n_243)
);

AOI21x1_ASAP7_75t_SL g245 ( 
.A1(n_221),
.A2(n_51),
.B(n_29),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_246),
.B(n_229),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_83),
.C(n_51),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_249),
.B(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_250),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_234),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_0),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_252),
.B(n_253),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_0),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_SL g267 ( 
.A(n_254),
.B(n_239),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_240),
.B(n_244),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_259),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_51),
.B1(n_83),
.B2(n_41),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_SL g275 ( 
.A1(n_257),
.A2(n_260),
.B(n_9),
.C(n_14),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_237),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_41),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_245),
.A2(n_0),
.B(n_1),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_228),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_266),
.B(n_267),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_228),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_242),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_271),
.B(n_272),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_239),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_41),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_274),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_1),
.Y(n_274)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_13),
.B(n_12),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_262),
.C(n_254),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_277),
.A2(n_278),
.B(n_280),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_262),
.C(n_253),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_265),
.C(n_263),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_37),
.B(n_29),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_284),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_29),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_282),
.A2(n_1),
.B(n_2),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_29),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_2),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_291),
.B(n_292),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_13),
.A3(n_12),
.B1(n_11),
.B2(n_10),
.C1(n_9),
.C2(n_7),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_283),
.A3(n_282),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_5),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_12),
.Y(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_3),
.B(n_4),
.C(n_6),
.D(n_8),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_297),
.B(n_293),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_8),
.C1(n_10),
.C2(n_286),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_296),
.C(n_4),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_3),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_299),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_8),
.Y(n_301)
);


endmodule