module real_jpeg_5038_n_20 (n_17, n_8, n_0, n_93, n_95, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_94, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_93;
input n_95;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_94;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_1),
.A2(n_18),
.B(n_85),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_1),
.B(n_18),
.C(n_33),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_2),
.B(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_5),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_6),
.A2(n_19),
.B(n_26),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_6),
.B(n_19),
.C(n_33),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_9),
.A2(n_13),
.B(n_31),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_11),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_11),
.B(n_16),
.C(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_12),
.A2(n_35),
.B(n_93),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g60 ( 
.A(n_12),
.B(n_61),
.C(n_95),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_13),
.B(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_14),
.A2(n_15),
.B(n_33),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_14),
.B(n_15),
.C(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_16),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_17),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

NAND3xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_29),
.C(n_31),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_40),
.B(n_41),
.Y(n_39)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_65),
.C(n_66),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_41),
.B(n_44),
.Y(n_45)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_87),
.B(n_89),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_42),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_44),
.Y(n_43)
);

NAND3xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_84),
.B(n_86),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_79),
.B(n_83),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B(n_77),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_69),
.B(n_73),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_68),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_63),
.B(n_67),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B(n_60),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_72),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_81),
.C(n_82),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_82),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_94),
.Y(n_59)
);


endmodule