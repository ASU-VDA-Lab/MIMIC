module fake_jpeg_4324_n_208 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_30),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_32),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_0),
.Y(n_46)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_14),
.B1(n_22),
.B2(n_27),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_41),
.B1(n_54),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_22),
.B1(n_27),
.B2(n_17),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_18),
.C(n_20),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_47),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_53),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_18),
.C(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_28),
.B(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_24),
.Y(n_53)
);

AO22x1_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_24),
.B1(n_21),
.B2(n_26),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_56),
.B1(n_65),
.B2(n_51),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_37),
.B1(n_30),
.B2(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_60),
.B(n_61),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_31),
.B1(n_16),
.B2(n_25),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_31),
.B1(n_29),
.B2(n_24),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_45),
.B(n_29),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_31),
.B1(n_35),
.B2(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_67),
.Y(n_88)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_73),
.Y(n_75)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_83),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_43),
.CI(n_47),
.CON(n_80),
.SN(n_80)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_80),
.B(n_85),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_90),
.B1(n_93),
.B2(n_79),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_91),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_59),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_69),
.B1(n_57),
.B2(n_61),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_87),
.B1(n_49),
.B2(n_42),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_50),
.B1(n_45),
.B2(n_48),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_56),
.B1(n_65),
.B2(n_68),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_32),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_50),
.B1(n_35),
.B2(n_34),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_62),
.C(n_71),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_106),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_82),
.B1(n_94),
.B2(n_89),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_111),
.Y(n_122)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_32),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_76),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_112),
.B(n_21),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_78),
.B(n_36),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_36),
.Y(n_112)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_84),
.Y(n_113)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_104),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_101),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_79),
.B1(n_81),
.B2(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_129),
.B1(n_112),
.B2(n_99),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_94),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_118),
.B(n_98),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_132),
.B1(n_35),
.B2(n_34),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_80),
.B(n_76),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_95),
.C(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_80),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_130),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_89),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_128),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_88),
.B(n_77),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_26),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_35),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_137),
.C(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_138),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_105),
.C(n_100),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_120),
.B1(n_116),
.B2(n_132),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_35),
.C(n_34),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_0),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_147),
.A2(n_116),
.B1(n_123),
.B2(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_148),
.B(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_0),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_149),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_149),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_155),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_159),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_118),
.B(n_125),
.C(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_118),
.B1(n_137),
.B2(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_136),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_142),
.B1(n_140),
.B2(n_135),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_158),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_118),
.B1(n_132),
.B2(n_126),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_145),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_144),
.C(n_124),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_163),
.C(n_161),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_134),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_173),
.Y(n_182)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_134),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_163),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_172),
.A2(n_174),
.B1(n_151),
.B2(n_160),
.Y(n_179)
);

OAI322xp33_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_118),
.A3(n_146),
.B1(n_130),
.B2(n_123),
.C1(n_115),
.C2(n_8),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_115),
.B(n_4),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_153),
.B(n_152),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_2),
.B(n_4),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_154),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_179),
.B1(n_170),
.B2(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_167),
.B(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_177),
.B(n_178),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_164),
.B(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_155),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_181),
.B(n_183),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_184),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_9),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_180),
.B1(n_172),
.B2(n_176),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_190),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_166),
.B1(n_165),
.B2(n_33),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_2),
.B(n_6),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_33),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_2),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_186),
.C(n_191),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_194),
.B(n_197),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_195),
.B(n_198),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_185),
.A2(n_7),
.B(n_9),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_196),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_9),
.B(n_10),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_189),
.B1(n_187),
.B2(n_197),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_33),
.C(n_12),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_10),
.A3(n_12),
.B1(n_13),
.B2(n_33),
.C1(n_199),
.C2(n_201),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_204),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_207),
.Y(n_208)
);


endmodule