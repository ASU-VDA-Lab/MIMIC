module fake_jpeg_28184_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx11_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_43),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_66),
.Y(n_74)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_62),
.Y(n_87)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_23),
.B1(n_31),
.B2(n_33),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_23),
.B1(n_45),
.B2(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_28),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_45),
.B1(n_41),
.B2(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_69),
.A2(n_53),
.B1(n_61),
.B2(n_60),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_70),
.A2(n_86),
.B1(n_104),
.B2(n_32),
.Y(n_121)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_71),
.B(n_77),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_76),
.Y(n_114)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_38),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_78),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_102),
.B1(n_53),
.B2(n_61),
.Y(n_113)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_49),
.B(n_21),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_100),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_53),
.A2(n_23),
.B1(n_44),
.B2(n_18),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_61),
.B1(n_51),
.B2(n_26),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_35),
.Y(n_96)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_28),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_105),
.Y(n_119)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_57),
.B(n_35),
.Y(n_100)
);

BUFx4f_ASAP7_75t_SL g101 ( 
.A(n_62),
.Y(n_101)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_49),
.A2(n_33),
.B1(n_19),
.B2(n_36),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_44),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_107),
.B(n_118),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_121),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_126),
.B1(n_99),
.B2(n_80),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_37),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_127),
.B(n_98),
.Y(n_141)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_49),
.B1(n_60),
.B2(n_19),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_37),
.Y(n_127)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_85),
.B1(n_91),
.B2(n_68),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_165),
.B1(n_109),
.B2(n_156),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_71),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_144),
.Y(n_185)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_155),
.B(n_16),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_87),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_147),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_129),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_149),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_69),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_95),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_145),
.B(n_146),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_84),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_39),
.C(n_101),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_154),
.C(n_161),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_79),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_151),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_108),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_36),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_157),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_118),
.A2(n_105),
.B(n_32),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_83),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_67),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_83),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_163),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_101),
.C(n_81),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_28),
.Y(n_162)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_82),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_26),
.B1(n_16),
.B2(n_29),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_166),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_147),
.A2(n_120),
.B1(n_115),
.B2(n_128),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_167),
.A2(n_184),
.B1(n_34),
.B2(n_22),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_106),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_180),
.B(n_183),
.Y(n_200)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_135),
.B1(n_124),
.B2(n_125),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_112),
.B1(n_106),
.B2(n_125),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_112),
.B1(n_122),
.B2(n_135),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_124),
.B(n_1),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_198),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_26),
.B1(n_16),
.B2(n_29),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_187),
.B(n_195),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_29),
.B(n_133),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_137),
.A2(n_148),
.B1(n_146),
.B2(n_151),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_193),
.B1(n_196),
.B2(n_139),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_145),
.A2(n_25),
.B1(n_24),
.B2(n_20),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_138),
.A2(n_0),
.B(n_1),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_25),
.B1(n_24),
.B2(n_20),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_138),
.Y(n_201)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_154),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_220),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_150),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_209),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_165),
.Y(n_210)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_214),
.Y(n_235)
);

NOR2x1_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_153),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_169),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_140),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_217),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_164),
.Y(n_219)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_180),
.B(n_11),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_140),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_223),
.C(n_224),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_46),
.C(n_40),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_46),
.C(n_40),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_20),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_226),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_167),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_170),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_172),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_172),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_20),
.Y(n_229)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_192),
.B1(n_179),
.B2(n_166),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_210),
.B1(n_200),
.B2(n_222),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_192),
.B(n_183),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_238),
.A2(n_0),
.B(n_1),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_252),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_179),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_228),
.A2(n_178),
.B1(n_195),
.B2(n_174),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_251),
.A2(n_254),
.B1(n_216),
.B2(n_191),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_187),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_202),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_256),
.A2(n_251),
.B1(n_249),
.B2(n_243),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_231),
.A2(n_212),
.B1(n_213),
.B2(n_201),
.Y(n_257)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_257),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_221),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_259),
.B(n_274),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_260),
.A2(n_263),
.B1(n_238),
.B2(n_234),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_184),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_270),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_208),
.B1(n_213),
.B2(n_220),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_205),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_267),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_203),
.C(n_223),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_269),
.C(n_273),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_224),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_230),
.A2(n_191),
.B(n_10),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_268),
.A2(n_252),
.B(n_231),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_46),
.C(n_40),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_34),
.C(n_22),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_275),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_270),
.B(n_237),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_281),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_264),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_284),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_285),
.B(n_2),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_263),
.A2(n_247),
.B1(n_236),
.B2(n_253),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_271),
.B1(n_243),
.B2(n_253),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_267),
.C(n_259),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_278),
.C(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_292),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_240),
.B1(n_234),
.B2(n_249),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_291),
.A2(n_34),
.B1(n_25),
.B2(n_24),
.Y(n_308)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_254),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_297),
.A2(n_304),
.B1(n_287),
.B2(n_25),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_250),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_302),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_301),
.C(n_278),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_255),
.C(n_245),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_280),
.B(n_246),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_272),
.B1(n_274),
.B2(n_232),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_303),
.A2(n_306),
.B1(n_279),
.B2(n_283),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_258),
.B1(n_254),
.B2(n_34),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_295),
.B(n_296),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_9),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_308),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_304),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_309),
.B(n_294),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_298),
.A2(n_288),
.B1(n_279),
.B2(n_285),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_315),
.Y(n_326)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_312),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_313),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_296),
.A2(n_24),
.B1(n_8),
.B2(n_4),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_7),
.C(n_12),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_307),
.C(n_297),
.Y(n_320)
);

XOR2x2_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_7),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_318),
.A2(n_8),
.B(n_14),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_7),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_320),
.B(n_322),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_324),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_323),
.A2(n_314),
.B(n_313),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_309),
.C(n_317),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_328),
.B(n_330),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_310),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_329),
.Y(n_333)
);

OAI21x1_ASAP7_75t_SL g335 ( 
.A1(n_333),
.A2(n_325),
.B(n_324),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_322),
.A3(n_334),
.B1(n_327),
.B2(n_6),
.C1(n_8),
.C2(n_9),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_4),
.B(n_9),
.C(n_12),
.Y(n_337)
);

O2A1O1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_4),
.B(n_12),
.C(n_2),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_338),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_339),
.B(n_3),
.Y(n_340)
);

NAND3xp33_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_3),
.C(n_318),
.Y(n_341)
);


endmodule