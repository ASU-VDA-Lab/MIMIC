module fake_jpeg_31525_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_15),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_0),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_56),
.Y(n_58)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_45),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_40),
.B1(n_4),
.B2(n_5),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_64),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_65),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_5),
.B(n_6),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_4),
.Y(n_79)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_47),
.C(n_37),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_13),
.C(n_16),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_43),
.B1(n_22),
.B2(n_23),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_83),
.Y(n_85)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_8),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_43),
.B1(n_24),
.B2(n_26),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_43),
.B1(n_21),
.B2(n_27),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_36),
.B1(n_17),
.B2(n_9),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_7),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_96),
.B1(n_30),
.B2(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_12),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_91),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_34),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_72),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_78),
.C(n_76),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_98),
.C(n_95),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_33),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_85),
.B1(n_86),
.B2(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_106),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_105),
.B(n_107),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_90),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_108),
.C(n_100),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_103),
.B(n_97),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);


endmodule