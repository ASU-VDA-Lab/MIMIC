module real_jpeg_5355_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_0),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_0),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_0),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_0),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_0),
.B(n_134),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_0),
.B(n_181),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_0),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_0),
.B(n_309),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_1),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_1),
.Y(n_186)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_1),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_1),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_1),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_2),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_3),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_3),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_3),
.B(n_186),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_3),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_3),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_3),
.B(n_387),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_3),
.B(n_143),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_4),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_4),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_4),
.B(n_53),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_4),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_4),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_4),
.B(n_212),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_5),
.Y(n_102)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_5),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_5),
.Y(n_145)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_6),
.Y(n_537)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_7),
.Y(n_188)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_7),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_7),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_8),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_8),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_8),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_8),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_8),
.B(n_59),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_8),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_8),
.B(n_373),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_8),
.B(n_418),
.Y(n_417)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_10),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_10),
.B(n_45),
.Y(n_168)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_10),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_10),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_10),
.B(n_325),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_10),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_10),
.B(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_11),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_11),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_11),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_12),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_12),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_12),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_12),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_12),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_12),
.B(n_202),
.Y(n_201)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_14),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_15),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_15),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_15),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_15),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_15),
.B(n_212),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_15),
.B(n_390),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_15),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_16),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_16),
.B(n_190),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_16),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_16),
.B(n_68),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_16),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_16),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_16),
.B(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_16),
.B(n_358),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_17),
.B(n_28),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_17),
.B(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_17),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_17),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_17),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_17),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_17),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_18),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_18),
.B(n_66),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_18),
.B(n_197),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_18),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_18),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_18),
.B(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_18),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_18),
.B(n_409),
.Y(n_408)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_535),
.B(n_538),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_41),
.B(n_77),
.C(n_534),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_24),
.B(n_48),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.C(n_35),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_26),
.A2(n_30),
.B1(n_40),
.B2(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_52),
.C(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_33),
.Y(n_192)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_34),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_34),
.Y(n_199)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_34),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_35),
.B(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_47),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_73),
.C(n_75),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_49),
.B(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_62),
.C(n_63),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_50),
.B(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_52),
.A2(n_57),
.B1(n_69),
.B2(n_108),
.Y(n_112)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_53),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_54),
.Y(n_356)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_55),
.Y(n_136)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_55),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_55),
.Y(n_391)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_55),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_64),
.C(n_69),
.Y(n_63)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_63),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_64),
.A2(n_65),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_69),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_69),
.A2(n_103),
.B1(n_104),
.B2(n_108),
.Y(n_504)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_72),
.Y(n_213)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_72),
.Y(n_336)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_72),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_119),
.B(n_533),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_116),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_79),
.B(n_116),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_113),
.C(n_114),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_80),
.A2(n_81),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_97),
.C(n_109),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_82),
.A2(n_83),
.B1(n_508),
.B2(n_510),
.Y(n_507)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_86),
.C(n_88),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.C(n_95),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_89),
.B(n_498),
.Y(n_497)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_498)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_97),
.A2(n_109),
.B1(n_110),
.B2(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_97),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.C(n_108),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_98),
.B(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_100),
.Y(n_262)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_103),
.A2(n_104),
.B1(n_201),
.B2(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_104),
.B(n_196),
.C(n_201),
.Y(n_505)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_107),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_107),
.Y(n_287)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_113),
.B(n_114),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_527),
.B(n_532),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_491),
.B(n_524),
.Y(n_120)
);

OAI21x1_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_292),
.B(n_490),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_241),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_123),
.B(n_241),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_193),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_124),
.B(n_194),
.C(n_223),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_166),
.C(n_175),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_125),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_140),
.C(n_155),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_126),
.B(n_476),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_132),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_133),
.C(n_137),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_131),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_131),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_134),
.Y(n_219)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_140),
.A2(n_141),
.B1(n_155),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.C(n_151),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_142),
.B(n_151),
.Y(n_466)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_145),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_146),
.B(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_155),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_156),
.B(n_158),
.C(n_163),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g376 ( 
.A(n_160),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_161),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_162),
.B(n_201),
.C(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_162),
.A2(n_163),
.B1(n_201),
.B2(n_204),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_166),
.B(n_175),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_174),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_167)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_172),
.C(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_169),
.A2(n_173),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_171),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_173),
.B(n_228),
.C(n_234),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_174),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_187),
.C(n_189),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_176),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_184),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_177),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_180),
.B(n_184),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_186),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_187),
.B(n_189),
.Y(n_270)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_192),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_223),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_205),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_195),
.B(n_206),
.C(n_222),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_203),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_214),
.B1(n_221),
.B2(n_222),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.C(n_211),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_211),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_215),
.B(n_217),
.C(n_220),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_235),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_225),
.B(n_227),
.C(n_235),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_229),
.B(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_239),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_248),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_243),
.B(n_246),
.Y(n_486)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_248),
.B(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_268),
.C(n_271),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_250),
.B(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_259),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_251),
.A2(n_252),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_254),
.A2(n_255),
.B(n_258),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_254),
.B(n_259),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.C(n_265),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_434)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_265),
.B(n_434),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_266),
.B(n_369),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_271),
.Y(n_480)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_283),
.C(n_288),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_273),
.B(n_468),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.C(n_280),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_274),
.B(n_446),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_276),
.A2(n_280),
.B1(n_281),
.B2(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_276),
.Y(n_447)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_283),
.B(n_288),
.Y(n_468)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_484),
.B(n_489),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_471),
.B(n_483),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_453),
.B(n_470),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_427),
.B(n_452),
.Y(n_295)
);

AOI21x1_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_395),
.B(n_426),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_361),
.B(n_394),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_338),
.B(n_360),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_316),
.B(n_337),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_313),
.B(n_315),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_311),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_311),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_308),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_308),
.Y(n_317)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_307),
.Y(n_323)
);

INVx3_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_318),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_326),
.B2(n_327),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_319),
.B(n_329),
.C(n_333),
.Y(n_359)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_324),
.Y(n_349)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_325),
.Y(n_348)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_333),
.B2(n_334),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_332),
.Y(n_370)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_359),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_359),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_350),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_349),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_349),
.C(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_346),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_342),
.B(n_346),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_350),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_351),
.B(n_380),
.C(n_381),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_357),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_357),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_364),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_378),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_365),
.B(n_379),
.C(n_382),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_368),
.C(n_371),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_374),
.B1(n_375),
.B2(n_377),
.Y(n_371)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_372),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_377),
.Y(n_404)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_382),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_385),
.Y(n_382)
);

MAJx2_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_389),
.C(n_392),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_389),
.B1(n_392),
.B2(n_393),
.Y(n_385)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_386),
.Y(n_392)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_389),
.Y(n_393)
);

INVx6_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_425),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_425),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_406),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_405),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_398),
.B(n_405),
.C(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_404),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_403),
.Y(n_399)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_400),
.Y(n_441)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_403),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_404),
.B(n_441),
.C(n_442),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_406),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_414),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_416),
.C(n_423),
.Y(n_430)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_407),
.Y(n_541)
);

FAx1_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_410),
.CI(n_411),
.CON(n_407),
.SN(n_407)
);

MAJx2_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_410),
.C(n_411),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_416),
.B1(n_423),
.B2(n_424),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_422),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_422),
.Y(n_437)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_424),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_450),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_450),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_439),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_431),
.C(n_439),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_435),
.B2(n_436),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_462),
.C(n_463),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_443),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_444),
.C(n_449),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_448),
.B2(n_449),
.Y(n_443)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_444),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_445),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_469),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_469),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_460),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_459),
.C(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_457),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_464),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_465),
.C(n_467),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_467),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_481),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_481),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_473),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_478),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_475),
.B(n_478),
.C(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_487),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_487),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_519),
.Y(n_491)
);

OAI21xp33_ASAP7_75t_L g524 ( 
.A1(n_492),
.A2(n_525),
.B(n_526),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_493),
.B(n_512),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_493),
.B(n_512),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_495),
.B1(n_501),
.B2(n_511),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_494),
.B(n_502),
.C(n_507),
.Y(n_531)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_497),
.C(n_499),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_496),
.B(n_515),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_497),
.A2(n_499),
.B1(n_500),
.B2(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_497),
.Y(n_516)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_501),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_507),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_505),
.C(n_506),
.Y(n_502)
);

FAx1_ASAP7_75t_SL g517 ( 
.A(n_503),
.B(n_505),
.CI(n_506),
.CON(n_517),
.SN(n_517)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_508),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_517),
.C(n_518),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_513),
.A2(n_514),
.B1(n_517),
.B2(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_517),
.Y(n_522)
);

BUFx24_ASAP7_75t_SL g542 ( 
.A(n_517),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_518),
.B(n_521),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_520),
.B(n_523),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_523),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_528),
.B(n_531),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_531),
.Y(n_532)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

BUFx12f_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_536),
.Y(n_539)
);

INVx13_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_540),
.Y(n_538)
);


endmodule