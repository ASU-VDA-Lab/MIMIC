module fake_jpeg_8353_n_32 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_32);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_32;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_15;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_7),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_13),
.B(n_2),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_8),
.Y(n_17)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_0),
.B(n_1),
.Y(n_18)
);

FAx1_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_17),
.CI(n_14),
.CON(n_26),
.SN(n_26)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_4),
.C(n_5),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_29),
.C(n_30),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_25),
.Y(n_30)
);

AO21x1_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_26),
.B(n_24),
.Y(n_32)
);


endmodule