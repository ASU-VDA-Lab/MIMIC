module fake_aes_7726_n_1362 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1362);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1362;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_298;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVxp33_ASAP7_75t_L g295 ( .A(n_115), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_95), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_253), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_250), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_6), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_150), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_280), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_58), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_252), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_13), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_175), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_181), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_66), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_208), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_195), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_36), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_248), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_56), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_139), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_271), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_138), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_94), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_98), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_171), .Y(n_318) );
INVxp33_ASAP7_75t_SL g319 ( .A(n_75), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_10), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_44), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_156), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_178), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_52), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_272), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_254), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_154), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_12), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_246), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_230), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_19), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_256), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_123), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_213), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_127), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_71), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_41), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_129), .Y(n_338) );
CKINVDCx16_ASAP7_75t_R g339 ( .A(n_206), .Y(n_339) );
INVxp33_ASAP7_75t_L g340 ( .A(n_126), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_93), .Y(n_341) );
INVxp67_ASAP7_75t_L g342 ( .A(n_134), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_64), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_293), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_87), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_7), .Y(n_346) );
INVxp67_ASAP7_75t_SL g347 ( .A(n_78), .Y(n_347) );
INVxp33_ASAP7_75t_SL g348 ( .A(n_199), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_80), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_113), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_135), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_3), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_165), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_99), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_270), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_67), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_14), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_279), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_15), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_119), .Y(n_360) );
INVxp33_ASAP7_75t_L g361 ( .A(n_240), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_184), .Y(n_362) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_64), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_108), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_192), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_236), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_288), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_200), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_18), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_191), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_216), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_32), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_83), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_116), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_1), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_7), .Y(n_376) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_84), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_223), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_131), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_88), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_71), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_100), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_106), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_51), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_258), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_247), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_261), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_58), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_109), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_70), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_267), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_25), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_57), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_215), .Y(n_394) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_130), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_260), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_237), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_76), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_282), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_11), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_269), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_251), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_46), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_76), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_235), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_292), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_8), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_56), .Y(n_408) );
BUFx3_ASAP7_75t_L g409 ( .A(n_193), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_110), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_2), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_174), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_245), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_274), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_65), .Y(n_415) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_186), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_4), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_225), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_204), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_196), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_161), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_72), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_275), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_222), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_3), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_153), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_2), .Y(n_427) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_74), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_103), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_50), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_60), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_234), .Y(n_432) );
INVxp33_ASAP7_75t_L g433 ( .A(n_198), .Y(n_433) );
CKINVDCx16_ASAP7_75t_R g434 ( .A(n_80), .Y(n_434) );
INVxp67_ASAP7_75t_L g435 ( .A(n_36), .Y(n_435) );
INVxp33_ASAP7_75t_L g436 ( .A(n_16), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_231), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_128), .B(n_217), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_101), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_243), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_327), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_362), .B(n_0), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_362), .B(n_0), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_327), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_327), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_428), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_300), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_414), .B(n_1), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_327), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_327), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_364), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_297), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_436), .B(n_4), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_364), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_297), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_364), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_322), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_322), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_364), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_295), .B(n_5), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_326), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_324), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_302), .B(n_5), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_364), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_396), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_389), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_340), .B(n_6), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_326), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_428), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_361), .B(n_8), .Y(n_470) );
INVx5_ASAP7_75t_L g471 ( .A(n_389), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_330), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_330), .Y(n_473) );
INVx3_ASAP7_75t_L g474 ( .A(n_428), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_471), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_462), .B(n_339), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_462), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_461), .B(n_433), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_460), .B(n_429), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_463), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_471), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_452), .B(n_455), .Y(n_482) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_444), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_465), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_465), .Y(n_485) );
BUFx4f_ASAP7_75t_L g486 ( .A(n_463), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_463), .Y(n_487) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_444), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_452), .A2(n_328), .B1(n_331), .B2(n_321), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_463), .B(n_302), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_452), .B(n_308), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_461), .B(n_301), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_463), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_453), .A2(n_319), .B1(n_434), .B2(n_325), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_463), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_453), .A2(n_328), .B1(n_331), .B2(n_321), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_468), .B(n_342), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_455), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_455), .Y(n_499) );
NOR2x1p5_ASAP7_75t_L g500 ( .A(n_442), .B(n_299), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_471), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_457), .B(n_320), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_457), .B(n_308), .Y(n_503) );
INVx4_ASAP7_75t_L g504 ( .A(n_465), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_453), .A2(n_384), .B1(n_427), .B2(n_336), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_471), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_457), .B(n_318), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_460), .A2(n_319), .B1(n_325), .B2(n_300), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_458), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_471), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_444), .Y(n_511) );
INVx4_ASAP7_75t_L g512 ( .A(n_465), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_444), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_458), .B(n_296), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_473), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_473), .Y(n_517) );
BUFx4_ASAP7_75t_L g518 ( .A(n_442), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_473), .B(n_320), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_498), .Y(n_520) );
INVx4_ASAP7_75t_L g521 ( .A(n_486), .Y(n_521) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_486), .Y(n_522) );
BUFx12f_ASAP7_75t_L g523 ( .A(n_476), .Y(n_523) );
BUFx3_ASAP7_75t_L g524 ( .A(n_484), .Y(n_524) );
INVx5_ASAP7_75t_L g525 ( .A(n_504), .Y(n_525) );
INVx5_ASAP7_75t_L g526 ( .A(n_504), .Y(n_526) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_500), .B(n_448), .Y(n_527) );
BUFx4f_ASAP7_75t_L g528 ( .A(n_476), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_502), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_477), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_477), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_478), .B(n_460), .Y(n_532) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_486), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_502), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_498), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_476), .B(n_447), .Y(n_536) );
INVx2_ASAP7_75t_SL g537 ( .A(n_500), .Y(n_537) );
BUFx8_ASAP7_75t_L g538 ( .A(n_518), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_486), .A2(n_447), .B1(n_412), .B2(n_351), .Y(n_539) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_484), .Y(n_540) );
AND2x6_ASAP7_75t_SL g541 ( .A(n_479), .B(n_448), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_479), .A2(n_470), .B1(n_443), .B2(n_467), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_479), .B(n_470), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_496), .A2(n_470), .B1(n_443), .B2(n_467), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_502), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_502), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_499), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_502), .Y(n_548) );
BUFx3_ASAP7_75t_L g549 ( .A(n_484), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_509), .B(n_468), .Y(n_550) );
INVx2_ASAP7_75t_SL g551 ( .A(n_518), .Y(n_551) );
BUFx3_ASAP7_75t_L g552 ( .A(n_485), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_509), .B(n_472), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_519), .Y(n_554) );
INVx4_ASAP7_75t_L g555 ( .A(n_490), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_515), .B(n_472), .Y(n_556) );
OR2x2_ASAP7_75t_SL g557 ( .A(n_508), .B(n_373), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_509), .B(n_296), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_499), .B(n_438), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_490), .B(n_336), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_505), .A2(n_412), .B1(n_351), .B2(n_299), .Y(n_561) );
INVx4_ASAP7_75t_L g562 ( .A(n_490), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_519), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_490), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_508), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_519), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_492), .B(n_323), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_497), .B(n_323), .Y(n_568) );
O2A1O1Ixp5_ASAP7_75t_L g569 ( .A1(n_482), .A2(n_487), .B(n_493), .C(n_480), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_519), .Y(n_570) );
INVx3_ASAP7_75t_L g571 ( .A(n_490), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_494), .A2(n_346), .B1(n_356), .B2(n_310), .Y(n_572) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_513), .Y(n_573) );
OAI21xp33_ASAP7_75t_L g574 ( .A1(n_480), .A2(n_348), .B(n_384), .Y(n_574) );
O2A1O1Ixp5_ASAP7_75t_L g575 ( .A1(n_487), .A2(n_395), .B(n_416), .C(n_371), .Y(n_575) );
INVx4_ASAP7_75t_L g576 ( .A(n_504), .Y(n_576) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_485), .Y(n_577) );
BUFx8_ASAP7_75t_L g578 ( .A(n_493), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_513), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_494), .B(n_375), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_516), .Y(n_582) );
NAND2x1p5_ASAP7_75t_L g583 ( .A(n_495), .B(n_427), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_495), .A2(n_431), .B1(n_430), .B2(n_307), .Y(n_584) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_516), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_489), .Y(n_586) );
AND2x4_ASAP7_75t_L g587 ( .A(n_489), .B(n_430), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_517), .B(n_348), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_491), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_517), .B(n_438), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_485), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_504), .B(n_298), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_512), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_512), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_512), .B(n_365), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_491), .B(n_431), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_503), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_503), .Y(n_598) );
INVxp67_ASAP7_75t_L g599 ( .A(n_507), .Y(n_599) );
OR2x6_ASAP7_75t_L g600 ( .A(n_507), .B(n_393), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_512), .A2(n_304), .B1(n_343), .B2(n_312), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_475), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_475), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_475), .B(n_347), .Y(n_604) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_530), .Y(n_605) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_578), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_560), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_599), .A2(n_373), .B1(n_346), .B2(n_356), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_528), .B(n_310), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_589), .B(n_369), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_560), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_578), .Y(n_612) );
INVx3_ASAP7_75t_SL g613 ( .A(n_551), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_531), .A2(n_369), .B1(n_398), .B2(n_392), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_562), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_536), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_578), .A2(n_377), .B1(n_363), .B2(n_392), .Y(n_617) );
AOI222xp33_ASAP7_75t_L g618 ( .A1(n_528), .A2(n_435), .B1(n_398), .B2(n_404), .C1(n_359), .C2(n_357), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_586), .A2(n_334), .B1(n_355), .B2(n_329), .Y(n_619) );
BUFx2_ASAP7_75t_L g620 ( .A(n_538), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_597), .B(n_329), .Y(n_621) );
O2A1O1Ixp5_ASAP7_75t_L g622 ( .A1(n_575), .A2(n_332), .B(n_341), .C(n_318), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_600), .Y(n_623) );
OA21x2_ASAP7_75t_L g624 ( .A1(n_569), .A2(n_335), .B(n_333), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_537), .B(n_349), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_520), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_520), .Y(n_627) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_600), .Y(n_628) );
INVx3_ASAP7_75t_L g629 ( .A(n_562), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_538), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_562), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_535), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_555), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_598), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_543), .B(n_334), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_586), .A2(n_352), .B1(n_376), .B2(n_372), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_557), .B(n_388), .Y(n_637) );
BUFx8_ASAP7_75t_L g638 ( .A(n_523), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_555), .Y(n_639) );
BUFx8_ASAP7_75t_L g640 ( .A(n_523), .Y(n_640) );
BUFx3_ASAP7_75t_L g641 ( .A(n_525), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_596), .B(n_355), .Y(n_642) );
CKINVDCx16_ASAP7_75t_R g643 ( .A(n_539), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_587), .A2(n_400), .B1(n_403), .B2(n_390), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_600), .B(n_407), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_538), .Y(n_646) );
NOR2xp67_ASAP7_75t_SL g647 ( .A(n_522), .B(n_378), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_587), .A2(n_571), .B1(n_564), .B2(n_529), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_535), .Y(n_649) );
OAI22x1_ASAP7_75t_L g650 ( .A1(n_561), .A2(n_378), .B1(n_413), .B2(n_391), .Y(n_650) );
INVx2_ASAP7_75t_SL g651 ( .A(n_596), .Y(n_651) );
INVx2_ASAP7_75t_SL g652 ( .A(n_596), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_583), .Y(n_653) );
BUFx2_ASAP7_75t_L g654 ( .A(n_541), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_588), .B(n_391), .Y(n_655) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_540), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_588), .B(n_532), .Y(n_657) );
BUFx4f_ASAP7_75t_L g658 ( .A(n_587), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_542), .B(n_413), .Y(n_659) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_540), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_564), .Y(n_661) );
BUFx8_ASAP7_75t_SL g662 ( .A(n_565), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_544), .B(n_421), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_583), .B(n_421), .Y(n_664) );
INVx2_ASAP7_75t_SL g665 ( .A(n_527), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_571), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_547), .A2(n_411), .B(n_415), .C(n_408), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_581), .B(n_417), .Y(n_668) );
AOI21xp33_ASAP7_75t_L g669 ( .A1(n_521), .A2(n_424), .B(n_426), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_559), .B(n_424), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_521), .B(n_422), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_547), .Y(n_672) );
NAND3x1_ASAP7_75t_L g673 ( .A(n_565), .B(n_425), .C(n_335), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_572), .A2(n_338), .B1(n_432), .B2(n_333), .Y(n_674) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_521), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_L g676 ( .A1(n_580), .A2(n_381), .B(n_337), .C(n_338), .Y(n_676) );
BUFx3_ASAP7_75t_L g677 ( .A(n_525), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_534), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_545), .B(n_337), .Y(n_679) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_540), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_546), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_548), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_604), .B(n_381), .Y(n_683) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_540), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_576), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_554), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_550), .A2(n_553), .B(n_573), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_563), .A2(n_428), .B1(n_439), .B2(n_432), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_604), .Y(n_689) );
AND2x6_ASAP7_75t_L g690 ( .A(n_522), .B(n_439), .Y(n_690) );
INVx4_ASAP7_75t_L g691 ( .A(n_522), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_566), .Y(n_692) );
BUFx2_ASAP7_75t_L g693 ( .A(n_522), .Y(n_693) );
AND2x6_ASAP7_75t_L g694 ( .A(n_533), .B(n_396), .Y(n_694) );
BUFx2_ASAP7_75t_L g695 ( .A(n_533), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_604), .B(n_428), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_570), .Y(n_697) );
INVx2_ASAP7_75t_SL g698 ( .A(n_579), .Y(n_698) );
INVx5_ASAP7_75t_L g699 ( .A(n_533), .Y(n_699) );
A2O1A1Ixp33_ASAP7_75t_L g700 ( .A1(n_580), .A2(n_305), .B(n_306), .C(n_303), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_585), .A2(n_501), .B(n_481), .Y(n_701) );
INVx1_ASAP7_75t_SL g702 ( .A(n_558), .Y(n_702) );
OAI22xp5_ASAP7_75t_SL g703 ( .A1(n_584), .A2(n_311), .B1(n_313), .B2(n_309), .Y(n_703) );
NAND2xp33_ASAP7_75t_L g704 ( .A(n_533), .B(n_481), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_582), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_582), .Y(n_706) );
OR2x6_ASAP7_75t_L g707 ( .A(n_576), .B(n_314), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_592), .A2(n_501), .B(n_481), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_559), .B(n_315), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_602), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g711 ( .A1(n_556), .A2(n_317), .B(n_344), .C(n_316), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_602), .Y(n_712) );
O2A1O1Ixp33_ASAP7_75t_L g713 ( .A1(n_590), .A2(n_350), .B(n_353), .C(n_345), .Y(n_713) );
INVx2_ASAP7_75t_SL g714 ( .A(n_590), .Y(n_714) );
NAND2x1p5_ASAP7_75t_L g715 ( .A(n_576), .B(n_401), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_584), .B(n_9), .Y(n_716) );
INVx2_ASAP7_75t_SL g717 ( .A(n_525), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_525), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_593), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_556), .B(n_354), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_593), .Y(n_721) );
CKINVDCx11_ASAP7_75t_R g722 ( .A(n_577), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_574), .B(n_358), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_603), .Y(n_724) );
BUFx3_ASAP7_75t_L g725 ( .A(n_526), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_601), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_634), .B(n_601), .Y(n_727) );
OAI21x1_ASAP7_75t_L g728 ( .A1(n_715), .A2(n_591), .B(n_594), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_726), .A2(n_595), .B1(n_568), .B2(n_567), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_616), .B(n_595), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_658), .A2(n_549), .B1(n_552), .B2(n_524), .Y(n_731) );
OAI211xp5_ASAP7_75t_L g732 ( .A1(n_617), .A2(n_592), .B(n_366), .C(n_367), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_658), .A2(n_594), .B1(n_549), .B2(n_552), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_605), .B(n_526), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_605), .Y(n_735) );
BUFx2_ASAP7_75t_SL g736 ( .A(n_606), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_623), .B(n_526), .Y(n_737) );
INVx3_ASAP7_75t_L g738 ( .A(n_641), .Y(n_738) );
OAI21x1_ASAP7_75t_L g739 ( .A1(n_715), .A2(n_591), .B(n_341), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_683), .Y(n_740) );
NAND2x1p5_ASAP7_75t_L g741 ( .A(n_607), .B(n_611), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_679), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_679), .Y(n_743) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_617), .A2(n_360), .B1(n_370), .B2(n_368), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_716), .Y(n_745) );
INVx3_ASAP7_75t_SL g746 ( .A(n_630), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_657), .A2(n_524), .B1(n_526), .B2(n_577), .Y(n_747) );
OAI221xp5_ASAP7_75t_L g748 ( .A1(n_636), .A2(n_420), .B1(n_374), .B2(n_379), .C(n_380), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_608), .A2(n_577), .B1(n_382), .B2(n_385), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_623), .B(n_577), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_628), .B(n_9), .Y(n_751) );
INVx3_ASAP7_75t_L g752 ( .A(n_641), .Y(n_752) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_646), .Y(n_753) );
OAI221xp5_ASAP7_75t_L g754 ( .A1(n_636), .A2(n_440), .B1(n_383), .B2(n_437), .C(n_387), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_626), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_651), .A2(n_406), .B1(n_410), .B2(n_394), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_653), .B(n_418), .Y(n_757) );
OAI221xp5_ASAP7_75t_L g758 ( .A1(n_637), .A2(n_419), .B1(n_423), .B2(n_386), .C(n_397), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_668), .A2(n_332), .B1(n_386), .B2(n_402), .C(n_397), .Y(n_759) );
OR2x6_ASAP7_75t_L g760 ( .A(n_606), .B(n_399), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_653), .B(n_10), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_652), .A2(n_409), .B1(n_401), .B2(n_402), .Y(n_762) );
INVx6_ASAP7_75t_L g763 ( .A(n_699), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_707), .A2(n_399), .B1(n_409), .B2(n_446), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_714), .B(n_11), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_707), .A2(n_469), .B1(n_474), .B2(n_446), .Y(n_766) );
AOI21xp33_ASAP7_75t_L g767 ( .A1(n_702), .A2(n_405), .B(n_389), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_626), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_703), .A2(n_469), .B1(n_474), .B2(n_446), .Y(n_769) );
AND2x4_ASAP7_75t_L g770 ( .A(n_612), .B(n_12), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_628), .B(n_13), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_612), .B(n_14), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_648), .A2(n_469), .B1(n_474), .B2(n_446), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g774 ( .A1(n_643), .A2(n_405), .B1(n_389), .B2(n_446), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_707), .A2(n_474), .B1(n_469), .B2(n_445), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_648), .B(n_15), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_689), .A2(n_474), .B1(n_469), .B2(n_405), .Y(n_777) );
AOI22xp33_ASAP7_75t_SL g778 ( .A1(n_654), .A2(n_405), .B1(n_389), .B2(n_471), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_627), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_610), .B(n_16), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_644), .A2(n_405), .B1(n_445), .B2(n_441), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_644), .B(n_17), .Y(n_782) );
BUFx2_ASAP7_75t_L g783 ( .A(n_638), .Y(n_783) );
OAI21x1_ASAP7_75t_L g784 ( .A1(n_627), .A2(n_445), .B(n_441), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_671), .Y(n_785) );
BUFx2_ASAP7_75t_R g786 ( .A(n_620), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_649), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_649), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_672), .Y(n_789) );
INVx1_ASAP7_75t_SL g790 ( .A(n_722), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_671), .Y(n_791) );
OR2x2_ASAP7_75t_L g792 ( .A(n_614), .B(n_17), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_705), .A2(n_445), .B1(n_449), .B2(n_441), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_672), .Y(n_794) );
AND2x4_ASAP7_75t_L g795 ( .A(n_665), .B(n_18), .Y(n_795) );
BUFx3_ASAP7_75t_L g796 ( .A(n_638), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_706), .A2(n_449), .B1(n_450), .B2(n_441), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_642), .A2(n_449), .B1(n_451), .B2(n_450), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_719), .Y(n_799) );
INVxp67_ASAP7_75t_L g800 ( .A(n_675), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_645), .A2(n_449), .B1(n_451), .B2(n_450), .Y(n_801) );
INVx2_ASAP7_75t_SL g802 ( .A(n_640), .Y(n_802) );
AOI222xp33_ASAP7_75t_L g803 ( .A1(n_650), .A2(n_450), .B1(n_451), .B2(n_454), .C1(n_456), .C2(n_459), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_696), .Y(n_804) );
BUFx3_ASAP7_75t_L g805 ( .A(n_722), .Y(n_805) );
AOI221xp5_ASAP7_75t_L g806 ( .A1(n_667), .A2(n_454), .B1(n_451), .B2(n_456), .C(n_466), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_687), .A2(n_466), .B1(n_454), .B2(n_456), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_678), .Y(n_808) );
AND2x4_ASAP7_75t_L g809 ( .A(n_615), .B(n_19), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_681), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_619), .A2(n_501), .B1(n_506), .B2(n_510), .Y(n_811) );
AO22x1_ASAP7_75t_SL g812 ( .A1(n_613), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_663), .A2(n_456), .B1(n_454), .B2(n_459), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_632), .A2(n_459), .B1(n_466), .B2(n_471), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_682), .A2(n_459), .B1(n_466), .B2(n_464), .Y(n_815) );
NAND2xp5_ASAP7_75t_SL g816 ( .A(n_656), .B(n_506), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_686), .A2(n_697), .B1(n_692), .B2(n_635), .Y(n_817) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_675), .Y(n_818) );
INVx3_ASAP7_75t_L g819 ( .A(n_677), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_719), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_664), .A2(n_471), .B1(n_506), .B2(n_510), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_639), .Y(n_822) );
BUFx3_ASAP7_75t_L g823 ( .A(n_677), .Y(n_823) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_656), .Y(n_824) );
OAI21x1_ASAP7_75t_L g825 ( .A1(n_708), .A2(n_510), .B(n_464), .Y(n_825) );
OR2x2_ASAP7_75t_L g826 ( .A(n_609), .B(n_20), .Y(n_826) );
AND2x4_ASAP7_75t_L g827 ( .A(n_615), .B(n_21), .Y(n_827) );
AND2x4_ASAP7_75t_L g828 ( .A(n_629), .B(n_22), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_709), .A2(n_464), .B1(n_444), .B2(n_471), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_659), .A2(n_464), .B1(n_444), .B2(n_488), .Y(n_830) );
OR2x6_ASAP7_75t_L g831 ( .A(n_640), .B(n_23), .Y(n_831) );
CKINVDCx6p67_ASAP7_75t_R g832 ( .A(n_613), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_721), .Y(n_833) );
BUFx2_ASAP7_75t_SL g834 ( .A(n_690), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_724), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_621), .A2(n_444), .B1(n_464), .B2(n_25), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_721), .Y(n_837) );
INVx6_ASAP7_75t_L g838 ( .A(n_699), .Y(n_838) );
INVx1_ASAP7_75t_SL g839 ( .A(n_690), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_661), .Y(n_840) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_690), .A2(n_694), .B1(n_673), .B2(n_625), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g842 ( .A1(n_674), .A2(n_23), .B1(n_24), .B2(n_26), .Y(n_842) );
AND2x4_ASAP7_75t_L g843 ( .A(n_629), .B(n_24), .Y(n_843) );
CKINVDCx9p33_ASAP7_75t_R g844 ( .A(n_693), .Y(n_844) );
OAI22xp33_ASAP7_75t_SL g845 ( .A1(n_670), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_845) );
CKINVDCx16_ASAP7_75t_R g846 ( .A(n_690), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_710), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_666), .Y(n_848) );
INVx1_ASAP7_75t_SL g849 ( .A(n_690), .Y(n_849) );
OAI22xp33_ASAP7_75t_L g850 ( .A1(n_720), .A2(n_27), .B1(n_28), .B2(n_29), .Y(n_850) );
CKINVDCx11_ASAP7_75t_R g851 ( .A(n_725), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_698), .A2(n_444), .B1(n_464), .B2(n_31), .Y(n_852) );
OAI221xp5_ASAP7_75t_L g853 ( .A1(n_618), .A2(n_464), .B1(n_30), .B2(n_31), .C(n_32), .Y(n_853) );
OAI22xp5_ASAP7_75t_SL g854 ( .A1(n_662), .A2(n_29), .B1(n_30), .B2(n_33), .Y(n_854) );
INVx4_ASAP7_75t_L g855 ( .A(n_699), .Y(n_855) );
AND2x4_ASAP7_75t_L g856 ( .A(n_725), .B(n_33), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_655), .A2(n_464), .B1(n_511), .B2(n_488), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_625), .B(n_667), .Y(n_858) );
INVx2_ASAP7_75t_SL g859 ( .A(n_699), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_832), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_858), .A2(n_662), .B1(n_669), .B2(n_633), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_735), .Y(n_862) );
INVx3_ASAP7_75t_SL g863 ( .A(n_796), .Y(n_863) );
BUFx2_ASAP7_75t_L g864 ( .A(n_831), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_835), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_744), .A2(n_633), .B1(n_631), .B2(n_694), .Y(n_866) );
INVx3_ASAP7_75t_L g867 ( .A(n_855), .Y(n_867) );
AOI22xp33_ASAP7_75t_SL g868 ( .A1(n_770), .A2(n_694), .B1(n_624), .B2(n_685), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_730), .B(n_700), .Y(n_869) );
AOI222xp33_ASAP7_75t_L g870 ( .A1(n_854), .A2(n_711), .B1(n_700), .B2(n_676), .C1(n_723), .C2(n_688), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_785), .A2(n_694), .B1(n_695), .B2(n_685), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_846), .A2(n_710), .B1(n_712), .B2(n_691), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_770), .B(n_711), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_772), .B(n_676), .Y(n_874) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_791), .A2(n_688), .B1(n_713), .B2(n_712), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_808), .Y(n_876) );
BUFx2_ASAP7_75t_L g877 ( .A(n_831), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_853), .A2(n_694), .B1(n_624), .B2(n_691), .Y(n_878) );
OR2x2_ASAP7_75t_SL g879 ( .A(n_792), .B(n_624), .Y(n_879) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_818), .Y(n_880) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_758), .A2(n_622), .B1(n_701), .B2(n_647), .C(n_717), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_810), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_745), .A2(n_718), .B1(n_704), .B2(n_684), .Y(n_883) );
OAI221xp5_ASAP7_75t_L g884 ( .A1(n_748), .A2(n_622), .B1(n_680), .B2(n_660), .C(n_656), .Y(n_884) );
AOI221xp5_ASAP7_75t_L g885 ( .A1(n_740), .A2(n_684), .B1(n_680), .B2(n_660), .C(n_656), .Y(n_885) );
BUFx4f_ASAP7_75t_L g886 ( .A(n_831), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_847), .Y(n_887) );
AOI22xp33_ASAP7_75t_SL g888 ( .A1(n_772), .A2(n_684), .B1(n_680), .B2(n_660), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_760), .A2(n_684), .B1(n_680), .B2(n_660), .Y(n_889) );
NAND3xp33_ASAP7_75t_L g890 ( .A(n_778), .B(n_488), .C(n_483), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_771), .A2(n_514), .B1(n_511), .B2(n_488), .Y(n_891) );
INVxp67_ASAP7_75t_L g892 ( .A(n_818), .Y(n_892) );
AOI22xp33_ASAP7_75t_SL g893 ( .A1(n_795), .A2(n_34), .B1(n_35), .B2(n_37), .Y(n_893) );
OAI221xp5_ASAP7_75t_L g894 ( .A1(n_754), .A2(n_514), .B1(n_511), .B2(n_488), .C(n_483), .Y(n_894) );
INVx4_ASAP7_75t_L g895 ( .A(n_783), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_795), .Y(n_896) );
CKINVDCx5p33_ASAP7_75t_R g897 ( .A(n_753), .Y(n_897) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_816), .A2(n_488), .B(n_483), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_856), .A2(n_34), .B1(n_35), .B2(n_37), .Y(n_899) );
OR2x2_ASAP7_75t_L g900 ( .A(n_826), .B(n_38), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_760), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_901) );
OAI221xp5_ASAP7_75t_L g902 ( .A1(n_729), .A2(n_817), .B1(n_841), .B2(n_780), .C(n_759), .Y(n_902) );
AND2x4_ASAP7_75t_L g903 ( .A(n_855), .B(n_39), .Y(n_903) );
OAI221xp5_ASAP7_75t_L g904 ( .A1(n_729), .A2(n_514), .B1(n_511), .B2(n_488), .C(n_483), .Y(n_904) );
OR2x6_ASAP7_75t_L g905 ( .A(n_834), .B(n_40), .Y(n_905) );
OAI221xp5_ASAP7_75t_L g906 ( .A1(n_817), .A2(n_514), .B1(n_511), .B2(n_483), .C(n_44), .Y(n_906) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_856), .A2(n_41), .B1(n_42), .B2(n_43), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_727), .B(n_42), .Y(n_908) );
AOI221xp5_ASAP7_75t_L g909 ( .A1(n_842), .A2(n_514), .B1(n_511), .B2(n_483), .C(n_47), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_809), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_842), .A2(n_514), .B1(n_511), .B2(n_483), .Y(n_911) );
AOI31xp33_ASAP7_75t_L g912 ( .A1(n_841), .A2(n_43), .A3(n_45), .B(n_46), .Y(n_912) );
OA21x2_ASAP7_75t_L g913 ( .A1(n_825), .A2(n_514), .B(n_90), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_771), .A2(n_45), .B1(n_47), .B2(n_48), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_780), .B(n_48), .Y(n_915) );
OAI211xp5_ASAP7_75t_L g916 ( .A1(n_774), .A2(n_49), .B(n_50), .C(n_51), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_809), .A2(n_49), .B1(n_52), .B2(n_53), .Y(n_917) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_800), .Y(n_918) );
AOI21xp5_ASAP7_75t_L g919 ( .A1(n_816), .A2(n_91), .B(n_89), .Y(n_919) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_805), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_920) );
AOI21xp33_ASAP7_75t_L g921 ( .A1(n_803), .A2(n_54), .B(n_55), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_760), .A2(n_57), .B1(n_59), .B2(n_60), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_827), .A2(n_59), .B1(n_61), .B2(n_62), .Y(n_923) );
AOI21xp5_ASAP7_75t_L g924 ( .A1(n_807), .A2(n_96), .B(n_92), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g925 ( .A(n_746), .Y(n_925) );
OAI211xp5_ASAP7_75t_L g926 ( .A1(n_774), .A2(n_732), .B(n_749), .C(n_769), .Y(n_926) );
OR2x2_ASAP7_75t_L g927 ( .A(n_751), .B(n_61), .Y(n_927) );
BUFx2_ASAP7_75t_L g928 ( .A(n_805), .Y(n_928) );
INVx4_ASAP7_75t_L g929 ( .A(n_851), .Y(n_929) );
HB1xp67_ASAP7_75t_L g930 ( .A(n_800), .Y(n_930) );
AOI221xp5_ASAP7_75t_L g931 ( .A1(n_850), .A2(n_62), .B1(n_63), .B2(n_65), .C(n_66), .Y(n_931) );
AOI322xp5_ASAP7_75t_L g932 ( .A1(n_850), .A2(n_63), .A3(n_67), .B1(n_68), .B2(n_69), .C1(n_70), .C2(n_72), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_827), .A2(n_843), .B1(n_828), .B2(n_782), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_756), .A2(n_68), .B1(n_69), .B2(n_73), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_828), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_843), .A2(n_77), .B1(n_78), .B2(n_79), .Y(n_936) );
OR2x2_ASAP7_75t_L g937 ( .A(n_741), .B(n_77), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_776), .A2(n_79), .B1(n_81), .B2(n_82), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_822), .Y(n_939) );
INVx8_ASAP7_75t_L g940 ( .A(n_734), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_742), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_941) );
OAI221xp5_ASAP7_75t_L g942 ( .A1(n_756), .A2(n_84), .B1(n_85), .B2(n_86), .C(n_97), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_743), .A2(n_85), .B1(n_86), .B2(n_102), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_799), .Y(n_944) );
INVx2_ASAP7_75t_L g945 ( .A(n_820), .Y(n_945) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_755), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_736), .A2(n_104), .B1(n_105), .B2(n_107), .Y(n_947) );
OAI211xp5_ASAP7_75t_SL g948 ( .A1(n_757), .A2(n_111), .B(n_112), .C(n_114), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_762), .A2(n_117), .B1(n_118), .B2(n_120), .Y(n_949) );
INVx4_ASAP7_75t_L g950 ( .A(n_851), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_833), .Y(n_951) );
OA21x2_ASAP7_75t_L g952 ( .A1(n_784), .A2(n_121), .B(n_122), .Y(n_952) );
OR2x2_ASAP7_75t_L g953 ( .A(n_741), .B(n_124), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_769), .A2(n_125), .B1(n_132), .B2(n_133), .Y(n_954) );
AO31x2_ASAP7_75t_L g955 ( .A1(n_836), .A2(n_136), .A3(n_137), .B(n_140), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_840), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_790), .B(n_141), .Y(n_957) );
OAI211xp5_ASAP7_75t_SL g958 ( .A1(n_801), .A2(n_142), .B(n_143), .C(n_144), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_804), .A2(n_145), .B1(n_146), .B2(n_147), .Y(n_959) );
AOI221xp5_ASAP7_75t_L g960 ( .A1(n_845), .A2(n_148), .B1(n_149), .B2(n_151), .C(n_152), .Y(n_960) );
AOI22xp33_ASAP7_75t_SL g961 ( .A1(n_839), .A2(n_155), .B1(n_157), .B2(n_158), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_761), .A2(n_159), .B1(n_160), .B2(n_162), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_737), .B(n_163), .Y(n_963) );
OR2x2_ASAP7_75t_L g964 ( .A(n_746), .B(n_164), .Y(n_964) );
AOI22xp33_ASAP7_75t_SL g965 ( .A1(n_849), .A2(n_166), .B1(n_167), .B2(n_168), .Y(n_965) );
INVxp67_ASAP7_75t_L g966 ( .A(n_768), .Y(n_966) );
OA21x2_ASAP7_75t_L g967 ( .A1(n_767), .A2(n_169), .B(n_170), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_848), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_750), .A2(n_172), .B1(n_173), .B2(n_176), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_802), .B(n_177), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_779), .B(n_294), .Y(n_971) );
BUFx12f_ASAP7_75t_L g972 ( .A(n_786), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_765), .Y(n_973) );
AOI21xp5_ASAP7_75t_L g974 ( .A1(n_857), .A2(n_179), .B(n_180), .Y(n_974) );
INVx3_ASAP7_75t_L g975 ( .A(n_763), .Y(n_975) );
OAI221xp5_ASAP7_75t_L g976 ( .A1(n_801), .A2(n_182), .B1(n_183), .B2(n_185), .C(n_187), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_787), .Y(n_977) );
A2O1A1Ixp33_ASAP7_75t_L g978 ( .A1(n_806), .A2(n_188), .B(n_189), .C(n_190), .Y(n_978) );
AOI31xp33_ASAP7_75t_L g979 ( .A1(n_778), .A2(n_194), .A3(n_197), .B(n_201), .Y(n_979) );
OAI22xp33_ASAP7_75t_L g980 ( .A1(n_764), .A2(n_202), .B1(n_203), .B2(n_205), .Y(n_980) );
OAI22xp33_ASAP7_75t_L g981 ( .A1(n_788), .A2(n_207), .B1(n_209), .B2(n_210), .Y(n_981) );
CKINVDCx5p33_ASAP7_75t_R g982 ( .A(n_844), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_837), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_977), .B(n_789), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_946), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_946), .B(n_794), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_886), .A2(n_823), .B1(n_762), .B2(n_821), .Y(n_987) );
NAND2xp5_ASAP7_75t_SL g988 ( .A(n_886), .B(n_859), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_966), .B(n_823), .Y(n_989) );
INVx2_ASAP7_75t_L g990 ( .A(n_887), .Y(n_990) );
AOI21x1_ASAP7_75t_L g991 ( .A1(n_913), .A2(n_739), .B(n_852), .Y(n_991) );
OAI21xp5_ASAP7_75t_L g992 ( .A1(n_902), .A2(n_781), .B(n_830), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_869), .B(n_738), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_966), .B(n_738), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_944), .Y(n_995) );
OAI221xp5_ASAP7_75t_SL g996 ( .A1(n_932), .A2(n_781), .B1(n_773), .B2(n_812), .C(n_813), .Y(n_996) );
INVx2_ASAP7_75t_L g997 ( .A(n_945), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_870), .A2(n_752), .B1(n_819), .B2(n_775), .Y(n_998) );
OAI33xp33_ASAP7_75t_L g999 ( .A1(n_901), .A2(n_798), .A3(n_766), .B1(n_814), .B2(n_731), .B3(n_844), .Y(n_999) );
INVx2_ASAP7_75t_L g1000 ( .A(n_951), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_873), .A2(n_752), .B1(n_819), .B2(n_773), .Y(n_1001) );
NAND3xp33_ASAP7_75t_L g1002 ( .A(n_960), .B(n_830), .C(n_857), .Y(n_1002) );
INVx2_ASAP7_75t_L g1003 ( .A(n_983), .Y(n_1003) );
AO21x2_ASAP7_75t_L g1004 ( .A1(n_884), .A2(n_728), .B(n_811), .Y(n_1004) );
INVx4_ASAP7_75t_R g1005 ( .A(n_910), .Y(n_1005) );
OAI33xp33_ASAP7_75t_L g1006 ( .A1(n_922), .A2(n_813), .A3(n_793), .B1(n_797), .B2(n_829), .B3(n_815), .Y(n_1006) );
OAI211xp5_ASAP7_75t_SL g1007 ( .A1(n_861), .A2(n_793), .B(n_797), .C(n_829), .Y(n_1007) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_933), .A2(n_747), .B1(n_733), .B2(n_777), .C(n_815), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_874), .B(n_838), .Y(n_1009) );
OAI22xp33_ASAP7_75t_L g1010 ( .A1(n_912), .A2(n_905), .B1(n_877), .B2(n_864), .Y(n_1010) );
NAND2xp5_ASAP7_75t_SL g1011 ( .A(n_888), .B(n_824), .Y(n_1011) );
AO221x1_ASAP7_75t_L g1012 ( .A1(n_872), .A2(n_824), .B1(n_838), .B2(n_763), .C(n_777), .Y(n_1012) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_880), .B(n_824), .Y(n_1013) );
AOI221xp5_ASAP7_75t_L g1014 ( .A1(n_931), .A2(n_747), .B1(n_733), .B2(n_824), .C(n_838), .Y(n_1014) );
AO21x2_ASAP7_75t_L g1015 ( .A1(n_904), .A2(n_763), .B(n_212), .Y(n_1015) );
AOI33xp33_ASAP7_75t_L g1016 ( .A1(n_893), .A2(n_211), .A3(n_214), .B1(n_218), .B2(n_219), .B3(n_220), .Y(n_1016) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_899), .A2(n_221), .B1(n_224), .B2(n_226), .C(n_227), .Y(n_1017) );
BUFx2_ASAP7_75t_L g1018 ( .A(n_905), .Y(n_1018) );
AOI33xp33_ASAP7_75t_L g1019 ( .A1(n_893), .A2(n_228), .A3(n_229), .B1(n_232), .B2(n_233), .B3(n_238), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_865), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_876), .B(n_239), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_882), .B(n_241), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_862), .B(n_291), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_956), .B(n_242), .Y(n_1024) );
INVx2_ASAP7_75t_L g1025 ( .A(n_913), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_952), .Y(n_1026) );
OAI33xp33_ASAP7_75t_L g1027 ( .A1(n_934), .A2(n_244), .A3(n_249), .B1(n_255), .B2(n_257), .B3(n_259), .Y(n_1027) );
INVx2_ASAP7_75t_L g1028 ( .A(n_952), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_968), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_939), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_880), .B(n_262), .Y(n_1031) );
OAI211xp5_ASAP7_75t_L g1032 ( .A1(n_899), .A2(n_263), .B(n_264), .C(n_265), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_918), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_879), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_905), .A2(n_266), .B1(n_268), .B2(n_273), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_888), .A2(n_276), .B1(n_277), .B2(n_278), .Y(n_1036) );
OAI221xp5_ASAP7_75t_L g1037 ( .A1(n_907), .A2(n_281), .B1(n_283), .B2(n_284), .C(n_285), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_921), .A2(n_286), .B1(n_287), .B2(n_289), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_911), .A2(n_290), .B1(n_907), .B2(n_900), .Y(n_1039) );
NAND3xp33_ASAP7_75t_L g1040 ( .A(n_920), .B(n_938), .C(n_935), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_918), .B(n_930), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_909), .A2(n_915), .B1(n_973), .B2(n_911), .Y(n_1042) );
NOR2xp33_ASAP7_75t_SL g1043 ( .A(n_972), .B(n_860), .Y(n_1043) );
NAND3xp33_ASAP7_75t_L g1044 ( .A(n_868), .B(n_916), .C(n_920), .Y(n_1044) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_982), .A2(n_903), .B1(n_929), .B2(n_950), .Y(n_1045) );
BUFx3_ASAP7_75t_L g1046 ( .A(n_863), .Y(n_1046) );
INVxp67_ASAP7_75t_SL g1047 ( .A(n_930), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_896), .B(n_892), .Y(n_1048) );
INVx2_ASAP7_75t_L g1049 ( .A(n_955), .Y(n_1049) );
CKINVDCx20_ASAP7_75t_R g1050 ( .A(n_863), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_908), .Y(n_1051) );
INVx2_ASAP7_75t_L g1052 ( .A(n_955), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_928), .A2(n_895), .B1(n_940), .B2(n_942), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_892), .B(n_927), .Y(n_1054) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_940), .B(n_937), .Y(n_1055) );
BUFx3_ASAP7_75t_L g1056 ( .A(n_940), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_895), .A2(n_903), .B1(n_914), .B2(n_866), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_955), .Y(n_1058) );
AOI221xp5_ASAP7_75t_L g1059 ( .A1(n_917), .A2(n_936), .B1(n_923), .B2(n_875), .C(n_941), .Y(n_1059) );
OR2x6_ASAP7_75t_L g1060 ( .A(n_889), .B(n_953), .Y(n_1060) );
OAI22xp33_ASAP7_75t_L g1061 ( .A1(n_979), .A2(n_929), .B1(n_950), .B2(n_964), .Y(n_1061) );
INVxp67_ASAP7_75t_SL g1062 ( .A(n_872), .Y(n_1062) );
OAI211xp5_ASAP7_75t_L g1063 ( .A1(n_868), .A2(n_943), .B(n_926), .C(n_957), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_955), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_975), .B(n_867), .Y(n_1065) );
INVx2_ASAP7_75t_L g1066 ( .A(n_967), .Y(n_1066) );
OA21x2_ASAP7_75t_L g1067 ( .A1(n_878), .A2(n_885), .B(n_890), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_867), .B(n_975), .Y(n_1068) );
OAI221xp5_ASAP7_75t_L g1069 ( .A1(n_878), .A2(n_906), .B1(n_891), .B2(n_881), .C(n_883), .Y(n_1069) );
INVx2_ASAP7_75t_L g1070 ( .A(n_967), .Y(n_1070) );
NAND3xp33_ASAP7_75t_L g1071 ( .A(n_961), .B(n_965), .C(n_883), .Y(n_1071) );
NAND3xp33_ASAP7_75t_L g1072 ( .A(n_961), .B(n_965), .C(n_947), .Y(n_1072) );
BUFx3_ASAP7_75t_L g1073 ( .A(n_925), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_980), .A2(n_958), .B1(n_948), .B2(n_970), .Y(n_1074) );
OAI22xp5_ASAP7_75t_SL g1075 ( .A1(n_897), .A2(n_871), .B1(n_976), .B2(n_894), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_963), .B(n_959), .Y(n_1076) );
OAI222xp33_ASAP7_75t_L g1077 ( .A1(n_980), .A2(n_981), .B1(n_949), .B2(n_974), .C1(n_954), .C2(n_969), .Y(n_1077) );
AOI33xp33_ASAP7_75t_L g1078 ( .A1(n_981), .A2(n_962), .A3(n_978), .B1(n_924), .B2(n_919), .B3(n_971), .Y(n_1078) );
OA21x2_ASAP7_75t_L g1079 ( .A1(n_898), .A2(n_825), .B(n_884), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_933), .A2(n_658), .B1(n_886), .B2(n_643), .Y(n_1080) );
HB1xp67_ASAP7_75t_L g1081 ( .A(n_880), .Y(n_1081) );
OA21x2_ASAP7_75t_L g1082 ( .A1(n_884), .A2(n_825), .B(n_878), .Y(n_1082) );
AND2x2_ASAP7_75t_SL g1083 ( .A(n_886), .B(n_846), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g1084 ( .A(n_880), .Y(n_1084) );
INVx3_ASAP7_75t_L g1085 ( .A(n_867), .Y(n_1085) );
NOR2xp33_ASAP7_75t_L g1086 ( .A(n_864), .B(n_565), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_977), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1034), .B(n_986), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1034), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1020), .Y(n_1090) );
INVx2_ASAP7_75t_SL g1091 ( .A(n_1013), .Y(n_1091) );
OAI31xp33_ASAP7_75t_L g1092 ( .A1(n_1010), .A2(n_1061), .A3(n_1018), .B(n_1080), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1020), .Y(n_1093) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_1039), .A2(n_1040), .B1(n_1018), .B2(n_1086), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_985), .B(n_1047), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1029), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_990), .Y(n_1097) );
OAI33xp33_ASAP7_75t_L g1098 ( .A1(n_1029), .A2(n_1030), .A3(n_1054), .B1(n_1051), .B2(n_1048), .B3(n_993), .Y(n_1098) );
INVx5_ASAP7_75t_SL g1099 ( .A(n_1083), .Y(n_1099) );
NAND3xp33_ASAP7_75t_L g1100 ( .A(n_1044), .B(n_1045), .C(n_1033), .Y(n_1100) );
CKINVDCx20_ASAP7_75t_R g1101 ( .A(n_1050), .Y(n_1101) );
INVx2_ASAP7_75t_L g1102 ( .A(n_990), .Y(n_1102) );
INVx2_ASAP7_75t_L g1103 ( .A(n_997), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1030), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_985), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_986), .B(n_1041), .Y(n_1106) );
NOR2xp33_ASAP7_75t_L g1107 ( .A(n_1050), .B(n_1046), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1087), .Y(n_1108) );
NOR2xp33_ASAP7_75t_L g1109 ( .A(n_1046), .B(n_1055), .Y(n_1109) );
NAND3xp33_ASAP7_75t_L g1110 ( .A(n_1044), .B(n_1019), .C(n_1016), .Y(n_1110) );
AO21x2_ASAP7_75t_L g1111 ( .A1(n_1026), .A2(n_1028), .B(n_1070), .Y(n_1111) );
NOR2xp67_ASAP7_75t_L g1112 ( .A(n_1071), .B(n_1072), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1041), .B(n_997), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1087), .B(n_1051), .Y(n_1114) );
NOR3xp33_ASAP7_75t_L g1115 ( .A(n_988), .B(n_1063), .C(n_996), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_1081), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1000), .Y(n_1117) );
OAI22xp5_ASAP7_75t_SL g1118 ( .A1(n_1083), .A2(n_1056), .B1(n_1073), .B2(n_1055), .Y(n_1118) );
OAI221xp5_ASAP7_75t_L g1119 ( .A1(n_1053), .A2(n_1057), .B1(n_1042), .B2(n_1059), .C(n_1001), .Y(n_1119) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_1084), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1000), .B(n_1003), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_995), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1123 ( .A(n_989), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1003), .B(n_995), .Y(n_1124) );
NOR3xp33_ASAP7_75t_L g1125 ( .A(n_999), .B(n_1065), .C(n_1017), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_984), .B(n_989), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1009), .B(n_984), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1049), .Y(n_1128) );
NAND3xp33_ASAP7_75t_L g1129 ( .A(n_1071), .B(n_1074), .C(n_1072), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1009), .B(n_1052), .Y(n_1130) );
AND2x4_ASAP7_75t_L g1131 ( .A(n_1085), .B(n_1060), .Y(n_1131) );
NAND4xp25_ASAP7_75t_L g1132 ( .A(n_1043), .B(n_998), .C(n_987), .D(n_992), .Y(n_1132) );
OAI22xp5_ASAP7_75t_SL g1133 ( .A1(n_1083), .A2(n_1056), .B1(n_1073), .B2(n_1075), .Y(n_1133) );
OAI211xp5_ASAP7_75t_L g1134 ( .A1(n_1068), .A2(n_1032), .B(n_1062), .C(n_1037), .Y(n_1134) );
INVx3_ASAP7_75t_L g1135 ( .A(n_1085), .Y(n_1135) );
INVx2_ASAP7_75t_L g1136 ( .A(n_1025), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_994), .B(n_1068), .Y(n_1137) );
OR2x2_ASAP7_75t_L g1138 ( .A(n_1013), .B(n_1064), .Y(n_1138) );
NAND2xp5_ASAP7_75t_SL g1139 ( .A(n_1085), .B(n_1031), .Y(n_1139) );
NAND2xp5_ASAP7_75t_SL g1140 ( .A(n_1031), .B(n_1075), .Y(n_1140) );
AND2x4_ASAP7_75t_L g1141 ( .A(n_1060), .B(n_1011), .Y(n_1141) );
INVx2_ASAP7_75t_L g1142 ( .A(n_1025), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1049), .Y(n_1143) );
NOR2xp33_ASAP7_75t_L g1144 ( .A(n_994), .B(n_1022), .Y(n_1144) );
NOR3xp33_ASAP7_75t_L g1145 ( .A(n_1007), .B(n_1006), .C(n_1035), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1052), .Y(n_1146) );
INVxp67_ASAP7_75t_SL g1147 ( .A(n_1058), .Y(n_1147) );
NOR2xp33_ASAP7_75t_L g1148 ( .A(n_1021), .B(n_1022), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1058), .B(n_1064), .Y(n_1149) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_1021), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1026), .Y(n_1151) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1028), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1060), .B(n_1082), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1060), .B(n_1082), .Y(n_1154) );
HB1xp67_ASAP7_75t_L g1155 ( .A(n_1023), .Y(n_1155) );
NOR2xp67_ASAP7_75t_L g1156 ( .A(n_1036), .B(n_1002), .Y(n_1156) );
INVx4_ASAP7_75t_L g1157 ( .A(n_1015), .Y(n_1157) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1066), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1082), .B(n_1012), .Y(n_1159) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1066), .Y(n_1160) );
OAI211xp5_ASAP7_75t_L g1161 ( .A1(n_1024), .A2(n_1038), .B(n_1014), .C(n_1008), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_1012), .A2(n_1076), .B1(n_1069), .B2(n_1002), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1070), .Y(n_1163) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1082), .Y(n_1164) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_1076), .A2(n_1027), .B1(n_1015), .B2(n_1067), .Y(n_1165) );
INVx2_ASAP7_75t_L g1166 ( .A(n_1079), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1004), .B(n_1067), .Y(n_1167) );
OAI211xp5_ASAP7_75t_L g1168 ( .A1(n_1067), .A2(n_1079), .B(n_991), .C(n_1005), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1067), .B(n_1015), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1005), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1078), .B(n_1004), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1004), .B(n_1079), .Y(n_1172) );
BUFx2_ASAP7_75t_L g1173 ( .A(n_1079), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_991), .Y(n_1174) );
OAI21xp5_ASAP7_75t_L g1175 ( .A1(n_1129), .A2(n_1077), .B(n_1112), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1095), .B(n_1106), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1177 ( .A(n_1095), .B(n_1106), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1130), .B(n_1088), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1090), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1130), .B(n_1088), .Y(n_1180) );
INVx1_ASAP7_75t_SL g1181 ( .A(n_1101), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1090), .Y(n_1182) );
OR2x6_ASAP7_75t_L g1183 ( .A(n_1141), .B(n_1131), .Y(n_1183) );
AND4x1_ASAP7_75t_L g1184 ( .A(n_1107), .B(n_1092), .C(n_1100), .D(n_1115), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1089), .B(n_1127), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1089), .B(n_1127), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1093), .Y(n_1187) );
INVx2_ASAP7_75t_L g1188 ( .A(n_1136), .Y(n_1188) );
HB1xp67_ASAP7_75t_L g1189 ( .A(n_1116), .Y(n_1189) );
NOR2xp33_ASAP7_75t_L g1190 ( .A(n_1132), .B(n_1094), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1113), .B(n_1096), .Y(n_1191) );
BUFx2_ASAP7_75t_L g1192 ( .A(n_1101), .Y(n_1192) );
OR2x2_ASAP7_75t_L g1193 ( .A(n_1123), .B(n_1138), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1113), .B(n_1108), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1104), .Y(n_1195) );
OAI22xp33_ASAP7_75t_SL g1196 ( .A1(n_1140), .A2(n_1119), .B1(n_1120), .B2(n_1109), .Y(n_1196) );
INVxp67_ASAP7_75t_SL g1197 ( .A(n_1150), .Y(n_1197) );
AND2x4_ASAP7_75t_L g1198 ( .A(n_1131), .B(n_1141), .Y(n_1198) );
NAND4xp25_ASAP7_75t_L g1199 ( .A(n_1162), .B(n_1110), .C(n_1156), .D(n_1145), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1138), .B(n_1105), .Y(n_1200) );
OAI221xp5_ASAP7_75t_L g1201 ( .A1(n_1133), .A2(n_1125), .B1(n_1155), .B2(n_1161), .C(n_1134), .Y(n_1201) );
OR2x2_ASAP7_75t_L g1202 ( .A(n_1126), .B(n_1091), .Y(n_1202) );
BUFx2_ASAP7_75t_L g1203 ( .A(n_1091), .Y(n_1203) );
NOR2xp33_ASAP7_75t_L g1204 ( .A(n_1098), .B(n_1114), .Y(n_1204) );
NAND4xp25_ASAP7_75t_L g1205 ( .A(n_1144), .B(n_1137), .C(n_1148), .D(n_1159), .Y(n_1205) );
INVx1_ASAP7_75t_SL g1206 ( .A(n_1124), .Y(n_1206) );
INVx1_ASAP7_75t_SL g1207 ( .A(n_1124), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1121), .B(n_1149), .Y(n_1208) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1136), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1122), .B(n_1121), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1149), .B(n_1167), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1117), .B(n_1097), .Y(n_1212) );
INVx1_ASAP7_75t_SL g1213 ( .A(n_1118), .Y(n_1213) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1142), .Y(n_1214) );
AND2x4_ASAP7_75t_L g1215 ( .A(n_1131), .B(n_1141), .Y(n_1215) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_1139), .A2(n_1099), .B1(n_1165), .B2(n_1170), .Y(n_1216) );
NAND4xp25_ASAP7_75t_SL g1217 ( .A(n_1159), .B(n_1168), .C(n_1154), .D(n_1153), .Y(n_1217) );
NOR2xp33_ASAP7_75t_L g1218 ( .A(n_1135), .B(n_1171), .Y(n_1218) );
OR2x2_ASAP7_75t_L g1219 ( .A(n_1097), .B(n_1102), .Y(n_1219) );
HB1xp67_ASAP7_75t_L g1220 ( .A(n_1102), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1103), .Y(n_1221) );
OR2x2_ASAP7_75t_L g1222 ( .A(n_1103), .B(n_1128), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1167), .B(n_1154), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1153), .B(n_1172), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1172), .B(n_1143), .Y(n_1225) );
NOR2x1_ASAP7_75t_L g1226 ( .A(n_1135), .B(n_1157), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1146), .B(n_1163), .Y(n_1227) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1146), .B(n_1163), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1151), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1142), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1135), .B(n_1151), .Y(n_1231) );
NAND4xp25_ASAP7_75t_L g1232 ( .A(n_1169), .B(n_1173), .C(n_1157), .D(n_1164), .Y(n_1232) );
INVx3_ASAP7_75t_SL g1233 ( .A(n_1157), .Y(n_1233) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1188), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1179), .Y(n_1235) );
OR2x6_ASAP7_75t_L g1236 ( .A(n_1183), .B(n_1164), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1211), .B(n_1173), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1182), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1187), .Y(n_1239) );
INVx1_ASAP7_75t_SL g1240 ( .A(n_1192), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1204), .B(n_1158), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1204), .B(n_1158), .Y(n_1242) );
INVxp67_ASAP7_75t_SL g1243 ( .A(n_1220), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1191), .B(n_1160), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1191), .B(n_1160), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1194), .B(n_1152), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1228), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1211), .B(n_1147), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1224), .B(n_1166), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1224), .B(n_1166), .Y(n_1250) );
NAND2xp5_ASAP7_75t_SL g1251 ( .A(n_1196), .B(n_1099), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1228), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1223), .B(n_1152), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1229), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1194), .B(n_1174), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1227), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1185), .B(n_1186), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1223), .B(n_1111), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1227), .Y(n_1259) );
OAI22xp5_ASAP7_75t_L g1260 ( .A1(n_1201), .A2(n_1099), .B1(n_1174), .B2(n_1111), .Y(n_1260) );
A2O1A1Ixp33_ASAP7_75t_L g1261 ( .A1(n_1190), .A2(n_1099), .B(n_1111), .C(n_1175), .Y(n_1261) );
INVxp67_ASAP7_75t_L g1262 ( .A(n_1189), .Y(n_1262) );
INVxp67_ASAP7_75t_SL g1263 ( .A(n_1197), .Y(n_1263) );
INVx1_ASAP7_75t_SL g1264 ( .A(n_1181), .Y(n_1264) );
NOR3xp33_ASAP7_75t_L g1265 ( .A(n_1199), .B(n_1190), .C(n_1213), .Y(n_1265) );
AOI322xp5_ASAP7_75t_L g1266 ( .A1(n_1185), .A2(n_1186), .A3(n_1178), .B1(n_1180), .B2(n_1206), .C1(n_1207), .C2(n_1200), .Y(n_1266) );
INVx1_ASAP7_75t_SL g1267 ( .A(n_1176), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1200), .B(n_1176), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1208), .B(n_1178), .Y(n_1269) );
NOR2xp33_ASAP7_75t_L g1270 ( .A(n_1240), .B(n_1184), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1241), .B(n_1180), .Y(n_1271) );
INVx1_ASAP7_75t_SL g1272 ( .A(n_1264), .Y(n_1272) );
NAND2x1_ASAP7_75t_L g1273 ( .A(n_1236), .B(n_1183), .Y(n_1273) );
OA21x2_ASAP7_75t_L g1274 ( .A1(n_1261), .A2(n_1232), .B(n_1218), .Y(n_1274) );
XNOR2xp5_ASAP7_75t_L g1275 ( .A(n_1265), .B(n_1205), .Y(n_1275) );
NOR2xp33_ASAP7_75t_SL g1276 ( .A(n_1263), .B(n_1203), .Y(n_1276) );
INVx1_ASAP7_75t_SL g1277 ( .A(n_1267), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1258), .B(n_1208), .Y(n_1278) );
NAND3xp33_ASAP7_75t_L g1279 ( .A(n_1260), .B(n_1218), .C(n_1216), .Y(n_1279) );
NAND3xp33_ASAP7_75t_L g1280 ( .A(n_1242), .B(n_1226), .C(n_1231), .Y(n_1280) );
OAI22xp5_ASAP7_75t_L g1281 ( .A1(n_1251), .A2(n_1177), .B1(n_1202), .B2(n_1183), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1235), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1235), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1258), .B(n_1225), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1238), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1269), .B(n_1225), .Y(n_1286) );
INVx1_ASAP7_75t_SL g1287 ( .A(n_1269), .Y(n_1287) );
OAI21xp5_ASAP7_75t_SL g1288 ( .A1(n_1266), .A2(n_1215), .B(n_1198), .Y(n_1288) );
NOR2xp33_ASAP7_75t_L g1289 ( .A(n_1262), .B(n_1177), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1249), .B(n_1183), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1238), .Y(n_1291) );
NAND2xp5_ASAP7_75t_SL g1292 ( .A(n_1243), .B(n_1233), .Y(n_1292) );
NOR2xp67_ASAP7_75t_SL g1293 ( .A(n_1248), .B(n_1193), .Y(n_1293) );
NOR2xp33_ASAP7_75t_L g1294 ( .A(n_1257), .B(n_1195), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1247), .Y(n_1295) );
INVx2_ASAP7_75t_SL g1296 ( .A(n_1248), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1247), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1249), .B(n_1215), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1252), .B(n_1259), .Y(n_1299) );
HB1xp67_ASAP7_75t_L g1300 ( .A(n_1253), .Y(n_1300) );
NOR3xp33_ASAP7_75t_SL g1301 ( .A(n_1255), .B(n_1217), .C(n_1210), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1252), .Y(n_1302) );
NAND2xp5_ASAP7_75t_SL g1303 ( .A(n_1234), .B(n_1233), .Y(n_1303) );
INVx2_ASAP7_75t_SL g1304 ( .A(n_1253), .Y(n_1304) );
XNOR2xp5_ASAP7_75t_L g1305 ( .A(n_1268), .B(n_1215), .Y(n_1305) );
XNOR2x2_ASAP7_75t_L g1306 ( .A(n_1244), .B(n_1193), .Y(n_1306) );
NOR2xp33_ASAP7_75t_L g1307 ( .A(n_1256), .B(n_1198), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1237), .B(n_1198), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1256), .Y(n_1309) );
NOR2x1_ASAP7_75t_L g1310 ( .A(n_1236), .B(n_1222), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1259), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1239), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1239), .Y(n_1313) );
NOR3xp33_ASAP7_75t_L g1314 ( .A(n_1254), .B(n_1212), .C(n_1221), .Y(n_1314) );
NOR2xp33_ASAP7_75t_L g1315 ( .A(n_1237), .B(n_1222), .Y(n_1315) );
AOI21xp5_ASAP7_75t_L g1316 ( .A1(n_1236), .A2(n_1219), .B(n_1214), .Y(n_1316) );
INVx1_ASAP7_75t_SL g1317 ( .A(n_1245), .Y(n_1317) );
AOI22xp5_ASAP7_75t_L g1318 ( .A1(n_1236), .A2(n_1209), .B1(n_1214), .B2(n_1230), .Y(n_1318) );
XOR2xp5_ASAP7_75t_SL g1319 ( .A(n_1250), .B(n_1219), .Y(n_1319) );
INVx2_ASAP7_75t_L g1320 ( .A(n_1304), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1299), .Y(n_1321) );
OAI21xp5_ASAP7_75t_SL g1322 ( .A1(n_1275), .A2(n_1288), .B(n_1281), .Y(n_1322) );
AND2x4_ASAP7_75t_L g1323 ( .A(n_1310), .B(n_1273), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1300), .Y(n_1324) );
OA33x2_ASAP7_75t_L g1325 ( .A1(n_1271), .A2(n_1275), .A3(n_1246), .B1(n_1306), .B2(n_1319), .B3(n_1301), .Y(n_1325) );
OAI22xp33_ASAP7_75t_L g1326 ( .A1(n_1276), .A2(n_1273), .B1(n_1292), .B2(n_1319), .Y(n_1326) );
AOI221xp5_ASAP7_75t_L g1327 ( .A1(n_1270), .A2(n_1289), .B1(n_1294), .B2(n_1293), .C(n_1279), .Y(n_1327) );
OAI211xp5_ASAP7_75t_SL g1328 ( .A1(n_1272), .A2(n_1277), .B(n_1303), .C(n_1318), .Y(n_1328) );
NOR2x1_ASAP7_75t_SL g1329 ( .A(n_1303), .B(n_1236), .Y(n_1329) );
INVx2_ASAP7_75t_SL g1330 ( .A(n_1304), .Y(n_1330) );
OAI22xp5_ASAP7_75t_SL g1331 ( .A1(n_1274), .A2(n_1287), .B1(n_1305), .B2(n_1296), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1285), .Y(n_1332) );
NOR3x1_ASAP7_75t_L g1333 ( .A(n_1322), .B(n_1280), .C(n_1296), .Y(n_1333) );
OAI322xp33_ASAP7_75t_L g1334 ( .A1(n_1326), .A2(n_1317), .A3(n_1307), .B1(n_1295), .B2(n_1297), .C1(n_1302), .C2(n_1315), .Y(n_1334) );
NOR3xp33_ASAP7_75t_L g1335 ( .A(n_1326), .B(n_1314), .C(n_1316), .Y(n_1335) );
NAND5xp2_ASAP7_75t_L g1336 ( .A(n_1327), .B(n_1307), .C(n_1290), .D(n_1315), .E(n_1274), .Y(n_1336) );
BUFx6f_ASAP7_75t_L g1337 ( .A(n_1330), .Y(n_1337) );
OAI221xp5_ASAP7_75t_SL g1338 ( .A1(n_1325), .A2(n_1290), .B1(n_1311), .B2(n_1309), .C(n_1308), .Y(n_1338) );
NOR3x1_ASAP7_75t_L g1339 ( .A(n_1331), .B(n_1274), .C(n_1293), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1321), .B(n_1286), .Y(n_1340) );
OA22x2_ASAP7_75t_L g1341 ( .A1(n_1323), .A2(n_1286), .B1(n_1298), .B2(n_1278), .Y(n_1341) );
NAND3xp33_ASAP7_75t_SL g1342 ( .A(n_1335), .B(n_1328), .C(n_1320), .Y(n_1342) );
NAND4xp25_ASAP7_75t_L g1343 ( .A(n_1333), .B(n_1328), .C(n_1323), .D(n_1324), .Y(n_1343) );
NOR4xp25_ASAP7_75t_L g1344 ( .A(n_1334), .B(n_1320), .C(n_1332), .D(n_1313), .Y(n_1344) );
OR2x2_ASAP7_75t_L g1345 ( .A(n_1340), .B(n_1278), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1337), .B(n_1284), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1337), .B(n_1284), .Y(n_1347) );
OAI22xp5_ASAP7_75t_L g1348 ( .A1(n_1346), .A2(n_1341), .B1(n_1338), .B2(n_1336), .Y(n_1348) );
AOI21xp5_ASAP7_75t_L g1349 ( .A1(n_1342), .A2(n_1329), .B(n_1274), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1347), .Y(n_1350) );
OAI221xp5_ASAP7_75t_L g1351 ( .A1(n_1343), .A2(n_1339), .B1(n_1312), .B2(n_1282), .C(n_1291), .Y(n_1351) );
INVx2_ASAP7_75t_L g1352 ( .A(n_1345), .Y(n_1352) );
INVx2_ASAP7_75t_SL g1353 ( .A(n_1350), .Y(n_1353) );
XNOR2xp5_ASAP7_75t_L g1354 ( .A(n_1349), .B(n_1344), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1352), .B(n_1283), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1351), .Y(n_1356) );
OR3x1_ASAP7_75t_L g1357 ( .A(n_1356), .B(n_1348), .C(n_1291), .Y(n_1357) );
BUFx2_ASAP7_75t_L g1358 ( .A(n_1353), .Y(n_1358) );
XNOR2xp5_ASAP7_75t_L g1359 ( .A(n_1357), .B(n_1354), .Y(n_1359) );
AOI221xp5_ASAP7_75t_L g1360 ( .A1(n_1358), .A2(n_1355), .B1(n_1285), .B2(n_1283), .C(n_1282), .Y(n_1360) );
INVxp67_ASAP7_75t_L g1361 ( .A(n_1359), .Y(n_1361) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_1361), .A2(n_1360), .B1(n_1250), .B2(n_1234), .Y(n_1362) );
endmodule