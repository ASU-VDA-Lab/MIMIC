module fake_jpeg_7115_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_34),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_40),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_13),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_32),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_28),
.B1(n_31),
.B2(n_25),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_68),
.B1(n_23),
.B2(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_16),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_61),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_49),
.B(n_9),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_25),
.B1(n_31),
.B2(n_16),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_27),
.C(n_21),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_19),
.B1(n_29),
.B2(n_26),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_62),
.B1(n_23),
.B2(n_21),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_28),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_29),
.B1(n_26),
.B2(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_39),
.A2(n_17),
.B1(n_27),
.B2(n_32),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_66),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_71),
.B(n_83),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_82),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_39),
.B(n_30),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_48),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_21),
.B1(n_27),
.B2(n_20),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_48),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_50),
.B1(n_61),
.B2(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_44),
.A2(n_61),
.B1(n_52),
.B2(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_20),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_53),
.Y(n_118)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_93),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_44),
.A2(n_21),
.B1(n_27),
.B2(n_30),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_49),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_111),
.Y(n_124)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_81),
.B1(n_74),
.B2(n_71),
.Y(n_121)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_105),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_53),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_118),
.Y(n_129)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_47),
.B1(n_92),
.B2(n_63),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_107),
.A2(n_83),
.B1(n_78),
.B2(n_75),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_134),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_73),
.B1(n_87),
.B2(n_88),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_80),
.B1(n_73),
.B2(n_86),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_139),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_51),
.B(n_69),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_133),
.B(n_137),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_57),
.B(n_59),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_86),
.B1(n_59),
.B2(n_65),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_69),
.B(n_89),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_79),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_98),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_53),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_101),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_95),
.A2(n_88),
.B1(n_103),
.B2(n_111),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_103),
.B1(n_76),
.B2(n_104),
.Y(n_157)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_138),
.B(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_154),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_152),
.A2(n_166),
.B(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_113),
.Y(n_156)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_125),
.B(n_30),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_134),
.B(n_98),
.Y(n_161)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_140),
.A2(n_141),
.B1(n_124),
.B2(n_120),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_163),
.A2(n_67),
.B1(n_27),
.B2(n_57),
.Y(n_191)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_168),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_130),
.B(n_115),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_172),
.B(n_152),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_121),
.B1(n_142),
.B2(n_133),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_173),
.A2(n_178),
.B1(n_190),
.B2(n_197),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_189),
.B(n_192),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_176),
.B(n_191),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_135),
.C(n_127),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_198),
.C(n_157),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_125),
.B1(n_127),
.B2(n_119),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_171),
.A2(n_146),
.B1(n_76),
.B2(n_145),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_179),
.A2(n_161),
.B(n_172),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_180),
.B(n_188),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_146),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_195),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_116),
.B1(n_112),
.B2(n_54),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_164),
.B1(n_165),
.B2(n_158),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_54),
.B1(n_109),
.B2(n_64),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_67),
.B(n_20),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_67),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_109),
.B1(n_132),
.B2(n_105),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_132),
.C(n_105),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_193),
.B(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_185),
.B(n_148),
.Y(n_200)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_214),
.B1(n_174),
.B2(n_190),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_115),
.Y(n_202)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_194),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_206),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_181),
.B(n_148),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_205),
.B(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_166),
.C(n_162),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_154),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_212),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_149),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_20),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_189),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_175),
.A2(n_150),
.B1(n_147),
.B2(n_155),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_158),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_217),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_221),
.B(n_192),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_220),
.C(n_160),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_184),
.C(n_177),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_162),
.B(n_168),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_181),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_222),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_167),
.Y(n_223)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_232),
.C(n_233),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_228),
.A2(n_230),
.B1(n_215),
.B2(n_201),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_241),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_178),
.B1(n_196),
.B2(n_198),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_191),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_239),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_162),
.C(n_157),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_180),
.C(n_196),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_20),
.C(n_18),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_219),
.C(n_211),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_18),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_18),
.Y(n_243)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_206),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_226),
.Y(n_248)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_256),
.C(n_4),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_SL g252 ( 
.A1(n_229),
.A2(n_204),
.B(n_215),
.C(n_207),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_252),
.A2(n_253),
.B(n_0),
.Y(n_270)
);

OAI21x1_ASAP7_75t_SL g253 ( 
.A1(n_233),
.A2(n_204),
.B(n_218),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_216),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_254),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_214),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_260),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_210),
.C(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_216),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_4),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_259),
.A2(n_261),
.B1(n_235),
.B2(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_239),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_274),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_267),
.B1(n_273),
.B2(n_271),
.Y(n_289)
);

OAI321xp33_ASAP7_75t_L g265 ( 
.A1(n_252),
.A2(n_242),
.A3(n_227),
.B1(n_238),
.B2(n_231),
.C(n_241),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_270),
.B(n_275),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_232),
.B1(n_234),
.B2(n_3),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_273),
.B1(n_247),
.B2(n_251),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_252),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_2),
.B(n_3),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_9),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_266),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_250),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_281),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_245),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_280),
.B(n_286),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_257),
.Y(n_280)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_247),
.Y(n_283)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_250),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_287),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_269),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_9),
.Y(n_287)
);

OAI21x1_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_8),
.B(n_12),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_8),
.B(n_12),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_4),
.Y(n_292)
);

A2O1A1O1Ixp25_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_268),
.B(n_263),
.C(n_267),
.D(n_11),
.Y(n_291)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_292),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_8),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_4),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_5),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_284),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_303),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_294),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_306),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_277),
.C(n_10),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_305),
.A2(n_10),
.B(n_13),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_293),
.B1(n_299),
.B2(n_277),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_309),
.C(n_307),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_302),
.A2(n_5),
.B(n_6),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_5),
.B(n_6),
.Y(n_311)
);

AO21x1_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_300),
.B(n_6),
.Y(n_314)
);

OAI211xp5_ASAP7_75t_SL g315 ( 
.A1(n_313),
.A2(n_314),
.B(n_312),
.C(n_310),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_6),
.B(n_7),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_7),
.C(n_267),
.Y(n_317)
);


endmodule