module fake_jpeg_3205_n_492 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_492);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_492;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_56),
.Y(n_104)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_53),
.Y(n_121)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_55),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_16),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_15),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_66),
.B(n_68),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_0),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_17),
.B(n_1),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_1),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_77),
.B(n_83),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_17),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_90),
.Y(n_111)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_2),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

AND2x4_ASAP7_75t_SL g87 ( 
.A(n_18),
.B(n_2),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_97),
.Y(n_99)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_3),
.Y(n_90)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

BUFx8_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g148 ( 
.A(n_94),
.Y(n_148)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

CKINVDCx11_ASAP7_75t_R g100 ( 
.A(n_94),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_100),
.B(n_117),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_101),
.B(n_115),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_29),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_29),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_57),
.B(n_50),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_119),
.B(n_123),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_50),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_28),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_124),
.B(n_125),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_28),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_32),
.C(n_20),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_11),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_82),
.A2(n_30),
.B1(n_46),
.B2(n_38),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_130),
.A2(n_134),
.B1(n_154),
.B2(n_159),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_49),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_133),
.B(n_144),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_84),
.A2(n_30),
.B1(n_46),
.B2(n_38),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_54),
.B(n_49),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_137),
.B(n_140),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_70),
.B(n_37),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_37),
.Y(n_142)
);

NAND2xp33_ASAP7_75t_SL g220 ( 
.A(n_142),
.B(n_118),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_97),
.Y(n_144)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_73),
.B(n_36),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_62),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_154)
);

BUFx10_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_91),
.A2(n_30),
.B1(n_27),
.B2(n_26),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_142),
.A2(n_34),
.B1(n_25),
.B2(n_40),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_161),
.B(n_202),
.Y(n_243)
);

BUFx2_ASAP7_75t_SL g164 ( 
.A(n_98),
.Y(n_164)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_151),
.A2(n_38),
.B1(n_46),
.B2(n_27),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_166),
.A2(n_173),
.B1(n_175),
.B2(n_196),
.Y(n_246)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_168),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_110),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_170),
.B(n_213),
.Y(n_254)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_171),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_27),
.B1(n_21),
.B2(n_26),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_99),
.B(n_26),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_177),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_106),
.A2(n_35),
.B1(n_44),
.B2(n_43),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_99),
.B(n_75),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_176),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_74),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_104),
.B(n_34),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_184),
.Y(n_232)
);

NOR2x1_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_89),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_180),
.B(n_215),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_108),
.A2(n_25),
.B1(n_35),
.B2(n_44),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_181),
.A2(n_186),
.B1(n_103),
.B2(n_116),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_L g183 ( 
.A1(n_130),
.A2(n_40),
.B1(n_36),
.B2(n_43),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_183),
.A2(n_187),
.B1(n_201),
.B2(n_215),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_120),
.B(n_39),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_185),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_39),
.B1(n_65),
.B2(n_88),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_47),
.B1(n_22),
.B2(n_7),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_126),
.B(n_5),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_200),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_199),
.Y(n_227)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_191),
.Y(n_268)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_136),
.A2(n_47),
.B1(n_6),
.B2(n_7),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

AOI32xp33_ASAP7_75t_L g199 ( 
.A1(n_111),
.A2(n_47),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_113),
.B(n_5),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_134),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_114),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_220),
.Y(n_252)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_204),
.Y(n_257)
);

INVx11_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_205),
.Y(n_265)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_207),
.Y(n_260)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_209),
.Y(n_269)
);

AO22x1_ASAP7_75t_SL g211 ( 
.A1(n_138),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_211)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_98),
.B(n_12),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_216),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_155),
.A2(n_13),
.B(n_148),
.C(n_122),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_141),
.B(n_13),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_121),
.C(n_118),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_112),
.A2(n_132),
.B1(n_105),
.B2(n_138),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_141),
.B(n_105),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_132),
.A2(n_122),
.B1(n_139),
.B2(n_127),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_217),
.A2(n_219),
.B1(n_150),
.B2(n_109),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_127),
.A2(n_131),
.B1(n_146),
.B2(n_156),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_155),
.A2(n_148),
.B(n_135),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_221),
.A2(n_213),
.B(n_183),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_121),
.B1(n_135),
.B2(n_109),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_222),
.A2(n_263),
.B1(n_240),
.B2(n_237),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_224),
.B(n_247),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_225),
.A2(n_276),
.B1(n_194),
.B2(n_209),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_176),
.A2(n_131),
.B1(n_146),
.B2(n_156),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_228),
.A2(n_261),
.B1(n_267),
.B2(n_163),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_178),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_229),
.B(n_230),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_189),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_161),
.A2(n_129),
.B1(n_116),
.B2(n_103),
.Y(n_231)
);

A2O1A1Ixp33_ASAP7_75t_SL g301 ( 
.A1(n_231),
.A2(n_228),
.B(n_252),
.C(n_224),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_172),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_234),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_184),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_239),
.B(n_274),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_172),
.B(n_129),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_244),
.B(n_250),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_249),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_195),
.B(n_210),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_188),
.B(n_177),
.C(n_176),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_251),
.B(n_259),
.C(n_243),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_169),
.B(n_180),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_253),
.B(n_258),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_179),
.B(n_206),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_256),
.B(n_229),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_200),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_203),
.B(n_174),
.C(n_216),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_203),
.A2(n_202),
.B1(n_187),
.B2(n_217),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_185),
.B(n_198),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_262),
.B(n_273),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_165),
.A2(n_221),
.B1(n_167),
.B2(n_211),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_171),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g316 ( 
.A(n_264),
.B(n_275),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_214),
.A2(n_201),
.B1(n_207),
.B2(n_211),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_193),
.B(n_162),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_191),
.B(n_162),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_204),
.A2(n_208),
.B1(n_205),
.B2(n_193),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_279),
.B(n_290),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_163),
.B(n_218),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_280),
.A2(n_317),
.B(n_301),
.Y(n_341)
);

BUFx24_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_281),
.Y(n_343)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_283),
.A2(n_286),
.B1(n_295),
.B2(n_305),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_274),
.B(n_272),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_284),
.A2(n_291),
.B(n_300),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_272),
.A2(n_223),
.B1(n_239),
.B2(n_245),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_236),
.Y(n_288)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_289),
.B(n_308),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_238),
.B(n_242),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_235),
.Y(n_292)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_230),
.B(n_248),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_293),
.B(n_294),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_236),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_223),
.A2(n_271),
.B1(n_242),
.B2(n_238),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_241),
.B(n_232),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_296),
.B(n_298),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_232),
.B(n_251),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_297),
.B(n_300),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_259),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_252),
.B(n_264),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g331 ( 
.A1(n_301),
.A2(n_240),
.B(n_226),
.Y(n_331)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_260),
.Y(n_302)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_302),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_252),
.B(n_264),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_303),
.B(n_268),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_271),
.A2(n_227),
.B1(n_243),
.B2(n_246),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_231),
.B(n_261),
.Y(n_307)
);

AND2x2_ASAP7_75t_SL g352 ( 
.A(n_307),
.B(n_317),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_255),
.B(n_266),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_233),
.Y(n_309)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_311),
.B(n_303),
.C(n_316),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_243),
.A2(n_267),
.B1(n_231),
.B2(n_225),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_312),
.A2(n_307),
.B1(n_285),
.B2(n_314),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_255),
.B(n_257),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_318),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_231),
.B(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_257),
.B(n_270),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_320),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_235),
.Y(n_320)
);

AND2x2_ASAP7_75t_SL g321 ( 
.A(n_237),
.B(n_268),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_321),
.Y(n_329)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_233),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_309),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_323),
.A2(n_226),
.B1(n_269),
.B2(n_312),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_326),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_269),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_327),
.B(n_358),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_321),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_330),
.B(n_333),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_331),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_290),
.B(n_295),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_336),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_337),
.A2(n_344),
.B(n_346),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_339),
.A2(n_342),
.B1(n_316),
.B2(n_289),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_341),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_307),
.A2(n_283),
.B1(n_305),
.B2(n_286),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_284),
.B(n_291),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_280),
.A2(n_317),
.B(n_285),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_285),
.A2(n_301),
.B1(n_296),
.B2(n_298),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_350),
.A2(n_361),
.B1(n_323),
.B2(n_282),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_313),
.C(n_318),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_297),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_360),
.Y(n_366)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_287),
.B(n_304),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_287),
.B(n_279),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_301),
.A2(n_316),
.B1(n_311),
.B2(n_306),
.Y(n_361)
);

OAI32xp33_ASAP7_75t_L g362 ( 
.A1(n_301),
.A2(n_293),
.A3(n_324),
.B1(n_294),
.B2(n_319),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_362),
.B(n_316),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_364),
.A2(n_372),
.B1(n_385),
.B2(n_390),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_365),
.B(n_382),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_362),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_359),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_379),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_332),
.A2(n_342),
.B1(n_339),
.B2(n_336),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_355),
.Y(n_374)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_348),
.B(n_308),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_375),
.B(n_378),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_326),
.C(n_331),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_322),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_334),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_332),
.A2(n_288),
.B1(n_322),
.B2(n_310),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_380),
.A2(n_328),
.B1(n_354),
.B2(n_331),
.Y(n_405)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_355),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_383),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_320),
.Y(n_382)
);

OAI32xp33_ASAP7_75t_L g383 ( 
.A1(n_345),
.A2(n_302),
.A3(n_321),
.B1(n_299),
.B2(n_281),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_346),
.A2(n_321),
.B1(n_281),
.B2(n_292),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_325),
.B(n_281),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_386),
.B(n_338),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_347),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_391),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_352),
.A2(n_333),
.B1(n_341),
.B2(n_325),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_352),
.A2(n_344),
.B1(n_337),
.B2(n_358),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_350),
.B(n_347),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_392),
.B(n_349),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_356),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_340),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_340),
.Y(n_394)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_359),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_395),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_396),
.A2(n_404),
.B1(n_405),
.B2(n_409),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_349),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_397),
.Y(n_431)
);

AOI322xp5_ASAP7_75t_SL g399 ( 
.A1(n_366),
.A2(n_353),
.A3(n_361),
.B1(n_356),
.B2(n_351),
.C1(n_329),
.C2(n_330),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_399),
.B(n_419),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_352),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_412),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_403),
.C(n_414),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_352),
.C(n_331),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_387),
.A2(n_335),
.B1(n_329),
.B2(n_328),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_373),
.A2(n_335),
.B1(n_354),
.B2(n_357),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_410),
.Y(n_432)
);

AND2x6_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_343),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_385),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_363),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_415),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_386),
.B(n_335),
.C(n_338),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_340),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_374),
.B(n_381),
.Y(n_419)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_421),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_422),
.A2(n_427),
.B1(n_429),
.B2(n_438),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_389),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_425),
.B(n_430),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_404),
.A2(n_372),
.B1(n_367),
.B2(n_364),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_408),
.A2(n_367),
.B1(n_368),
.B2(n_370),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_369),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_388),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_407),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_400),
.C(n_412),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_436),
.B(n_437),
.C(n_433),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_403),
.B(n_384),
.C(n_370),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_408),
.A2(n_380),
.B1(n_373),
.B2(n_384),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_406),
.Y(n_439)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_439),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_420),
.A2(n_373),
.B(n_369),
.Y(n_440)
);

OAI21xp33_ASAP7_75t_L g456 ( 
.A1(n_440),
.A2(n_437),
.B(n_422),
.Y(n_456)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_398),
.Y(n_441)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_441),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_424),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_429),
.A2(n_432),
.B1(n_438),
.B2(n_427),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_443),
.A2(n_455),
.B1(n_457),
.B2(n_428),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_398),
.Y(n_444)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_444),
.Y(n_461)
);

XOR2x1_ASAP7_75t_SL g445 ( 
.A(n_435),
.B(n_415),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_446),
.C(n_448),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_414),
.C(n_420),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_413),
.C(n_407),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_451),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_446),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_434),
.A2(n_406),
.B1(n_377),
.B2(n_411),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_453),
.A2(n_426),
.B1(n_417),
.B2(n_394),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_371),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_454),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_432),
.A2(n_383),
.B1(n_371),
.B2(n_418),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_456),
.A2(n_448),
.B(n_445),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_440),
.A2(n_379),
.B1(n_395),
.B2(n_417),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_442),
.C(n_447),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_460),
.A2(n_461),
.B1(n_463),
.B2(n_462),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_462),
.A2(n_464),
.B1(n_469),
.B2(n_463),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_443),
.A2(n_428),
.B1(n_424),
.B2(n_394),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_470),
.Y(n_471)
);

AOI322xp5_ASAP7_75t_L g468 ( 
.A1(n_450),
.A2(n_454),
.A3(n_449),
.B1(n_444),
.B2(n_451),
.C1(n_458),
.C2(n_453),
.Y(n_468)
);

INVx11_ASAP7_75t_L g472 ( 
.A(n_468),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_455),
.A2(n_449),
.B1(n_457),
.B2(n_452),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_476),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_474),
.B(n_475),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_447),
.C(n_465),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_469),
.A2(n_461),
.B1(n_464),
.B2(n_470),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_478),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_460),
.C(n_466),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_476),
.A2(n_472),
.B(n_478),
.Y(n_482)
);

AOI21x1_ASAP7_75t_SL g484 ( 
.A1(n_482),
.A2(n_483),
.B(n_481),
.Y(n_484)
);

INVx13_ASAP7_75t_L g483 ( 
.A(n_473),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_484),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_482),
.B(n_474),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_485),
.A2(n_486),
.B(n_480),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_475),
.Y(n_486)
);

AO21x1_ASAP7_75t_L g489 ( 
.A1(n_488),
.A2(n_471),
.B(n_472),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_489),
.A2(n_487),
.B(n_484),
.Y(n_490)
);

OAI321xp33_ASAP7_75t_L g491 ( 
.A1(n_490),
.A2(n_466),
.A3(n_483),
.B1(n_480),
.B2(n_477),
.C(n_471),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g492 ( 
.A(n_491),
.Y(n_492)
);


endmodule