module fake_jpeg_21940_n_206 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

OR2x2_ASAP7_75t_SL g15 ( 
.A(n_8),
.B(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVxp67_ASAP7_75t_SL g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_1),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_22),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_14),
.B1(n_18),
.B2(n_24),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_50),
.B(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_43),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_25),
.B1(n_14),
.B2(n_24),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_52),
.B1(n_53),
.B2(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_41),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_18),
.B1(n_25),
.B2(n_15),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_18),
.B1(n_25),
.B2(n_15),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_18),
.B1(n_23),
.B2(n_17),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_26),
.B1(n_23),
.B2(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_60),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_40),
.B1(n_43),
.B2(n_54),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_44),
.B1(n_50),
.B2(n_41),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_22),
.B1(n_20),
.B2(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_37),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_70),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_81),
.B1(n_56),
.B2(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_78),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_34),
.B(n_51),
.C(n_53),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_80),
.B1(n_85),
.B2(n_88),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_39),
.B1(n_38),
.B2(n_45),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_35),
.B(n_47),
.C(n_27),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_45),
.B1(n_32),
.B2(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_93),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_101),
.B1(n_74),
.B2(n_88),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_69),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_98),
.C(n_79),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_99),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_49),
.C(n_70),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_103),
.Y(n_113)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_69),
.B1(n_36),
.B2(n_37),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_49),
.B(n_65),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_55),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_101),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_74),
.B1(n_81),
.B2(n_75),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_116),
.B1(n_101),
.B2(n_102),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_120),
.C(n_123),
.Y(n_126)
);

XNOR2x2_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_78),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_118),
.B(n_92),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_95),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_79),
.C(n_76),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_87),
.C(n_89),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_106),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_121),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_127),
.B(n_136),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_135),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_97),
.C(n_102),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_109),
.C(n_86),
.Y(n_149)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_138),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_134),
.A2(n_137),
.B(n_141),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_93),
.B(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_139),
.B(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_83),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_118),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_153),
.Y(n_168)
);

AOI321xp33_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_108),
.A3(n_116),
.B1(n_124),
.B2(n_123),
.C(n_109),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_19),
.B(n_22),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_154),
.C(n_155),
.Y(n_160)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_141),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_19),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_71),
.C(n_66),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_19),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_36),
.C(n_30),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_129),
.C(n_125),
.Y(n_164)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_163),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_140),
.B1(n_129),
.B2(n_133),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_154),
.C(n_156),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_149),
.A2(n_1),
.B(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_167),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_155),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_170),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_146),
.B(n_145),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_171),
.A2(n_168),
.B(n_163),
.C(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_2),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_19),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_178),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_19),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_20),
.C(n_13),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_159),
.B(n_165),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_183),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_185),
.B1(n_187),
.B2(n_7),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_168),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_157),
.B1(n_13),
.B2(n_4),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_186),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_172),
.B(n_175),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_190),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_171),
.B(n_170),
.C(n_179),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_184),
.A2(n_6),
.B(n_7),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_7),
.C(n_8),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_194),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_199),
.Y(n_202)
);

AO21x2_ASAP7_75t_SL g197 ( 
.A1(n_191),
.A2(n_9),
.B(n_11),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_197),
.A2(n_9),
.B(n_11),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_195),
.A2(n_9),
.B(n_11),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_200),
.A2(n_202),
.B(n_197),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_197),
.C(n_198),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_204),
.Y(n_206)
);


endmodule