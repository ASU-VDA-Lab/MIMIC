module fake_netlist_1_2990_n_729 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_729);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_729;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
HB1xp67_ASAP7_75t_L g84 ( .A(n_27), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_21), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_10), .Y(n_86) );
BUFx2_ASAP7_75t_L g87 ( .A(n_34), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_43), .Y(n_88) );
INVx4_ASAP7_75t_R g89 ( .A(n_33), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_45), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_50), .Y(n_91) );
INVxp33_ASAP7_75t_SL g92 ( .A(n_42), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_78), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_20), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_52), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_79), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_63), .Y(n_98) );
INVx3_ASAP7_75t_L g99 ( .A(n_28), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_26), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_38), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_73), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_62), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_3), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_81), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_69), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_70), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_77), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_23), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_37), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_49), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_47), .Y(n_114) );
INVxp33_ASAP7_75t_SL g115 ( .A(n_44), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_1), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_13), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_41), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_32), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_82), .Y(n_120) );
OR2x2_ASAP7_75t_L g121 ( .A(n_4), .B(n_0), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_65), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_83), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_71), .Y(n_124) );
OR2x2_ASAP7_75t_L g125 ( .A(n_66), .B(n_75), .Y(n_125) );
INVxp33_ASAP7_75t_SL g126 ( .A(n_59), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_68), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_30), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_14), .Y(n_129) );
INVxp67_ASAP7_75t_SL g130 ( .A(n_58), .Y(n_130) );
NOR2xp67_ASAP7_75t_L g131 ( .A(n_24), .B(n_74), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_35), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_88), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_99), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_90), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_85), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_109), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_99), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_91), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_99), .Y(n_142) );
NOR2xp33_ASAP7_75t_R g143 ( .A(n_109), .B(n_80), .Y(n_143) );
NOR2xp33_ASAP7_75t_R g144 ( .A(n_101), .B(n_76), .Y(n_144) );
NOR2xp33_ASAP7_75t_R g145 ( .A(n_127), .B(n_72), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_91), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_100), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_100), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_94), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_113), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_93), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_87), .B(n_1), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_87), .Y(n_153) );
INVxp33_ASAP7_75t_SL g154 ( .A(n_84), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_113), .Y(n_155) );
NOR2xp33_ASAP7_75t_R g156 ( .A(n_110), .B(n_64), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_93), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_92), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_95), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_95), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_96), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_106), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_85), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_115), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_110), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_117), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_104), .B(n_2), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_96), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_121), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_97), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_142), .Y(n_173) );
BUFx8_ASAP7_75t_SL g174 ( .A(n_149), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_154), .B(n_126), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
NAND2x1p5_ASAP7_75t_L g177 ( .A(n_167), .B(n_125), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
OAI22xp33_ASAP7_75t_L g179 ( .A1(n_169), .A2(n_121), .B1(n_104), .B2(n_112), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_166), .Y(n_181) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_139), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_133), .B(n_116), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_137), .Y(n_184) );
NAND2x1p5_ASAP7_75t_L g185 ( .A(n_167), .B(n_125), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_153), .B(n_114), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_158), .B(n_114), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_162), .B(n_164), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_140), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_140), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_163), .B(n_116), .Y(n_191) );
INVxp67_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_140), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_140), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_143), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_140), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_147), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_147), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_133), .A2(n_112), .B1(n_129), .B2(n_86), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_134), .B(n_129), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_144), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_134), .B(n_123), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
NAND2x1p5_ASAP7_75t_L g204 ( .A(n_136), .B(n_132), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_148), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_148), .Y(n_207) );
INVx1_ASAP7_75t_SL g208 ( .A(n_145), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_136), .B(n_132), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_150), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_150), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_138), .B(n_118), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_155), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_138), .B(n_118), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
AOI22xp33_ASAP7_75t_SL g218 ( .A1(n_141), .A2(n_97), .B1(n_98), .B2(n_102), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_155), .Y(n_219) );
BUFx2_ASAP7_75t_L g220 ( .A(n_141), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_146), .B(n_123), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_156), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_146), .B(n_111), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_151), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_151), .A2(n_111), .B1(n_102), .B2(n_128), .Y(n_225) );
AND2x6_ASAP7_75t_L g226 ( .A(n_157), .B(n_119), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_157), .A2(n_119), .B1(n_103), .B2(n_128), .Y(n_227) );
INVxp67_ASAP7_75t_SL g228 ( .A(n_159), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_159), .B(n_108), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_165), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_160), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_165), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_165), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_192), .B(n_170), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_171), .Y(n_235) );
NOR2xp33_ASAP7_75t_R g236 ( .A(n_195), .B(n_170), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_173), .Y(n_237) );
NOR2xp33_ASAP7_75t_SL g238 ( .A(n_188), .B(n_105), .Y(n_238) );
NOR2xp33_ASAP7_75t_R g239 ( .A(n_181), .B(n_168), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_173), .Y(n_240) );
CKINVDCx16_ASAP7_75t_R g241 ( .A(n_182), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_220), .B(n_168), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_220), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_173), .Y(n_244) );
NOR2xp33_ASAP7_75t_R g245 ( .A(n_222), .B(n_160), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_204), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_184), .A2(n_161), .B1(n_130), .B2(n_98), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_173), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_197), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_171), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_228), .B(n_161), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_172), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_184), .B(n_120), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_226), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_172), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_204), .Y(n_256) );
INVxp67_ASAP7_75t_L g257 ( .A(n_174), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_204), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_183), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_226), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_183), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_175), .A2(n_120), .B1(n_103), .B2(n_124), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_230), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_226), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_183), .Y(n_265) );
BUFx10_ASAP7_75t_L g266 ( .A(n_187), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_197), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_226), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_177), .B(n_124), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_191), .B(n_122), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_177), .A2(n_122), .B1(n_108), .B2(n_107), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_177), .B(n_107), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_230), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_205), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_226), .Y(n_275) );
NOR2xp33_ASAP7_75t_R g276 ( .A(n_201), .B(n_165), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_201), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_226), .Y(n_278) );
NOR2xp33_ASAP7_75t_R g279 ( .A(n_208), .B(n_61), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_185), .B(n_2), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_191), .B(n_131), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_205), .Y(n_282) );
AO22x1_ASAP7_75t_L g283 ( .A1(n_226), .A2(n_89), .B1(n_4), .B2(n_5), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_232), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_232), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_180), .Y(n_286) );
NAND3xp33_ASAP7_75t_L g287 ( .A(n_186), .B(n_3), .C(n_5), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_206), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_185), .B(n_6), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_185), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_206), .Y(n_291) );
NOR2xp33_ASAP7_75t_SL g292 ( .A(n_179), .B(n_6), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_210), .B(n_7), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_183), .B(n_7), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_180), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_180), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_200), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_210), .B(n_8), .Y(n_298) );
NOR3xp33_ASAP7_75t_SL g299 ( .A(n_225), .B(n_8), .C(n_9), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_203), .Y(n_300) );
NOR2x1_ASAP7_75t_L g301 ( .A(n_200), .B(n_9), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_207), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_259), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_290), .B(n_200), .Y(n_304) );
CKINVDCx6p67_ASAP7_75t_R g305 ( .A(n_290), .Y(n_305) );
AOI21x1_ASAP7_75t_L g306 ( .A1(n_256), .A2(n_231), .B(n_224), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_252), .Y(n_307) );
AOI222xp33_ASAP7_75t_L g308 ( .A1(n_270), .A2(n_199), .B1(n_216), .B2(n_214), .C1(n_200), .C2(n_223), .Y(n_308) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_246), .B(n_216), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_246), .B(n_214), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_239), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_254), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_258), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_241), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_234), .B(n_224), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_261), .Y(n_316) );
INVx5_ASAP7_75t_L g317 ( .A(n_254), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_264), .Y(n_318) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_292), .A2(n_229), .B1(n_231), .B2(n_221), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_243), .B(n_219), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_251), .A2(n_196), .B(n_193), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_280), .B(n_219), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_254), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_252), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_254), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_255), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_265), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_254), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_280), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_257), .Y(n_330) );
NAND2x2_ASAP7_75t_L g331 ( .A(n_269), .B(n_218), .Y(n_331) );
INVx2_ASAP7_75t_SL g332 ( .A(n_293), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_293), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_297), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_277), .B(n_202), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_293), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_275), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_275), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_255), .Y(n_339) );
NAND2xp33_ASAP7_75t_L g340 ( .A(n_275), .B(n_193), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_270), .A2(n_227), .B1(n_215), .B2(n_207), .C(n_212), .Y(n_341) );
NOR2xp67_ASAP7_75t_SL g342 ( .A(n_275), .B(n_213), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_245), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_298), .B(n_213), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_236), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_277), .Y(n_346) );
BUFx8_ASAP7_75t_SL g347 ( .A(n_298), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_242), .B(n_215), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g349 ( .A1(n_298), .A2(n_176), .B1(n_178), .B2(n_212), .Y(n_349) );
CKINVDCx11_ASAP7_75t_R g350 ( .A(n_266), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_272), .B(n_211), .Y(n_351) );
INVx4_ASAP7_75t_L g352 ( .A(n_275), .Y(n_352) );
INVx4_ASAP7_75t_L g353 ( .A(n_264), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_274), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_270), .B(n_211), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_315), .A2(n_281), .B1(n_271), .B2(n_299), .C(n_253), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_354), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_333), .A2(n_289), .B1(n_294), .B2(n_262), .Y(n_358) );
BUFx3_ASAP7_75t_L g359 ( .A(n_317), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_SL g360 ( .A1(n_319), .A2(n_288), .B(n_274), .C(n_282), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_315), .B(n_282), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_307), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_331), .A2(n_281), .B1(n_301), .B2(n_266), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_304), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_331), .A2(n_281), .B1(n_266), .B2(n_238), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_307), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_355), .B(n_288), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_329), .A2(n_249), .B1(n_267), .B2(n_287), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_306), .A2(n_233), .B(n_217), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_324), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g371 ( .A1(n_332), .A2(n_302), .B1(n_291), .B2(n_235), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_347), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_308), .B(n_291), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_317), .Y(n_374) );
BUFx12f_ASAP7_75t_L g375 ( .A(n_350), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_324), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_322), .A2(n_267), .B1(n_249), .B2(n_247), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_326), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_322), .A2(n_249), .B1(n_267), .B2(n_302), .Y(n_379) );
INVx4_ASAP7_75t_L g380 ( .A(n_317), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g381 ( .A1(n_332), .A2(n_235), .B1(n_250), .B2(n_209), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_322), .A2(n_250), .B1(n_278), .B2(n_260), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_347), .A2(n_278), .B1(n_260), .B2(n_268), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_335), .A2(n_178), .B1(n_176), .B2(n_209), .C(n_198), .Y(n_384) );
AOI21xp33_ASAP7_75t_L g385 ( .A1(n_336), .A2(n_203), .B(n_198), .Y(n_385) );
INVx4_ASAP7_75t_L g386 ( .A(n_317), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_326), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_356), .A2(n_346), .B1(n_350), .B2(n_311), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_375), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_373), .A2(n_349), .B1(n_344), .B2(n_309), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_367), .B(n_344), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_370), .Y(n_392) );
AOI21xp33_ASAP7_75t_L g393 ( .A1(n_358), .A2(n_313), .B(n_343), .Y(n_393) );
AOI22xp33_ASAP7_75t_SL g394 ( .A1(n_372), .A2(n_345), .B1(n_346), .B2(n_314), .Y(n_394) );
OAI22xp33_ASAP7_75t_L g395 ( .A1(n_372), .A2(n_314), .B1(n_345), .B2(n_305), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_375), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_362), .Y(n_398) );
INVx4_ASAP7_75t_L g399 ( .A(n_380), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_380), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g401 ( .A1(n_361), .A2(n_321), .B(n_339), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_362), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_367), .B(n_361), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_L g404 ( .A1(n_358), .A2(n_309), .B(n_348), .C(n_355), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_356), .A2(n_330), .B1(n_320), .B2(n_341), .C(n_310), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_363), .A2(n_330), .B1(n_313), .B2(n_334), .C(n_303), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_373), .A2(n_305), .B1(n_310), .B2(n_351), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_366), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_357), .B(n_310), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_365), .B(n_304), .Y(n_410) );
INVxp67_ASAP7_75t_L g411 ( .A(n_384), .Y(n_411) );
OAI21x1_ASAP7_75t_L g412 ( .A1(n_369), .A2(n_339), .B(n_217), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_371), .A2(n_304), .B1(n_320), .B2(n_316), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_384), .A2(n_320), .B1(n_327), .B2(n_276), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_370), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_398), .Y(n_416) );
INVx4_ASAP7_75t_L g417 ( .A(n_399), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_398), .Y(n_418) );
OR2x6_ASAP7_75t_L g419 ( .A(n_413), .B(n_375), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_405), .A2(n_371), .B1(n_357), .B2(n_381), .Y(n_420) );
AND2x6_ASAP7_75t_SL g421 ( .A(n_389), .B(n_366), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_404), .A2(n_368), .B(n_381), .Y(n_422) );
NOR3xp33_ASAP7_75t_SL g423 ( .A(n_396), .B(n_385), .C(n_376), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_403), .B(n_364), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_409), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_402), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_413), .A2(n_364), .B1(n_379), .B2(n_382), .Y(n_427) );
BUFx3_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_403), .B(n_376), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_397), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_391), .B(n_378), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_390), .A2(n_378), .B1(n_387), .B2(n_377), .Y(n_432) );
INVx5_ASAP7_75t_SL g433 ( .A(n_409), .Y(n_433) );
INVx11_ASAP7_75t_L g434 ( .A(n_394), .Y(n_434) );
INVxp67_ASAP7_75t_L g435 ( .A(n_409), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_402), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_408), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_388), .B(n_197), .C(n_198), .D(n_385), .Y(n_438) );
BUFx4f_ASAP7_75t_L g439 ( .A(n_409), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_391), .B(n_387), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_406), .A2(n_383), .B1(n_360), .B2(n_176), .C(n_178), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_411), .A2(n_283), .B1(n_387), .B2(n_380), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_392), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_399), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_408), .B(n_197), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_392), .Y(n_446) );
OAI33xp33_ASAP7_75t_L g447 ( .A1(n_395), .A2(n_194), .A3(n_196), .B1(n_233), .B2(n_217), .B3(n_248), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_400), .Y(n_448) );
NOR2xp33_ASAP7_75t_R g449 ( .A(n_400), .B(n_359), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_410), .B(n_283), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_407), .A2(n_386), .B1(n_380), .B2(n_374), .Y(n_451) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_412), .A2(n_369), .B(n_233), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_443), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_416), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_431), .B(n_392), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_428), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_429), .B(n_415), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_418), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_426), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_443), .B(n_415), .Y(n_460) );
OAI33xp33_ASAP7_75t_L g461 ( .A1(n_436), .A2(n_390), .A3(n_194), .B1(n_12), .B2(n_13), .B3(n_14), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_428), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_437), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_446), .Y(n_464) );
INVx4_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_452), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_449), .Y(n_467) );
OAI21xp33_ASAP7_75t_L g468 ( .A1(n_419), .A2(n_393), .B(n_414), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_430), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_440), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_430), .B(n_415), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_419), .B(n_400), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_452), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_419), .A2(n_399), .B1(n_400), .B2(n_401), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_424), .B(n_399), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_448), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_448), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_432), .B(n_401), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_423), .B(n_386), .C(n_203), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_432), .B(n_412), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_417), .B(n_374), .Y(n_481) );
OAI33xp33_ASAP7_75t_L g482 ( .A1(n_427), .A2(n_10), .A3(n_11), .B1(n_12), .B2(n_15), .B3(n_16), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_450), .A2(n_386), .B1(n_374), .B2(n_359), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_417), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_445), .B(n_359), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_433), .B(n_198), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_425), .Y(n_487) );
AOI221xp5_ASAP7_75t_SL g488 ( .A1(n_435), .A2(n_176), .B1(n_178), .B2(n_244), .C(n_237), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_444), .Y(n_489) );
NOR2x1_ASAP7_75t_L g490 ( .A(n_438), .B(n_386), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_449), .Y(n_491) );
NOR2x1_ASAP7_75t_L g492 ( .A(n_441), .B(n_352), .Y(n_492) );
AOI33xp33_ASAP7_75t_L g493 ( .A1(n_420), .A2(n_11), .A3(n_15), .B1(n_16), .B2(n_17), .B3(n_18), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_451), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_421), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_442), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_439), .B(n_420), .Y(n_497) );
NAND2x1p5_ASAP7_75t_L g498 ( .A(n_439), .B(n_317), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_433), .B(n_17), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_444), .B(n_18), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_433), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_450), .B(n_19), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_423), .Y(n_503) );
NAND4xp25_ASAP7_75t_L g504 ( .A(n_422), .B(n_203), .C(n_20), .D(n_21), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_434), .B(n_19), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_447), .B(n_369), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_416), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_454), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_454), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_475), .B(n_22), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_502), .B(n_504), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_458), .Y(n_512) );
NOR2x1_ASAP7_75t_L g513 ( .A(n_465), .B(n_352), .Y(n_513) );
OAI22xp33_ASAP7_75t_L g514 ( .A1(n_504), .A2(n_352), .B1(n_328), .B2(n_353), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_475), .B(n_25), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_458), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_459), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_470), .B(n_29), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_459), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_500), .B(n_31), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_469), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_456), .B(n_240), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_465), .B(n_279), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_463), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_465), .B(n_338), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_495), .B(n_36), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_462), .B(n_240), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_507), .B(n_237), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_455), .B(n_244), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_457), .B(n_248), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_453), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_453), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_499), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_453), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_463), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_507), .Y(n_536) );
AND4x1_ASAP7_75t_L g537 ( .A(n_505), .B(n_342), .C(n_40), .D(n_46), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_471), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_490), .A2(n_338), .B(n_337), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_471), .B(n_39), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_497), .B(n_48), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_485), .B(n_51), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_464), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_481), .Y(n_544) );
NAND2xp33_ASAP7_75t_R g545 ( .A(n_491), .B(n_53), .Y(n_545) );
NOR3xp33_ASAP7_75t_L g546 ( .A(n_482), .B(n_180), .C(n_189), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_497), .B(n_54), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_464), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_460), .B(n_55), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_460), .B(n_56), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_464), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_496), .B(n_57), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_484), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_465), .B(n_328), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_484), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_496), .B(n_189), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_489), .B(n_189), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_489), .B(n_189), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_499), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_468), .B(n_190), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_485), .B(n_328), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_472), .B(n_190), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_478), .B(n_190), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_478), .B(n_190), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_461), .A2(n_263), .B1(n_285), .B2(n_273), .C(n_284), .Y(n_565) );
AOI31xp33_ASAP7_75t_L g566 ( .A1(n_467), .A2(n_353), .A3(n_325), .B(n_323), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_473), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_481), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_472), .B(n_300), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_477), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_487), .B(n_300), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_476), .Y(n_572) );
OAI31xp33_ASAP7_75t_L g573 ( .A1(n_514), .A2(n_468), .A3(n_467), .B(n_503), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_521), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_544), .B(n_477), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_532), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_538), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_521), .Y(n_578) );
AOI321xp33_ASAP7_75t_L g579 ( .A1(n_511), .A2(n_490), .A3(n_503), .B1(n_474), .B2(n_491), .C(n_494), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_538), .B(n_494), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_508), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_568), .B(n_533), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_532), .Y(n_583) );
AO21x1_ASAP7_75t_L g584 ( .A1(n_514), .A2(n_476), .B(n_506), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_509), .Y(n_585) );
AOI21xp33_ASAP7_75t_L g586 ( .A1(n_511), .A2(n_488), .B(n_501), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_545), .A2(n_494), .B1(n_501), .B2(n_487), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_512), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_523), .A2(n_493), .B(n_492), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_516), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_517), .B(n_480), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_559), .B(n_480), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_526), .A2(n_473), .B1(n_466), .B2(n_483), .C(n_479), .Y(n_593) );
AOI21xp33_ASAP7_75t_SL g594 ( .A1(n_545), .A2(n_498), .B(n_483), .Y(n_594) );
INVxp33_ASAP7_75t_L g595 ( .A(n_526), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_519), .B(n_473), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_546), .A2(n_492), .B1(n_506), .B2(n_466), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_567), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_553), .B(n_486), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_523), .A2(n_479), .B(n_486), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_524), .B(n_498), .Y(n_601) );
NOR2xp67_ASAP7_75t_L g602 ( .A(n_525), .B(n_498), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_535), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g604 ( .A1(n_520), .A2(n_312), .B(n_323), .C(n_325), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_536), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_555), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g607 ( .A1(n_552), .A2(n_340), .B(n_318), .C(n_273), .Y(n_607) );
AOI221x1_ASAP7_75t_L g608 ( .A1(n_560), .A2(n_353), .B1(n_338), .B2(n_337), .C(n_318), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_572), .B(n_263), .Y(n_609) );
INVx2_ASAP7_75t_SL g610 ( .A(n_554), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_548), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_541), .B(n_547), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_520), .B(n_318), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_543), .B(n_300), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_551), .B(n_284), .Y(n_615) );
AOI322xp5_ASAP7_75t_L g616 ( .A1(n_510), .A2(n_340), .A3(n_268), .B1(n_312), .B2(n_285), .C1(n_337), .C2(n_338), .Y(n_616) );
NOR2x1_ASAP7_75t_L g617 ( .A(n_513), .B(n_337), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_543), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_561), .A2(n_337), .B1(n_338), .B2(n_300), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_570), .B(n_300), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_540), .A2(n_286), .B1(n_295), .B2(n_296), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_563), .B(n_295), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_567), .Y(n_623) );
OAI21xp5_ASAP7_75t_SL g624 ( .A1(n_566), .A2(n_296), .B(n_537), .Y(n_624) );
AOI221x1_ASAP7_75t_L g625 ( .A1(n_560), .A2(n_546), .B1(n_564), .B2(n_556), .C(n_558), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_554), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_525), .A2(n_539), .B(n_515), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_531), .B(n_534), .Y(n_628) );
OAI211xp5_ASAP7_75t_SL g629 ( .A1(n_562), .A2(n_550), .B(n_549), .C(n_569), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_534), .B(n_530), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_610), .Y(n_631) );
NAND2xp33_ASAP7_75t_SL g632 ( .A(n_626), .B(n_542), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_574), .B(n_571), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_576), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_576), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_618), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_583), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_606), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_592), .B(n_518), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_581), .Y(n_640) );
INVxp33_ASAP7_75t_L g641 ( .A(n_594), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_582), .B(n_522), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_585), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_588), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_595), .B(n_586), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_590), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_587), .B(n_527), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_578), .B(n_529), .Y(n_648) );
INVx2_ASAP7_75t_SL g649 ( .A(n_577), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_611), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_575), .B(n_557), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_603), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_591), .B(n_528), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_628), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_612), .B(n_565), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_598), .B(n_623), .Y(n_656) );
INVx3_ASAP7_75t_L g657 ( .A(n_605), .Y(n_657) );
INVxp67_ASAP7_75t_SL g658 ( .A(n_598), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_580), .B(n_630), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_624), .A2(n_573), .B(n_593), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_623), .B(n_599), .Y(n_661) );
NOR2xp33_ASAP7_75t_SL g662 ( .A(n_602), .B(n_627), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_596), .B(n_601), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_614), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_584), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_609), .Y(n_666) );
XNOR2x2_ASAP7_75t_L g667 ( .A(n_593), .B(n_627), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_597), .B(n_625), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_597), .B(n_612), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_615), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_620), .B(n_589), .Y(n_671) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_660), .B(n_629), .C(n_600), .Y(n_672) );
INVxp67_ASAP7_75t_L g673 ( .A(n_645), .Y(n_673) );
INVx1_ASAP7_75t_SL g674 ( .A(n_631), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_655), .A2(n_629), .B1(n_613), .B2(n_622), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_663), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_656), .B(n_669), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_641), .B(n_621), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_663), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_671), .Y(n_680) );
NOR2xp33_ASAP7_75t_SL g681 ( .A(n_662), .B(n_617), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_656), .B(n_619), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_660), .A2(n_607), .B(n_604), .C(n_579), .Y(n_683) );
NAND2xp33_ASAP7_75t_SL g684 ( .A(n_665), .B(n_608), .Y(n_684) );
XOR2xp5_ASAP7_75t_L g685 ( .A(n_667), .B(n_616), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_638), .Y(n_686) );
AOI21xp5_ASAP7_75t_SL g687 ( .A1(n_668), .A2(n_607), .B(n_667), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_657), .A2(n_642), .B1(n_647), .B2(n_658), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_653), .B(n_661), .Y(n_689) );
NOR2xp67_ASAP7_75t_L g690 ( .A(n_657), .B(n_635), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_638), .Y(n_691) );
XOR2xp5_ASAP7_75t_L g692 ( .A(n_651), .B(n_639), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_634), .B(n_632), .C(n_635), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_673), .B(n_659), .Y(n_694) );
AOI222xp33_ASAP7_75t_L g695 ( .A1(n_680), .A2(n_661), .B1(n_639), .B2(n_648), .C1(n_651), .C2(n_666), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_676), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_672), .A2(n_646), .B1(n_644), .B2(n_643), .C(n_652), .Y(n_697) );
OAI221xp5_ASAP7_75t_SL g698 ( .A1(n_685), .A2(n_642), .B1(n_633), .B2(n_666), .C(n_664), .Y(n_698) );
NAND2xp33_ASAP7_75t_SL g699 ( .A(n_688), .B(n_649), .Y(n_699) );
NAND2x1p5_ASAP7_75t_L g700 ( .A(n_690), .B(n_649), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g701 ( .A(n_674), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_678), .A2(n_646), .B1(n_652), .B2(n_640), .Y(n_702) );
CKINVDCx16_ASAP7_75t_R g703 ( .A(n_681), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_692), .Y(n_704) );
NOR2xp33_ASAP7_75t_R g705 ( .A(n_678), .B(n_670), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_679), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_677), .B(n_644), .Y(n_707) );
AND4x1_ASAP7_75t_L g708 ( .A(n_687), .B(n_640), .C(n_643), .D(n_670), .Y(n_708) );
XNOR2xp5_ASAP7_75t_L g709 ( .A(n_693), .B(n_664), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_683), .A2(n_650), .B(n_654), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_684), .A2(n_636), .B(n_637), .Y(n_711) );
OAI211xp5_ASAP7_75t_L g712 ( .A1(n_675), .A2(n_636), .B(n_637), .C(n_684), .Y(n_712) );
INVx2_ASAP7_75t_SL g713 ( .A(n_689), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_682), .B(n_686), .C(n_691), .Y(n_714) );
OAI321xp33_ASAP7_75t_L g715 ( .A1(n_675), .A2(n_683), .A3(n_665), .B1(n_668), .B2(n_688), .C(n_673), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_701), .Y(n_716) );
XNOR2xp5_ASAP7_75t_L g717 ( .A(n_704), .B(n_708), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_703), .A2(n_698), .B1(n_700), .B2(n_710), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g719 ( .A(n_705), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_697), .B(n_714), .Y(n_720) );
OAI211xp5_ASAP7_75t_SL g721 ( .A1(n_718), .A2(n_712), .B(n_715), .C(n_695), .Y(n_721) );
NAND3xp33_ASAP7_75t_SL g722 ( .A(n_719), .B(n_699), .C(n_711), .Y(n_722) );
NOR3xp33_ASAP7_75t_L g723 ( .A(n_720), .B(n_715), .C(n_694), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_722), .Y(n_724) );
AOI211xp5_ASAP7_75t_L g725 ( .A1(n_721), .A2(n_717), .B(n_716), .C(n_709), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_724), .Y(n_726) );
OR2x2_ASAP7_75t_L g727 ( .A(n_725), .B(n_723), .Y(n_727) );
AOI322xp5_ASAP7_75t_L g728 ( .A1(n_726), .A2(n_716), .A3(n_702), .B1(n_713), .B2(n_696), .C1(n_706), .C2(n_707), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_728), .A2(n_727), .B(n_700), .Y(n_729) );
endmodule