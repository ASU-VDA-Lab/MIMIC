module fake_jpeg_7426_n_210 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_210);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_26),
.Y(n_44)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_27),
.A2(n_17),
.B1(n_15),
.B2(n_22),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_32),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_48),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_23),
.B1(n_17),
.B2(n_22),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_46),
.B1(n_50),
.B2(n_26),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_27),
.A2(n_23),
.B1(n_17),
.B2(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_15),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_26),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_25),
.B1(n_24),
.B2(n_15),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_19),
.B1(n_21),
.B2(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_64),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_59),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_29),
.B(n_20),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_63),
.B1(n_67),
.B2(n_36),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_39),
.B1(n_33),
.B2(n_31),
.Y(n_85)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_45),
.Y(n_71)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_75),
.B(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_72),
.Y(n_100)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_12),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_73),
.Y(n_98)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_58),
.B(n_16),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_39),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_68),
.B1(n_72),
.B2(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_16),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_57),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_89),
.C(n_59),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_63),
.B1(n_56),
.B2(n_65),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_35),
.B1(n_30),
.B2(n_47),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_53),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_91),
.B1(n_80),
.B2(n_47),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_95),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_96),
.B(n_85),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_64),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_58),
.B(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_59),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_59),
.B(n_78),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_103),
.B(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_73),
.B1(n_75),
.B2(n_78),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_97),
.B1(n_91),
.B2(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_114),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_121),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_116),
.B(n_117),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_69),
.B(n_66),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_70),
.B(n_47),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_120),
.B1(n_94),
.B2(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_95),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_111),
.B1(n_120),
.B2(n_109),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_126),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_128),
.Y(n_153)
);

NAND2x1_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_87),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_98),
.B1(n_99),
.B2(n_97),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_104),
.B1(n_35),
.B2(n_70),
.Y(n_154)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_89),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_104),
.B(n_70),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_145),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_116),
.B1(n_112),
.B2(n_119),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_114),
.C(n_107),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_151),
.C(n_126),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_117),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_35),
.B1(n_0),
.B2(n_2),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_155),
.A2(n_128),
.B1(n_123),
.B2(n_136),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_161),
.C(n_162),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_163),
.B1(n_166),
.B2(n_155),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_149),
.A2(n_124),
.B(n_135),
.C(n_137),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_158),
.A2(n_0),
.B1(n_35),
.B2(n_2),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_168),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_151),
.C(n_152),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_129),
.C(n_134),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_129),
.B(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_147),
.B(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_140),
.B1(n_123),
.B2(n_126),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_159),
.B(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_175),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_SL g184 ( 
.A1(n_173),
.A2(n_176),
.B(n_158),
.C(n_4),
.Y(n_184)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_1),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_2),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_168),
.B(n_1),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_3),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_165),
.B(n_158),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_181),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_185),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_184),
.A2(n_170),
.B1(n_176),
.B2(n_183),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_172),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_188),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_70),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_189),
.A2(n_193),
.B1(n_4),
.B2(n_7),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_7),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_177),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_192),
.B(n_189),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_177),
.C(n_6),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_198),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_11),
.C(n_6),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

AOI322xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_201),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_185),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_191),
.B(n_8),
.C(n_9),
.Y(n_202)
);

FAx1_ASAP7_75t_SL g201 ( 
.A(n_195),
.B(n_11),
.CI(n_8),
.CON(n_201),
.SN(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_202),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_201),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_205),
.B(n_203),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_207),
.C(n_9),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_10),
.Y(n_210)
);


endmodule