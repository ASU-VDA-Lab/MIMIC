module fake_netlist_6_1383_n_1735 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1735);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1735;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_40),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_109),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_129),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_76),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_100),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_38),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_21),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_18),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_11),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_42),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_40),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_5),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_147),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_18),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_39),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_106),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_126),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_52),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_3),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_37),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_94),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_24),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_52),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_139),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_9),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_101),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_8),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_25),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_35),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_51),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_96),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_62),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_55),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_29),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_103),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_30),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_43),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_32),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_44),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_87),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_128),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_16),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_7),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_61),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_59),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_118),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_127),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_91),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_78),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_112),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_119),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_65),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_20),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_57),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_35),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_29),
.Y(n_220)
);

CKINVDCx11_ASAP7_75t_R g221 ( 
.A(n_27),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_50),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_110),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_71),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_70),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_136),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_46),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_154),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_84),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_42),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_28),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_145),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_24),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_124),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_108),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_62),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_80),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_138),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_20),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_43),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_11),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_143),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_65),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_57),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_53),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_13),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_85),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_54),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_131),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_54),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_149),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_10),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_6),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_15),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_153),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_19),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_98),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_68),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_13),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_36),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_46),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_4),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_64),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_104),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_92),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_81),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_82),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_90),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_107),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_150),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_75),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_148),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_99),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_8),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_58),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_12),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_72),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_67),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_102),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_48),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_64),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_59),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_68),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_7),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_16),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_15),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_4),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_67),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_30),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_33),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_38),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_61),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_3),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_141),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_120),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_21),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_23),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_60),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_63),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_44),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_51),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_45),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_83),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_117),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_105),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_36),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_1),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_151),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_27),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_240),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_221),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_158),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_240),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_240),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_160),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_240),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_240),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_243),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_167),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_161),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_262),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_167),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_168),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_262),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_188),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_202),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_262),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_173),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_262),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_283),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_202),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_214),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_175),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_283),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_178),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_202),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_192),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_183),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_192),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_186),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_245),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_250),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_291),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_248),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_288),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_248),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_248),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_287),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_287),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_193),
.Y(n_358)
);

BUFx2_ASAP7_75t_SL g359 ( 
.A(n_159),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_187),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_279),
.B(n_0),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_196),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_198),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_210),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_287),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_212),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_214),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_299),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_234),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_299),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_299),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g372 ( 
.A(n_302),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_218),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_190),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_156),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_218),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_218),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_226),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_166),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_190),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_228),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_166),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_232),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_169),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_169),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_324),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_310),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_337),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_310),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_279),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_187),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_337),
.Y(n_395)
);

INVx5_ASAP7_75t_L g396 ( 
.A(n_337),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_207),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_314),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_346),
.B(n_224),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_329),
.B(n_234),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_315),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_329),
.B(n_336),
.Y(n_403)
);

OA21x2_ASAP7_75t_L g404 ( 
.A1(n_367),
.A2(n_181),
.B(n_171),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_317),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_336),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_352),
.B(n_200),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_320),
.A2(n_307),
.B1(n_256),
.B2(n_200),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_318),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_318),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_322),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_367),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_367),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_322),
.B(n_224),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_323),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_326),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_328),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_328),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_369),
.B(n_159),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_330),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_324),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_361),
.B(n_181),
.C(n_171),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_330),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_361),
.B(n_224),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_369),
.B(n_163),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_165),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_332),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_372),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_332),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_333),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_371),
.B(n_234),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_333),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_319),
.A2(n_256),
.B1(n_301),
.B2(n_189),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_334),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_334),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_335),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_335),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_339),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_339),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_376),
.B(n_294),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_340),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_359),
.B(n_237),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_340),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_341),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_341),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_343),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_376),
.B(n_242),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_343),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_379),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_391),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_446),
.B(n_375),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_404),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_403),
.B(n_312),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_408),
.B(n_316),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_403),
.B(n_321),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_404),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_403),
.B(n_325),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_407),
.B(n_331),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_416),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_408),
.B(n_338),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_342),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_436),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_407),
.B(n_345),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_432),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_415),
.B(n_294),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_404),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_436),
.Y(n_477)
);

BUFx4f_ASAP7_75t_L g478 ( 
.A(n_404),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_413),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_409),
.B(n_327),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_399),
.B(n_347),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_420),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_413),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_447),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_432),
.B(n_358),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_413),
.Y(n_486)
);

INVx5_ASAP7_75t_L g487 ( 
.A(n_413),
.Y(n_487)
);

NAND3xp33_ASAP7_75t_SL g488 ( 
.A(n_409),
.B(n_348),
.C(n_319),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_391),
.B(n_401),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_447),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_401),
.B(n_377),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_413),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_401),
.B(n_362),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_447),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_447),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_387),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_386),
.B(n_320),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_436),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_432),
.B(n_363),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_387),
.Y(n_500)
);

BUFx8_ASAP7_75t_SL g501 ( 
.A(n_429),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_436),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_389),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_427),
.A2(n_354),
.B1(n_344),
.B2(n_217),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_435),
.B(n_377),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_L g506 ( 
.A(n_429),
.B(n_364),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_389),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_399),
.B(n_366),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_452),
.B(n_378),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_422),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_438),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_428),
.B(n_381),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_428),
.B(n_383),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_413),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_435),
.B(n_179),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_413),
.Y(n_518)
);

AO22x2_ASAP7_75t_L g519 ( 
.A1(n_427),
.A2(n_354),
.B1(n_217),
.B2(n_207),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_435),
.B(n_179),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_386),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_422),
.B(n_204),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_SL g523 ( 
.A(n_424),
.B(n_311),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_438),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_424),
.B(n_374),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_444),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_438),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_441),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_413),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_437),
.B(n_348),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_441),
.Y(n_531)
);

BUFx8_ASAP7_75t_SL g532 ( 
.A(n_444),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_392),
.Y(n_533)
);

OR2x6_ASAP7_75t_L g534 ( 
.A(n_425),
.B(n_294),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_425),
.B(n_238),
.Y(n_535)
);

INVx4_ASAP7_75t_SL g536 ( 
.A(n_415),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_444),
.A2(n_224),
.B1(n_227),
.B2(n_254),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_441),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_430),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_430),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_415),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_441),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_397),
.B(n_255),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_393),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_397),
.B(n_360),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_437),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_415),
.A2(n_233),
.B1(n_254),
.B2(n_246),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_393),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_415),
.A2(n_189),
.B1(n_194),
.B2(n_206),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_397),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_450),
.B(n_269),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_414),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_414),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_431),
.B(n_204),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_431),
.B(n_360),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_415),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_450),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_398),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_431),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_394),
.A2(n_194),
.B1(n_206),
.B2(n_209),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_R g561 ( 
.A(n_454),
.B(n_162),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_454),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_431),
.B(n_157),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_414),
.Y(n_564)
);

NAND3xp33_ASAP7_75t_L g565 ( 
.A(n_394),
.B(n_295),
.C(n_214),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_451),
.B(n_351),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_414),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_431),
.B(n_374),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_398),
.Y(n_569)
);

NOR2x1p5_ASAP7_75t_L g570 ( 
.A(n_451),
.B(n_197),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_400),
.B(n_205),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_400),
.A2(n_272),
.B1(n_222),
.B2(n_220),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_417),
.B(n_380),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_451),
.B(n_295),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_417),
.B(n_418),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_414),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_418),
.B(n_205),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_419),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_419),
.B(n_421),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_453),
.B(n_247),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_442),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_420),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_421),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_423),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_453),
.A2(n_209),
.B1(n_216),
.B2(n_219),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_423),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_433),
.B(n_211),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_433),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_434),
.B(n_380),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_420),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_453),
.B(n_295),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_434),
.B(n_211),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_445),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_445),
.B(n_213),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_449),
.A2(n_216),
.B1(n_219),
.B2(n_227),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_414),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_449),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_420),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_390),
.A2(n_301),
.B1(n_260),
.B2(n_259),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_390),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_442),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_390),
.B(n_213),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_402),
.B(n_223),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_550),
.B(n_349),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_511),
.B(n_489),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_541),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_510),
.B(n_402),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_478),
.B(n_556),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_539),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_457),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_457),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_470),
.B(n_402),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_478),
.B(n_164),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_466),
.B(n_405),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_550),
.B(n_349),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_534),
.A2(n_157),
.B1(n_270),
.B2(n_170),
.Y(n_616)
);

AND2x2_ASAP7_75t_SL g617 ( 
.A(n_481),
.B(n_164),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_497),
.B(n_382),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_459),
.A2(n_274),
.B(n_246),
.C(n_239),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_539),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_478),
.B(n_164),
.Y(n_621)
);

NOR2x1p5_ASAP7_75t_L g622 ( 
.A(n_488),
.B(n_172),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_556),
.B(n_526),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_459),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_458),
.B(n_463),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_472),
.B(n_405),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_545),
.Y(n_627)
);

NOR2xp67_ASAP7_75t_L g628 ( 
.A(n_456),
.B(n_249),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_L g629 ( 
.A(n_464),
.B(n_164),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_465),
.A2(n_264),
.B1(n_235),
.B2(n_271),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_526),
.B(n_405),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_493),
.B(n_406),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_539),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_578),
.B(n_406),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_516),
.B(n_223),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_541),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_578),
.B(n_406),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_520),
.A2(n_229),
.B1(n_277),
.B2(n_225),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_586),
.B(n_410),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_506),
.A2(n_229),
.B1(n_277),
.B2(n_257),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_586),
.B(n_410),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_491),
.B(n_410),
.Y(n_642)
);

NAND3xp33_ASAP7_75t_L g643 ( 
.A(n_504),
.B(n_176),
.C(n_174),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_491),
.B(n_411),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_464),
.B(n_475),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_455),
.B(n_164),
.Y(n_646)
);

INVx8_ASAP7_75t_L g647 ( 
.A(n_574),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_534),
.A2(n_225),
.B1(n_170),
.B2(n_201),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_475),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_455),
.B(n_164),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_484),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_484),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_497),
.B(n_382),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_521),
.B(n_505),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_455),
.B(n_251),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_505),
.B(n_411),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_522),
.B(n_411),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_476),
.A2(n_233),
.B(n_239),
.C(n_261),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_476),
.B(n_251),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_496),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_R g661 ( 
.A(n_473),
.B(n_350),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_496),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_490),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_501),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_557),
.B(n_177),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_490),
.Y(n_666)
);

AO221x1_ASAP7_75t_L g667 ( 
.A1(n_519),
.A2(n_251),
.B1(n_261),
.B2(n_274),
.C(n_276),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_535),
.A2(n_305),
.B1(n_303),
.B2(n_308),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_521),
.B(n_350),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_559),
.B(n_600),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_559),
.B(n_600),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_557),
.B(n_251),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_561),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_525),
.Y(n_674)
);

AOI222xp33_ASAP7_75t_L g675 ( 
.A1(n_546),
.A2(n_276),
.B1(n_281),
.B2(n_282),
.C1(n_292),
.C2(n_185),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_474),
.Y(n_676)
);

AO221x1_ASAP7_75t_L g677 ( 
.A1(n_519),
.A2(n_572),
.B1(n_251),
.B2(n_281),
.C(n_282),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_525),
.Y(n_678)
);

AND2x6_ASAP7_75t_SL g679 ( 
.A(n_534),
.B(n_292),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_570),
.B(n_201),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_494),
.B(n_412),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_494),
.B(n_412),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_495),
.B(n_474),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_495),
.B(n_440),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_500),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_474),
.B(n_440),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_562),
.B(n_536),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_562),
.B(n_251),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_474),
.B(n_440),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_500),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_573),
.B(n_384),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_503),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_603),
.B(n_215),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_534),
.B(n_215),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_503),
.B(n_235),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_568),
.A2(n_264),
.B1(n_267),
.B2(n_270),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_540),
.Y(n_697)
);

AND2x6_ASAP7_75t_SL g698 ( 
.A(n_530),
.B(n_384),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_507),
.B(n_267),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_507),
.B(n_271),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_517),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_517),
.B(n_304),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_513),
.B(n_180),
.Y(n_703)
);

NAND2x1p5_ASAP7_75t_L g704 ( 
.A(n_563),
.B(n_304),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_533),
.B(n_420),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_514),
.B(n_182),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_533),
.B(n_420),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_568),
.B(n_385),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_544),
.B(n_420),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_589),
.B(n_290),
.C(n_191),
.Y(n_710)
);

BUFx6f_ASAP7_75t_SL g711 ( 
.A(n_540),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_583),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_544),
.B(n_420),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_548),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_548),
.B(n_426),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_558),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_558),
.B(n_426),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_569),
.Y(n_718)
);

INVx8_ASAP7_75t_L g719 ( 
.A(n_574),
.Y(n_719)
);

AND2x6_ASAP7_75t_SL g720 ( 
.A(n_530),
.B(n_385),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_569),
.B(n_426),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_536),
.B(n_265),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_536),
.B(n_266),
.Y(n_723)
);

O2A1O1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_602),
.A2(n_357),
.B(n_370),
.C(n_368),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_584),
.B(n_426),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_584),
.B(n_426),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_588),
.B(n_426),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_588),
.B(n_426),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_536),
.B(n_351),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_L g730 ( 
.A(n_565),
.B(n_268),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_515),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_593),
.B(n_426),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_593),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_597),
.B(n_439),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_597),
.Y(n_735)
);

OAI21xp33_ASAP7_75t_L g736 ( 
.A1(n_599),
.A2(n_289),
.B(n_195),
.Y(n_736)
);

AOI221xp5_ASAP7_75t_L g737 ( 
.A1(n_546),
.A2(n_519),
.B1(n_480),
.B2(n_543),
.C(n_599),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_594),
.B(n_439),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_509),
.A2(n_273),
.B1(n_184),
.B2(n_286),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_461),
.B(n_353),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_554),
.B(n_439),
.Y(n_741)
);

AO221x1_ASAP7_75t_L g742 ( 
.A1(n_519),
.A2(n_365),
.B1(n_355),
.B2(n_356),
.C(n_370),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_555),
.B(n_439),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_566),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_571),
.A2(n_296),
.B1(n_203),
.B2(n_208),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_563),
.B(n_414),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_563),
.B(n_439),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_563),
.A2(n_443),
.B1(n_442),
.B2(n_388),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_551),
.B(n_199),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_583),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_468),
.A2(n_298),
.B1(n_231),
.B2(n_236),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_R g752 ( 
.A(n_473),
.B(n_230),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_575),
.B(n_439),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_579),
.B(n_439),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_583),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_577),
.B(n_587),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_592),
.B(n_414),
.Y(n_757)
);

INVx8_ASAP7_75t_L g758 ( 
.A(n_532),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_515),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_537),
.A2(n_306),
.B1(n_244),
.B2(n_252),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_480),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_566),
.B(n_479),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_L g763 ( 
.A(n_515),
.B(n_241),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_460),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_479),
.B(n_439),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_574),
.A2(n_443),
.B1(n_442),
.B2(n_388),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_460),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_580),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_479),
.B(n_448),
.Y(n_769)
);

NOR2x1p5_ASAP7_75t_L g770 ( 
.A(n_565),
.B(n_253),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_483),
.B(n_448),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_483),
.B(n_448),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_L g773 ( 
.A(n_547),
.B(n_309),
.C(n_263),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_483),
.B(n_448),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_629),
.A2(n_482),
.B(n_598),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_629),
.A2(n_482),
.B(n_598),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_660),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_744),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_625),
.B(n_549),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_676),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_617),
.A2(n_574),
.B1(n_591),
.B2(n_499),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_SL g782 ( 
.A1(n_619),
.A2(n_601),
.B(n_462),
.C(n_581),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_676),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_654),
.B(n_485),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_741),
.A2(n_590),
.B(n_598),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_625),
.B(n_605),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_744),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_613),
.A2(n_590),
.B(n_482),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_617),
.A2(n_574),
.B1(n_591),
.B2(n_523),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_669),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_R g791 ( 
.A(n_712),
.B(n_258),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_613),
.A2(n_590),
.B(n_582),
.Y(n_792)
);

INVx11_ASAP7_75t_L g793 ( 
.A(n_711),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_627),
.B(n_591),
.Y(n_794)
);

AOI21x1_ASAP7_75t_L g795 ( 
.A1(n_621),
.A2(n_601),
.B(n_462),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_660),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_621),
.A2(n_582),
.B(n_515),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_759),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_608),
.A2(n_731),
.B(n_762),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_662),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_610),
.B(n_486),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_662),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_610),
.B(n_486),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_SL g804 ( 
.A(n_675),
.B(n_560),
.C(n_585),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_670),
.Y(n_805)
);

NOR3xp33_ASAP7_75t_L g806 ( 
.A(n_737),
.B(n_293),
.C(n_278),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_729),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_692),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_608),
.A2(n_582),
.B(n_515),
.Y(n_809)
);

NOR2xp67_ASAP7_75t_L g810 ( 
.A(n_664),
.B(n_595),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_607),
.A2(n_591),
.B1(n_492),
.B2(n_529),
.Y(n_811)
);

AOI211xp5_ASAP7_75t_L g812 ( 
.A1(n_749),
.A2(n_300),
.B(n_280),
.C(n_284),
.Y(n_812)
);

NAND2xp33_ASAP7_75t_L g813 ( 
.A(n_647),
.B(n_518),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_731),
.A2(n_683),
.B(n_645),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_731),
.A2(n_645),
.B(n_671),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_747),
.A2(n_596),
.B(n_518),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_659),
.A2(n_492),
.B(n_529),
.Y(n_817)
);

NOR2x1p5_ASAP7_75t_L g818 ( 
.A(n_712),
.B(n_275),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_756),
.A2(n_591),
.B1(n_492),
.B2(n_529),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_635),
.B(n_564),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_674),
.B(n_285),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_753),
.A2(n_553),
.B(n_552),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_635),
.B(n_564),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_612),
.B(n_564),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_692),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_614),
.B(n_567),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_659),
.A2(n_567),
.B(n_581),
.Y(n_827)
);

OR2x6_ASAP7_75t_L g828 ( 
.A(n_758),
.B(n_353),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_626),
.B(n_632),
.Y(n_829)
);

AND2x6_ASAP7_75t_L g830 ( 
.A(n_611),
.B(n_518),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_754),
.A2(n_576),
.B(n_553),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_611),
.B(n_518),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_686),
.A2(n_576),
.B(n_553),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_674),
.B(n_297),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_624),
.B(n_518),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_606),
.B(n_636),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_689),
.A2(n_576),
.B(n_553),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_624),
.B(n_552),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_743),
.A2(n_524),
.B(n_469),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_746),
.A2(n_576),
.B(n_553),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_746),
.A2(n_596),
.B(n_576),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_678),
.B(n_467),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_623),
.A2(n_552),
.B(n_596),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_623),
.A2(n_552),
.B(n_596),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_649),
.A2(n_687),
.B1(n_690),
.B2(n_685),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_649),
.A2(n_477),
.B1(n_467),
.B2(n_542),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_693),
.A2(n_355),
.B(n_356),
.C(n_357),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_729),
.B(n_552),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_729),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_657),
.B(n_469),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_718),
.B(n_596),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_759),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_738),
.A2(n_487),
.B(n_388),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_759),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_691),
.B(n_471),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_665),
.B(n_471),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_757),
.A2(n_487),
.B(n_395),
.Y(n_857)
);

AOI21xp33_ASAP7_75t_L g858 ( 
.A1(n_749),
.A2(n_0),
.B(n_1),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_718),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_733),
.Y(n_860)
);

NOR2xp67_ASAP7_75t_L g861 ( 
.A(n_750),
.B(n_69),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_701),
.B(n_477),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_619),
.A2(n_542),
.B(n_538),
.C(n_531),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_714),
.B(n_498),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_658),
.A2(n_538),
.B(n_531),
.C(n_528),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_716),
.B(n_498),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_733),
.B(n_528),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_735),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_735),
.B(n_502),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_651),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_SL g871 ( 
.A(n_604),
.B(n_365),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_652),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_757),
.A2(n_487),
.B(n_395),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_755),
.B(n_502),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_703),
.A2(n_527),
.B1(n_524),
.B2(n_512),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_703),
.A2(n_368),
.B(n_508),
.C(n_512),
.Y(n_876)
);

CKINVDCx8_ASAP7_75t_R g877 ( 
.A(n_698),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_618),
.Y(n_878)
);

NOR2x1_ASAP7_75t_L g879 ( 
.A(n_687),
.B(n_508),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_663),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_759),
.A2(n_487),
.B(n_395),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_628),
.B(n_443),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_768),
.A2(n_443),
.B1(n_395),
.B2(n_388),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_642),
.B(n_448),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_644),
.B(n_448),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_647),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_666),
.Y(n_887)
);

BUFx4f_ASAP7_75t_L g888 ( 
.A(n_758),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_615),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_758),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_646),
.A2(n_487),
.B(n_396),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_765),
.A2(n_771),
.B(n_769),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_656),
.B(n_448),
.Y(n_893)
);

OAI321xp33_ASAP7_75t_L g894 ( 
.A1(n_638),
.A2(n_2),
.A3(n_5),
.B1(n_6),
.B2(n_9),
.C(n_10),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_764),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_706),
.A2(n_448),
.B(n_487),
.C(n_396),
.Y(n_896)
);

AOI21x1_ASAP7_75t_L g897 ( 
.A1(n_681),
.A2(n_396),
.B(n_146),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_SL g898 ( 
.A(n_697),
.B(n_142),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_665),
.B(n_2),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_680),
.B(n_396),
.Y(n_900)
);

AOI21x1_ASAP7_75t_L g901 ( 
.A1(n_682),
.A2(n_396),
.B(n_135),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_646),
.A2(n_396),
.B(n_133),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_772),
.A2(n_396),
.B(n_132),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_650),
.A2(n_396),
.B(n_130),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_708),
.B(n_12),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_764),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_647),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_774),
.A2(n_396),
.B(n_125),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_647),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_680),
.B(n_123),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_680),
.B(n_14),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_631),
.A2(n_616),
.B1(n_648),
.B2(n_640),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_767),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_684),
.A2(n_121),
.B(n_116),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_634),
.B(n_637),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_767),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_639),
.B(n_14),
.Y(n_917)
);

NOR2x1p5_ASAP7_75t_L g918 ( 
.A(n_653),
.B(n_17),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_650),
.A2(n_115),
.B(n_114),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_SL g920 ( 
.A(n_711),
.B(n_113),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_705),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_641),
.B(n_17),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_707),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_722),
.A2(n_111),
.B(n_95),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_609),
.B(n_22),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_661),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_722),
.A2(n_93),
.B(n_89),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_723),
.A2(n_88),
.B(n_86),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_688),
.B(n_22),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_688),
.B(n_23),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_719),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_704),
.A2(n_79),
.B1(n_74),
.B2(n_73),
.Y(n_932)
);

NOR2xp67_ASAP7_75t_L g933 ( 
.A(n_620),
.B(n_633),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_723),
.A2(n_25),
.B(n_26),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_709),
.A2(n_26),
.B(n_28),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_713),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_719),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_706),
.B(n_31),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_719),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_715),
.A2(n_31),
.B(n_32),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_672),
.B(n_33),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_658),
.A2(n_34),
.B(n_37),
.C(n_39),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_717),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_721),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_725),
.A2(n_726),
.B(n_734),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_710),
.B(n_41),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_655),
.A2(n_41),
.B(n_45),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_727),
.A2(n_47),
.B(n_48),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_736),
.B(n_47),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_704),
.A2(n_66),
.B1(n_50),
.B2(n_53),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_728),
.A2(n_49),
.B(n_55),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_672),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_732),
.A2(n_56),
.B(n_60),
.Y(n_953)
);

OAI21xp33_ASAP7_75t_L g954 ( 
.A1(n_751),
.A2(n_63),
.B(n_66),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_655),
.A2(n_719),
.B(n_748),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_740),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_695),
.A2(n_700),
.B(n_702),
.Y(n_957)
);

BUFx4f_ASAP7_75t_L g958 ( 
.A(n_694),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_699),
.B(n_742),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_696),
.B(n_677),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_786),
.B(n_661),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_829),
.B(n_740),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_800),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_878),
.B(n_761),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_871),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_899),
.B(n_745),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_859),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_860),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_805),
.B(n_694),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_938),
.A2(n_668),
.B(n_739),
.C(n_730),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_949),
.A2(n_630),
.B(n_622),
.C(n_763),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_779),
.B(n_694),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_868),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_796),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_805),
.B(n_643),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_931),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_784),
.B(n_679),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_775),
.A2(n_763),
.B(n_766),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_802),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_949),
.A2(n_760),
.B(n_770),
.C(n_724),
.Y(n_980)
);

BUFx4_ASAP7_75t_SL g981 ( 
.A(n_890),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_R g982 ( 
.A(n_926),
.B(n_720),
.Y(n_982)
);

OR2x6_ASAP7_75t_SL g983 ( 
.A(n_950),
.B(n_773),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_858),
.A2(n_667),
.B(n_752),
.C(n_806),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_793),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_888),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_812),
.B(n_752),
.Y(n_987)
);

INVx4_ASAP7_75t_L g988 ( 
.A(n_937),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_915),
.B(n_856),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_886),
.B(n_907),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_856),
.B(n_842),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_842),
.B(n_778),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_SL g993 ( 
.A1(n_877),
.A2(n_790),
.B1(n_889),
.B2(n_946),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_SL g994 ( 
.A(n_806),
.B(n_946),
.C(n_954),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_776),
.A2(n_957),
.B(n_792),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_808),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_804),
.B(n_794),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_825),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_888),
.Y(n_999)
);

OA22x2_ASAP7_75t_L g1000 ( 
.A1(n_947),
.A2(n_952),
.B1(n_789),
.B2(n_828),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_821),
.B(n_834),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_931),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_925),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_821),
.B(n_834),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_787),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_SL g1006 ( 
.A1(n_794),
.A2(n_919),
.B(n_902),
.C(n_904),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_956),
.B(n_917),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_810),
.A2(n_912),
.B1(n_781),
.B2(n_956),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_958),
.B(n_807),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_798),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_855),
.B(n_905),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_955),
.A2(n_845),
.B1(n_907),
.B2(n_909),
.Y(n_1012)
);

NOR2x1_ASAP7_75t_L g1013 ( 
.A(n_886),
.B(n_909),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_SL g1014 ( 
.A(n_894),
.B(n_905),
.C(n_911),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_795),
.A2(n_809),
.B(n_892),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_788),
.A2(n_814),
.B(n_826),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_870),
.B(n_872),
.Y(n_1017)
);

NAND2x1p5_ASAP7_75t_L g1018 ( 
.A(n_937),
.B(n_939),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_807),
.Y(n_1019)
);

OAI22x1_ASAP7_75t_L g1020 ( 
.A1(n_918),
.A2(n_818),
.B1(n_836),
.B2(n_910),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_880),
.B(n_887),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_799),
.A2(n_785),
.B(n_824),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_922),
.A2(n_941),
.B(n_930),
.C(n_929),
.Y(n_1023)
);

NAND3xp33_ASAP7_75t_SL g1024 ( 
.A(n_791),
.B(n_934),
.C(n_920),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_820),
.A2(n_823),
.B1(n_819),
.B2(n_783),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_921),
.B(n_936),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_797),
.A2(n_815),
.B(n_831),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_822),
.A2(n_816),
.B(n_837),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_923),
.B(n_943),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_945),
.A2(n_893),
.B(n_885),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_849),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_944),
.B(n_850),
.Y(n_1032)
);

CKINVDCx16_ASAP7_75t_R g1033 ( 
.A(n_791),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_895),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_906),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_960),
.A2(n_959),
.B1(n_932),
.B2(n_951),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_913),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_798),
.Y(n_1038)
);

OAI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_898),
.A2(n_935),
.B(n_953),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_SL g1040 ( 
.A1(n_876),
.A2(n_896),
.B(n_832),
.C(n_835),
.Y(n_1040)
);

O2A1O1Ixp5_ASAP7_75t_L g1041 ( 
.A1(n_876),
.A2(n_811),
.B(n_851),
.C(n_897),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_780),
.A2(n_783),
.B1(n_937),
.B2(n_939),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_SL g1043 ( 
.A1(n_839),
.A2(n_882),
.B(n_891),
.C(n_817),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_916),
.Y(n_1044)
);

BUFx8_ASAP7_75t_L g1045 ( 
.A(n_937),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_942),
.A2(n_874),
.B(n_847),
.C(n_782),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_862),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_874),
.B(n_780),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_884),
.A2(n_813),
.B(n_833),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_939),
.A2(n_848),
.B1(n_866),
.B2(n_864),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_958),
.A2(n_928),
.B(n_927),
.C(n_924),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_940),
.A2(n_948),
.B1(n_900),
.B2(n_801),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_939),
.A2(n_848),
.B1(n_798),
.B2(n_852),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_867),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_900),
.B(n_838),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_840),
.A2(n_841),
.B(n_844),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_851),
.A2(n_838),
.B(n_835),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_828),
.B(n_933),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_828),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_869),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_798),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_801),
.B(n_803),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_883),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_861),
.B(n_847),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_863),
.A2(n_865),
.B(n_879),
.C(n_875),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_852),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_803),
.B(n_832),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_782),
.A2(n_846),
.B(n_827),
.C(n_914),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_852),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_852),
.B(n_854),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_854),
.A2(n_843),
.B1(n_853),
.B2(n_873),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_857),
.A2(n_881),
.B(n_830),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_854),
.A2(n_830),
.B1(n_901),
.B2(n_903),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_854),
.B(n_830),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_908),
.A2(n_478),
.B(n_645),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_830),
.B(n_786),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_830),
.A2(n_478),
.B(n_645),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_775),
.A2(n_478),
.B(n_645),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_800),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_798),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_775),
.A2(n_478),
.B(n_645),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_786),
.A2(n_829),
.B1(n_779),
.B2(n_617),
.Y(n_1082)
);

CKINVDCx6p67_ASAP7_75t_R g1083 ( 
.A(n_890),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_777),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_SL g1085 ( 
.A1(n_856),
.A2(n_625),
.B(n_456),
.C(n_481),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_800),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_777),
.Y(n_1087)
);

OR2x6_ASAP7_75t_L g1088 ( 
.A(n_937),
.B(n_758),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_786),
.B(n_673),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_786),
.B(n_829),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_878),
.B(n_627),
.Y(n_1091)
);

AOI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_806),
.A2(n_737),
.B1(n_546),
.B2(n_488),
.C(n_804),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_926),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_786),
.A2(n_625),
.B1(n_806),
.B2(n_481),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_786),
.A2(n_829),
.B1(n_779),
.B2(n_617),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_798),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_878),
.B(n_627),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_786),
.A2(n_625),
.B(n_938),
.C(n_779),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_784),
.B(n_654),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_798),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_777),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_786),
.B(n_829),
.Y(n_1102)
);

OAI22x1_ASAP7_75t_L g1103 ( 
.A1(n_918),
.A2(n_530),
.B1(n_480),
.B2(n_546),
.Y(n_1103)
);

INVx5_ASAP7_75t_L g1104 ( 
.A(n_830),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_878),
.Y(n_1105)
);

INVxp67_ASAP7_75t_SL g1106 ( 
.A(n_786),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_786),
.B(n_829),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_1033),
.Y(n_1108)
);

OA21x2_ASAP7_75t_L g1109 ( 
.A1(n_1041),
.A2(n_1015),
.B(n_1030),
.Y(n_1109)
);

OAI21xp33_ASAP7_75t_L g1110 ( 
.A1(n_1094),
.A2(n_1092),
.B(n_1004),
.Y(n_1110)
);

BUFx10_ASAP7_75t_L g1111 ( 
.A(n_964),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_997),
.A2(n_1025),
.A3(n_1098),
.B(n_1065),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_997),
.A2(n_1095),
.A3(n_1082),
.B(n_1073),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1085),
.A2(n_994),
.B(n_966),
.C(n_1090),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_1105),
.Y(n_1115)
);

OR2x6_ASAP7_75t_L g1116 ( 
.A(n_1088),
.B(n_990),
.Y(n_1116)
);

AND2x6_ASAP7_75t_L g1117 ( 
.A(n_990),
.B(n_1013),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_995),
.A2(n_1107),
.B(n_1102),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_971),
.A2(n_984),
.B(n_980),
.C(n_1008),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_994),
.A2(n_964),
.B1(n_977),
.B2(n_987),
.Y(n_1120)
);

AOI221xp5_ASAP7_75t_L g1121 ( 
.A1(n_1014),
.A2(n_991),
.B1(n_1103),
.B2(n_1106),
.C(n_993),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_977),
.A2(n_1099),
.B1(n_965),
.B2(n_961),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1105),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1028),
.A2(n_1078),
.B(n_1081),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1017),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1022),
.A2(n_1016),
.B(n_978),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_989),
.A2(n_1011),
.B(n_962),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1027),
.A2(n_1056),
.B(n_1049),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1106),
.A2(n_1075),
.B(n_1043),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_1083),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1001),
.B(n_1089),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1012),
.A2(n_1071),
.B(n_1057),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1091),
.B(n_1097),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1021),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1026),
.B(n_1032),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1047),
.B(n_1029),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1006),
.A2(n_1051),
.B(n_1068),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1005),
.Y(n_1138)
);

BUFx12f_ASAP7_75t_L g1139 ( 
.A(n_985),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_972),
.A2(n_1076),
.B(n_1036),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1091),
.B(n_1097),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1006),
.A2(n_1077),
.B(n_1023),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1035),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_992),
.B(n_1054),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1003),
.B(n_969),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_969),
.B(n_975),
.Y(n_1146)
);

AOI221x1_ASAP7_75t_L g1147 ( 
.A1(n_1039),
.A2(n_970),
.B1(n_1024),
.B2(n_1020),
.C(n_1050),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1000),
.A2(n_1036),
.B1(n_1007),
.B2(n_1014),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1072),
.A2(n_1041),
.B(n_1062),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1046),
.A2(n_1002),
.B(n_976),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1040),
.A2(n_1104),
.B(n_1052),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1045),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_963),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1055),
.A2(n_1048),
.A3(n_1063),
.B(n_1053),
.Y(n_1154)
);

AOI221x1_ASAP7_75t_L g1155 ( 
.A1(n_1024),
.A2(n_975),
.B1(n_1064),
.B2(n_1055),
.C(n_1048),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1104),
.A2(n_1052),
.B(n_1060),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1031),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1093),
.Y(n_1158)
);

AO32x2_ASAP7_75t_L g1159 ( 
.A1(n_1042),
.A2(n_983),
.A3(n_988),
.B1(n_1067),
.B2(n_968),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_976),
.A2(n_1002),
.B(n_1074),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1104),
.A2(n_1070),
.B(n_1009),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1031),
.B(n_1086),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_974),
.B(n_1087),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_967),
.B(n_973),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1079),
.B(n_998),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_979),
.B(n_1084),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1044),
.A2(n_1101),
.B(n_996),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1019),
.B(n_1034),
.Y(n_1168)
);

AOI221xp5_ASAP7_75t_SL g1169 ( 
.A1(n_1058),
.A2(n_1069),
.B1(n_1019),
.B2(n_1038),
.C(n_1100),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1061),
.B(n_986),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1104),
.A2(n_1018),
.B(n_1096),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1066),
.A2(n_999),
.B(n_1059),
.C(n_1100),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1018),
.A2(n_1066),
.B(n_988),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1088),
.A2(n_1045),
.B(n_982),
.C(n_981),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_982),
.B(n_1088),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1010),
.A2(n_1038),
.B(n_1080),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_981),
.Y(n_1177)
);

CKINVDCx6p67_ASAP7_75t_R g1178 ( 
.A(n_1010),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1010),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1038),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1096),
.B(n_1100),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1096),
.A2(n_1100),
.B(n_995),
.Y(n_1182)
);

AOI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1012),
.A2(n_1049),
.B(n_1025),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_997),
.A2(n_1095),
.B(n_1082),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1017),
.Y(n_1185)
);

CKINVDCx11_ASAP7_75t_R g1186 ( 
.A(n_1033),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1094),
.A2(n_327),
.B1(n_994),
.B2(n_1004),
.Y(n_1187)
);

AOI31xp67_ASAP7_75t_L g1188 ( 
.A1(n_1008),
.A2(n_1000),
.A3(n_1094),
.B(n_427),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1017),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_994),
.A2(n_1092),
.B1(n_806),
.B2(n_997),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_SL g1191 ( 
.A1(n_1092),
.A2(n_737),
.B1(n_949),
.B2(n_638),
.C(n_745),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1015),
.A2(n_1028),
.B(n_995),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_997),
.A2(n_1025),
.A3(n_1098),
.B(n_1065),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1099),
.B(n_654),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1015),
.A2(n_1028),
.B(n_995),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_SL g1196 ( 
.A1(n_1006),
.A2(n_1085),
.B(n_1098),
.C(n_970),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1015),
.A2(n_1028),
.B(n_995),
.Y(n_1197)
);

AOI221xp5_ASAP7_75t_SL g1198 ( 
.A1(n_1092),
.A2(n_737),
.B1(n_949),
.B2(n_638),
.C(n_745),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1105),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1107),
.B(n_1090),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1017),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1017),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1083),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1017),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_995),
.A2(n_1030),
.B(n_786),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1105),
.Y(n_1206)
);

AOI221x1_ASAP7_75t_L g1207 ( 
.A1(n_994),
.A2(n_806),
.B1(n_997),
.B2(n_1039),
.C(n_938),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1094),
.A2(n_1102),
.B(n_1107),
.C(n_1090),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1083),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1107),
.B(n_1090),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_995),
.A2(n_1030),
.B(n_786),
.Y(n_1211)
);

CKINVDCx8_ASAP7_75t_R g1212 ( 
.A(n_1033),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1015),
.A2(n_1028),
.B(n_995),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1107),
.B(n_1090),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1107),
.B(n_1090),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1094),
.A2(n_1098),
.B(n_786),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1015),
.A2(n_1028),
.B(n_995),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_995),
.A2(n_1030),
.B(n_786),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1083),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1107),
.B(n_1090),
.Y(n_1220)
);

NAND2x1_ASAP7_75t_L g1221 ( 
.A(n_990),
.B(n_988),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_995),
.A2(n_1030),
.B(n_786),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_SL g1223 ( 
.A(n_1033),
.B(n_888),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1015),
.A2(n_1028),
.B(n_995),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1015),
.A2(n_1028),
.B(n_995),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_997),
.A2(n_1025),
.A3(n_1098),
.B(n_1065),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1037),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1017),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_997),
.A2(n_1025),
.A3(n_1098),
.B(n_1065),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_SL g1230 ( 
.A1(n_1006),
.A2(n_1085),
.B(n_1098),
.C(n_970),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1017),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1015),
.A2(n_1028),
.B(n_995),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_995),
.A2(n_1030),
.B(n_786),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_995),
.A2(n_1030),
.B(n_786),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1037),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_995),
.A2(n_1030),
.B(n_786),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_990),
.Y(n_1237)
);

NAND2x1p5_ASAP7_75t_L g1238 ( 
.A(n_990),
.B(n_886),
.Y(n_1238)
);

BUFx10_ASAP7_75t_L g1239 ( 
.A(n_964),
.Y(n_1239)
);

AO32x2_ASAP7_75t_L g1240 ( 
.A1(n_1082),
.A2(n_1095),
.A3(n_1025),
.B1(n_1073),
.B2(n_1012),
.Y(n_1240)
);

NAND3xp33_ASAP7_75t_SL g1241 ( 
.A(n_1094),
.B(n_812),
.C(n_1092),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1001),
.B(n_1004),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1107),
.B(n_1090),
.Y(n_1243)
);

AOI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1012),
.A2(n_1049),
.B(n_1025),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_L g1245 ( 
.A(n_1093),
.B(n_609),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_995),
.A2(n_1030),
.B(n_786),
.Y(n_1246)
);

NAND3x1_ASAP7_75t_L g1247 ( 
.A(n_1092),
.B(n_806),
.C(n_737),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1094),
.A2(n_1098),
.B(n_786),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1001),
.B(n_1004),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1015),
.A2(n_1028),
.B(n_995),
.Y(n_1250)
);

INVx8_ASAP7_75t_L g1251 ( 
.A(n_1116),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1241),
.A2(n_1190),
.B1(n_1110),
.B2(n_1187),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1241),
.A2(n_1190),
.B1(n_1120),
.B2(n_1121),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1115),
.Y(n_1254)
);

INVx4_ASAP7_75t_L g1255 ( 
.A(n_1116),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1121),
.A2(n_1249),
.B1(n_1242),
.B2(n_1148),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1143),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1242),
.A2(n_1249),
.B1(n_1184),
.B2(n_1216),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1248),
.A2(n_1146),
.B1(n_1133),
.B2(n_1122),
.Y(n_1259)
);

BUFx10_ASAP7_75t_L g1260 ( 
.A(n_1158),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_1116),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1133),
.A2(n_1194),
.B1(n_1127),
.B2(n_1141),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1153),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1123),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1206),
.Y(n_1265)
);

OAI22x1_ASAP7_75t_SL g1266 ( 
.A1(n_1108),
.A2(n_1177),
.B1(n_1186),
.B2(n_1212),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1131),
.A2(n_1140),
.B1(n_1200),
.B2(n_1210),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1214),
.A2(n_1220),
.B1(n_1215),
.B2(n_1243),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1111),
.A2(n_1239),
.B1(n_1145),
.B2(n_1135),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1139),
.Y(n_1270)
);

OAI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1223),
.A2(n_1207),
.B1(n_1144),
.B2(n_1136),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1125),
.A2(n_1204),
.B1(n_1202),
.B2(n_1231),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1164),
.Y(n_1273)
);

NAND2x1p5_ASAP7_75t_L g1274 ( 
.A(n_1237),
.B(n_1221),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1160),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1134),
.A2(n_1228),
.B1(n_1185),
.B2(n_1201),
.Y(n_1276)
);

CKINVDCx9p33_ASAP7_75t_R g1277 ( 
.A(n_1170),
.Y(n_1277)
);

CKINVDCx6p67_ASAP7_75t_R g1278 ( 
.A(n_1152),
.Y(n_1278)
);

BUFx12f_ASAP7_75t_L g1279 ( 
.A(n_1175),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1199),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1247),
.A2(n_1189),
.B1(n_1191),
.B2(n_1198),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1245),
.A2(n_1119),
.B1(n_1208),
.B2(n_1164),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1165),
.Y(n_1283)
);

INVx5_ASAP7_75t_L g1284 ( 
.A(n_1117),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1208),
.A2(n_1165),
.B1(n_1172),
.B2(n_1162),
.Y(n_1285)
);

OAI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1155),
.A2(n_1147),
.B1(n_1237),
.B2(n_1235),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1178),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1157),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1227),
.Y(n_1289)
);

CKINVDCx6p67_ASAP7_75t_R g1290 ( 
.A(n_1130),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1203),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_R g1292 ( 
.A1(n_1166),
.A2(n_1163),
.B1(n_1157),
.B2(n_1174),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1137),
.A2(n_1166),
.B1(n_1142),
.B2(n_1118),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1167),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1114),
.A2(n_1174),
.B(n_1151),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1159),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1179),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1142),
.A2(n_1118),
.B1(n_1156),
.B2(n_1151),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_1181),
.Y(n_1299)
);

INVx4_ASAP7_75t_L g1300 ( 
.A(n_1117),
.Y(n_1300)
);

BUFx12f_ASAP7_75t_L g1301 ( 
.A(n_1209),
.Y(n_1301)
);

OAI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_1114),
.A2(n_1156),
.B(n_1129),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1238),
.A2(n_1168),
.B1(n_1161),
.B2(n_1219),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1129),
.A2(n_1161),
.B1(n_1117),
.B2(n_1149),
.Y(n_1304)
);

BUFx8_ASAP7_75t_L g1305 ( 
.A(n_1117),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_1180),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1117),
.A2(n_1188),
.B1(n_1238),
.B2(n_1126),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1205),
.A2(n_1233),
.B1(n_1246),
.B2(n_1236),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1205),
.A2(n_1233),
.B1(n_1246),
.B2(n_1236),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1211),
.A2(n_1234),
.B1(n_1222),
.B2(n_1218),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1211),
.A2(n_1234),
.B1(n_1222),
.B2(n_1218),
.Y(n_1311)
);

INVx6_ASAP7_75t_L g1312 ( 
.A(n_1169),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1173),
.A2(n_1244),
.B1(n_1183),
.B2(n_1171),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1112),
.B(n_1226),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1182),
.A2(n_1126),
.B1(n_1109),
.B2(n_1176),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1182),
.A2(n_1109),
.B1(n_1128),
.B2(n_1124),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1192),
.A2(n_1197),
.B1(n_1232),
.B2(n_1225),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1132),
.A2(n_1112),
.B1(n_1229),
.B2(n_1226),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1154),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1193),
.B(n_1229),
.Y(n_1320)
);

INVx6_ASAP7_75t_L g1321 ( 
.A(n_1154),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1195),
.A2(n_1217),
.B1(n_1224),
.B2(n_1250),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1159),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1159),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1159),
.Y(n_1325)
);

NAND2x1p5_ASAP7_75t_L g1326 ( 
.A(n_1213),
.B(n_1193),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1196),
.A2(n_1230),
.B1(n_1226),
.B2(n_1229),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1229),
.B(n_1113),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_SL g1329 ( 
.A(n_1196),
.Y(n_1329)
);

INVx6_ASAP7_75t_L g1330 ( 
.A(n_1230),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1113),
.B(n_1240),
.Y(n_1331)
);

BUFx8_ASAP7_75t_L g1332 ( 
.A(n_1240),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1113),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1240),
.A2(n_1094),
.B1(n_1210),
.B2(n_1200),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1240),
.A2(n_1241),
.B1(n_1190),
.B2(n_994),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1133),
.A2(n_408),
.B1(n_1004),
.B2(n_327),
.Y(n_1336)
);

OAI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1120),
.A2(n_408),
.B1(n_1094),
.B2(n_1187),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1241),
.A2(n_1247),
.B1(n_1110),
.B2(n_1190),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1115),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1116),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1116),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1206),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1150),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1157),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1241),
.A2(n_1190),
.B1(n_994),
.B2(n_1110),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1138),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1200),
.A2(n_1094),
.B1(n_1214),
.B2(n_1210),
.Y(n_1347)
);

CKINVDCx11_ASAP7_75t_R g1348 ( 
.A(n_1212),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1241),
.A2(n_1190),
.B1(n_994),
.B2(n_1110),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1241),
.A2(n_1190),
.B1(n_994),
.B2(n_1110),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1115),
.Y(n_1351)
);

INVx6_ASAP7_75t_L g1352 ( 
.A(n_1116),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1138),
.Y(n_1353)
);

INVx6_ASAP7_75t_L g1354 ( 
.A(n_1116),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1241),
.A2(n_1190),
.B1(n_994),
.B2(n_1110),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1241),
.A2(n_1190),
.B1(n_994),
.B2(n_1110),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1186),
.Y(n_1357)
);

BUFx12f_ASAP7_75t_L g1358 ( 
.A(n_1186),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1241),
.A2(n_1190),
.B1(n_994),
.B2(n_1110),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1120),
.B(n_1094),
.Y(n_1360)
);

INVx6_ASAP7_75t_L g1361 ( 
.A(n_1116),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1200),
.A2(n_1094),
.B1(n_1214),
.B2(n_1210),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1133),
.A2(n_408),
.B1(n_1004),
.B2(n_327),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1190),
.B(n_997),
.Y(n_1364)
);

AOI21xp33_ASAP7_75t_L g1365 ( 
.A1(n_1190),
.A2(n_1001),
.B(n_1085),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1138),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1190),
.A2(n_480),
.B(n_1187),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1116),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1241),
.A2(n_1190),
.B1(n_994),
.B2(n_1110),
.Y(n_1369)
);

INVx6_ASAP7_75t_L g1370 ( 
.A(n_1116),
.Y(n_1370)
);

CKINVDCx9p33_ASAP7_75t_R g1371 ( 
.A(n_1133),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1200),
.A2(n_1094),
.B1(n_1214),
.B2(n_1210),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1298),
.A2(n_1316),
.B(n_1326),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1284),
.B(n_1300),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1264),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1326),
.A2(n_1309),
.B(n_1308),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1252),
.A2(n_1364),
.B1(n_1360),
.B2(n_1253),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_SL g1378 ( 
.A1(n_1300),
.A2(n_1295),
.B(n_1282),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1302),
.A2(n_1313),
.B(n_1360),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1288),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1364),
.B(n_1334),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1333),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1344),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1255),
.B(n_1261),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1348),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1314),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1344),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1314),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1367),
.B(n_1338),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1320),
.Y(n_1390)
);

BUFx2_ASAP7_75t_SL g1391 ( 
.A(n_1284),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1320),
.Y(n_1392)
);

AOI21xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1337),
.A2(n_1350),
.B(n_1369),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1254),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1267),
.B(n_1347),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1275),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1328),
.Y(n_1397)
);

AOI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1318),
.A2(n_1303),
.B(n_1285),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1310),
.A2(n_1311),
.B(n_1322),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1305),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1305),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1293),
.A2(n_1327),
.B(n_1331),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1319),
.B(n_1323),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1362),
.B(n_1372),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1317),
.A2(n_1343),
.B(n_1315),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1321),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1323),
.Y(n_1407)
);

INVxp67_ASAP7_75t_L g1408 ( 
.A(n_1265),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1305),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1324),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1304),
.A2(n_1335),
.B(n_1325),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1345),
.A2(n_1355),
.B1(n_1349),
.B2(n_1359),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1332),
.A2(n_1329),
.B1(n_1330),
.B2(n_1312),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1257),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1294),
.A2(n_1366),
.B(n_1257),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1366),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1348),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1312),
.A2(n_1330),
.B1(n_1273),
.B2(n_1283),
.Y(n_1418)
);

A2O1A1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1356),
.A2(n_1365),
.B(n_1336),
.C(n_1363),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1296),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1268),
.B(n_1258),
.Y(n_1421)
);

OR2x6_ASAP7_75t_L g1422 ( 
.A(n_1251),
.B(n_1341),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1259),
.A2(n_1281),
.B1(n_1256),
.B2(n_1292),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1262),
.B(n_1299),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1342),
.B(n_1339),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1263),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1272),
.A2(n_1276),
.B1(n_1312),
.B2(n_1269),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1330),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1346),
.Y(n_1429)
);

OR2x6_ASAP7_75t_L g1430 ( 
.A(n_1251),
.B(n_1352),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1353),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1332),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1332),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1255),
.B(n_1368),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1341),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1329),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1274),
.A2(n_1289),
.B(n_1307),
.Y(n_1437)
);

OAI211xp5_ASAP7_75t_L g1438 ( 
.A1(n_1419),
.A2(n_1371),
.B(n_1291),
.C(n_1280),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1404),
.A2(n_1271),
.B(n_1286),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1426),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1395),
.B(n_1351),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1415),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1423),
.A2(n_1306),
.B1(n_1312),
.B2(n_1370),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1426),
.Y(n_1444)
);

A2O1A1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1393),
.A2(n_1251),
.B(n_1340),
.C(n_1306),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1425),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1386),
.B(n_1254),
.Y(n_1447)
);

AOI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1393),
.A2(n_1339),
.B1(n_1280),
.B2(n_1266),
.C(n_1289),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1408),
.B(n_1260),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1389),
.B(n_1385),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1386),
.B(n_1340),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1381),
.B(n_1380),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1412),
.A2(n_1395),
.B(n_1421),
.C(n_1427),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1412),
.A2(n_1251),
.B(n_1277),
.C(n_1287),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_SL g1455 ( 
.A1(n_1421),
.A2(n_1370),
.B(n_1361),
.C(n_1354),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1420),
.B(n_1297),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1377),
.A2(n_1357),
.B(n_1270),
.Y(n_1457)
);

A2O1A1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1413),
.A2(n_1287),
.B(n_1354),
.C(n_1352),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1417),
.B(n_1260),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1375),
.B(n_1361),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1427),
.A2(n_1361),
.B1(n_1352),
.B2(n_1354),
.Y(n_1461)
);

NOR2x1_ASAP7_75t_SL g1462 ( 
.A(n_1391),
.B(n_1358),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1394),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1379),
.A2(n_1354),
.B1(n_1352),
.B2(n_1357),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1424),
.B(n_1260),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1376),
.A2(n_1270),
.B(n_1279),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1383),
.B(n_1297),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1424),
.A2(n_1278),
.B1(n_1290),
.B2(n_1279),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1374),
.B(n_1301),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1387),
.B(n_1287),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1376),
.A2(n_1287),
.B(n_1290),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1388),
.B(n_1278),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1403),
.Y(n_1473)
);

INVxp67_ASAP7_75t_L g1474 ( 
.A(n_1429),
.Y(n_1474)
);

AND2x6_ASAP7_75t_L g1475 ( 
.A(n_1428),
.B(n_1291),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1379),
.A2(n_1301),
.B1(n_1384),
.B2(n_1434),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1373),
.A2(n_1405),
.B(n_1399),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1388),
.B(n_1390),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1390),
.B(n_1392),
.Y(n_1479)
);

AND2x2_ASAP7_75t_SL g1480 ( 
.A(n_1402),
.B(n_1381),
.Y(n_1480)
);

AOI221x1_ASAP7_75t_SL g1481 ( 
.A1(n_1436),
.A2(n_1429),
.B1(n_1431),
.B2(n_1392),
.C(n_1397),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1407),
.B(n_1410),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1406),
.B(n_1384),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_R g1484 ( 
.A(n_1400),
.B(n_1401),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1398),
.A2(n_1399),
.B(n_1437),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1400),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1398),
.A2(n_1399),
.B(n_1437),
.Y(n_1487)
);

INVxp67_ASAP7_75t_SL g1488 ( 
.A(n_1442),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1440),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1444),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1473),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1480),
.B(n_1397),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1438),
.A2(n_1433),
.B1(n_1432),
.B2(n_1428),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1442),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1452),
.B(n_1420),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1480),
.B(n_1478),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1479),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1474),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1482),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1482),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1450),
.B(n_1435),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1477),
.B(n_1396),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1477),
.B(n_1396),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1481),
.B(n_1379),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1447),
.B(n_1379),
.Y(n_1505)
);

OAI222xp33_ASAP7_75t_L g1506 ( 
.A1(n_1453),
.A2(n_1433),
.B1(n_1432),
.B2(n_1422),
.C1(n_1430),
.C2(n_1436),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1477),
.B(n_1396),
.Y(n_1507)
);

AOI222xp33_ASAP7_75t_L g1508 ( 
.A1(n_1439),
.A2(n_1378),
.B1(n_1409),
.B2(n_1431),
.C1(n_1416),
.C2(n_1414),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1456),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1456),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1471),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1483),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1465),
.A2(n_1378),
.B1(n_1435),
.B2(n_1434),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1496),
.B(n_1485),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1511),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1496),
.B(n_1487),
.Y(n_1516)
);

AND2x2_ASAP7_75t_SL g1517 ( 
.A(n_1511),
.B(n_1466),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1502),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1492),
.B(n_1463),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1505),
.B(n_1494),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1496),
.B(n_1502),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1505),
.B(n_1451),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1503),
.B(n_1466),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1503),
.B(n_1466),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1504),
.A2(n_1457),
.B1(n_1443),
.B2(n_1448),
.C(n_1461),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1491),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1498),
.B(n_1476),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1503),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1498),
.B(n_1464),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1495),
.B(n_1471),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1489),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1508),
.A2(n_1441),
.B1(n_1446),
.B2(n_1475),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1489),
.Y(n_1533)
);

OAI33xp33_ASAP7_75t_L g1534 ( 
.A1(n_1504),
.A2(n_1418),
.A3(n_1468),
.B1(n_1460),
.B2(n_1470),
.B3(n_1467),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1490),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1488),
.A2(n_1507),
.B(n_1382),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1508),
.A2(n_1475),
.B1(n_1411),
.B2(n_1402),
.Y(n_1537)
);

AOI221xp5_ASAP7_75t_L g1538 ( 
.A1(n_1506),
.A2(n_1454),
.B1(n_1418),
.B2(n_1445),
.C(n_1455),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1520),
.B(n_1509),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1531),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1521),
.B(n_1512),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1531),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1521),
.B(n_1512),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1536),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1515),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1525),
.A2(n_1493),
.B1(n_1454),
.B2(n_1475),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1531),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1533),
.Y(n_1548)
);

NAND2xp33_ASAP7_75t_SL g1549 ( 
.A(n_1532),
.B(n_1484),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1533),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1533),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1520),
.B(n_1510),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1535),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1521),
.B(n_1512),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1518),
.B(n_1497),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1519),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1536),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1518),
.B(n_1497),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1520),
.B(n_1499),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1538),
.B(n_1445),
.Y(n_1560)
);

NOR3xp33_ASAP7_75t_SL g1561 ( 
.A(n_1534),
.B(n_1459),
.C(n_1493),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1536),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1525),
.A2(n_1475),
.B1(n_1513),
.B2(n_1411),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1536),
.Y(n_1564)
);

NAND4xp75_ASAP7_75t_L g1565 ( 
.A(n_1538),
.B(n_1449),
.C(n_1472),
.D(n_1501),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1518),
.B(n_1500),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1536),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1536),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1540),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1545),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1545),
.B(n_1515),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1541),
.B(n_1515),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1540),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1561),
.B(n_1519),
.Y(n_1574)
);

XNOR2x2_ASAP7_75t_L g1575 ( 
.A(n_1565),
.B(n_1526),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1541),
.B(n_1528),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1541),
.B(n_1528),
.Y(n_1577)
);

NAND2x1p5_ASAP7_75t_L g1578 ( 
.A(n_1545),
.B(n_1517),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1542),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1544),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1542),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1560),
.A2(n_1532),
.B(n_1537),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1561),
.B(n_1522),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1544),
.Y(n_1584)
);

NAND2xp33_ASAP7_75t_R g1585 ( 
.A(n_1565),
.B(n_1469),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1560),
.A2(n_1537),
.B(n_1517),
.Y(n_1586)
);

INVxp33_ASAP7_75t_L g1587 ( 
.A(n_1546),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1547),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1539),
.B(n_1552),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1555),
.B(n_1522),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1552),
.B(n_1530),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1543),
.B(n_1523),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1555),
.B(n_1522),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1544),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1555),
.B(n_1522),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1548),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1543),
.B(n_1523),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1564),
.Y(n_1598)
);

NAND4xp75_ASAP7_75t_L g1599 ( 
.A(n_1546),
.B(n_1517),
.C(n_1529),
.D(n_1523),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1554),
.B(n_1523),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1558),
.B(n_1514),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1558),
.B(n_1514),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1548),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1603),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1569),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1578),
.B(n_1554),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1578),
.B(n_1554),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1583),
.B(n_1550),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1569),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1578),
.B(n_1558),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1578),
.B(n_1566),
.Y(n_1611)
);

NOR3xp33_ASAP7_75t_L g1612 ( 
.A(n_1599),
.B(n_1549),
.C(n_1534),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1576),
.B(n_1577),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1583),
.B(n_1550),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1587),
.B(n_1556),
.Y(n_1615)
);

AOI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1587),
.A2(n_1549),
.B1(n_1563),
.B2(n_1529),
.C(n_1557),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1574),
.B(n_1551),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1581),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1576),
.B(n_1517),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1574),
.B(n_1582),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1575),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1582),
.B(n_1486),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1581),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1576),
.B(n_1517),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1577),
.B(n_1566),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1601),
.B(n_1552),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1601),
.B(n_1559),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1586),
.B(n_1486),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1599),
.A2(n_1563),
.B1(n_1458),
.B2(n_1527),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1571),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1570),
.B(n_1551),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1586),
.B(n_1602),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1603),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1575),
.B(n_1527),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1602),
.B(n_1559),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1573),
.B(n_1553),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1603),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1577),
.B(n_1566),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1604),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1620),
.B(n_1599),
.Y(n_1640)
);

A2O1A1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1612),
.A2(n_1575),
.B(n_1585),
.C(n_1458),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1615),
.Y(n_1642)
);

NAND4xp25_ASAP7_75t_L g1643 ( 
.A(n_1620),
.B(n_1585),
.C(n_1570),
.D(n_1595),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1604),
.Y(n_1644)
);

AO21x1_ASAP7_75t_L g1645 ( 
.A1(n_1634),
.A2(n_1571),
.B(n_1573),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1613),
.B(n_1571),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1621),
.A2(n_1562),
.B1(n_1568),
.B2(n_1557),
.C(n_1571),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1605),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1612),
.A2(n_1524),
.B1(n_1572),
.B2(n_1516),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1605),
.Y(n_1650)
);

XOR2x2_ASAP7_75t_L g1651 ( 
.A(n_1622),
.B(n_1462),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1609),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1613),
.B(n_1571),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1609),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1618),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1628),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1618),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1623),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1623),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1633),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1613),
.B(n_1572),
.Y(n_1661)
);

AOI211x1_ASAP7_75t_L g1662 ( 
.A1(n_1629),
.A2(n_1572),
.B(n_1590),
.C(n_1595),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1621),
.Y(n_1663)
);

AOI211xp5_ASAP7_75t_L g1664 ( 
.A1(n_1641),
.A2(n_1616),
.B(n_1629),
.C(n_1632),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1641),
.A2(n_1616),
.B1(n_1632),
.B2(n_1617),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1666)
);

NAND3xp33_ASAP7_75t_SL g1667 ( 
.A(n_1645),
.B(n_1617),
.C(n_1614),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1656),
.B(n_1608),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1649),
.A2(n_1608),
.B1(n_1614),
.B2(n_1630),
.Y(n_1669)
);

CKINVDCx20_ASAP7_75t_R g1670 ( 
.A(n_1651),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1646),
.Y(n_1671)
);

OAI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1640),
.A2(n_1630),
.B1(n_1626),
.B2(n_1627),
.C(n_1635),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1662),
.B(n_1630),
.Y(n_1673)
);

AOI211xp5_ASAP7_75t_L g1674 ( 
.A1(n_1645),
.A2(n_1611),
.B(n_1610),
.C(n_1619),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1646),
.B(n_1638),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1639),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1644),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1660),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1653),
.A2(n_1625),
.B1(n_1638),
.B2(n_1624),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_SL g1680 ( 
.A(n_1643),
.B(n_1637),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1653),
.B(n_1625),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1661),
.B(n_1626),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1666),
.Y(n_1683)
);

AOI211xp5_ASAP7_75t_L g1684 ( 
.A1(n_1665),
.A2(n_1647),
.B(n_1659),
.C(n_1658),
.Y(n_1684)
);

OAI222xp33_ASAP7_75t_L g1685 ( 
.A1(n_1669),
.A2(n_1661),
.B1(n_1611),
.B2(n_1610),
.C1(n_1627),
.C2(n_1635),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1664),
.A2(n_1651),
.B1(n_1655),
.B2(n_1654),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1667),
.A2(n_1650),
.B(n_1648),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1677),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1674),
.A2(n_1657),
.B(n_1652),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_L g1690 ( 
.A(n_1680),
.B(n_1637),
.C(n_1633),
.Y(n_1690)
);

AOI21xp33_ASAP7_75t_L g1691 ( 
.A1(n_1672),
.A2(n_1637),
.B(n_1633),
.Y(n_1691)
);

O2A1O1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1677),
.A2(n_1570),
.B(n_1624),
.C(n_1619),
.Y(n_1692)
);

NAND2x1_ASAP7_75t_L g1693 ( 
.A(n_1675),
.B(n_1570),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1678),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1687),
.A2(n_1680),
.B(n_1670),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1688),
.B(n_1671),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1686),
.A2(n_1673),
.B1(n_1668),
.B2(n_1676),
.C(n_1681),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1683),
.B(n_1682),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1684),
.B(n_1679),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1694),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1692),
.B(n_1690),
.Y(n_1701)
);

NAND2xp33_ASAP7_75t_SL g1702 ( 
.A(n_1693),
.B(n_1570),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1689),
.Y(n_1703)
);

AOI211x1_ASAP7_75t_SL g1704 ( 
.A1(n_1695),
.A2(n_1691),
.B(n_1685),
.C(n_1692),
.Y(n_1704)
);

NOR3xp33_ASAP7_75t_L g1705 ( 
.A(n_1703),
.B(n_1607),
.C(n_1606),
.Y(n_1705)
);

OAI321xp33_ASAP7_75t_L g1706 ( 
.A1(n_1701),
.A2(n_1699),
.A3(n_1697),
.B1(n_1696),
.B2(n_1698),
.C(n_1700),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1702),
.A2(n_1619),
.B(n_1624),
.C(n_1606),
.Y(n_1707)
);

OAI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1703),
.A2(n_1607),
.B1(n_1636),
.B2(n_1625),
.C(n_1593),
.Y(n_1708)
);

OAI21xp33_ASAP7_75t_L g1709 ( 
.A1(n_1705),
.A2(n_1631),
.B(n_1636),
.Y(n_1709)
);

AOI211xp5_ASAP7_75t_L g1710 ( 
.A1(n_1706),
.A2(n_1631),
.B(n_1568),
.C(n_1562),
.Y(n_1710)
);

OAI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1708),
.A2(n_1589),
.B1(n_1593),
.B2(n_1590),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_L g1712 ( 
.A(n_1704),
.B(n_1631),
.C(n_1589),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1707),
.A2(n_1631),
.B1(n_1564),
.B2(n_1567),
.C(n_1598),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1705),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1714),
.B(n_1592),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1712),
.Y(n_1716)
);

NOR2xp67_ASAP7_75t_L g1717 ( 
.A(n_1709),
.B(n_1579),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1710),
.Y(n_1718)
);

NOR3x2_ASAP7_75t_L g1719 ( 
.A(n_1711),
.B(n_1589),
.C(n_1591),
.Y(n_1719)
);

AOI21xp33_ASAP7_75t_L g1720 ( 
.A1(n_1716),
.A2(n_1713),
.B(n_1594),
.Y(n_1720)
);

AND4x1_ASAP7_75t_L g1721 ( 
.A(n_1718),
.B(n_1600),
.C(n_1597),
.D(n_1592),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1715),
.B(n_1579),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1721),
.A2(n_1717),
.B1(n_1719),
.B2(n_1591),
.C(n_1594),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1723),
.Y(n_1724)
);

INVxp33_ASAP7_75t_L g1725 ( 
.A(n_1724),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1724),
.B(n_1722),
.Y(n_1726)
);

AOI21xp33_ASAP7_75t_L g1727 ( 
.A1(n_1725),
.A2(n_1726),
.B(n_1720),
.Y(n_1727)
);

OAI22x1_ASAP7_75t_L g1728 ( 
.A1(n_1726),
.A2(n_1719),
.B1(n_1588),
.B2(n_1596),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1727),
.A2(n_1584),
.B(n_1580),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1728),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1730),
.Y(n_1731)
);

OAI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1731),
.A2(n_1729),
.B(n_1584),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1732),
.Y(n_1733)
);

AOI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1733),
.A2(n_1584),
.B1(n_1598),
.B2(n_1580),
.C(n_1594),
.Y(n_1734)
);

AOI211xp5_ASAP7_75t_L g1735 ( 
.A1(n_1734),
.A2(n_1580),
.B(n_1598),
.C(n_1584),
.Y(n_1735)
);


endmodule