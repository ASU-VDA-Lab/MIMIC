module fake_jpeg_10500_n_116 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_116);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_59),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_0),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_1),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_62),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_71),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_49),
.B1(n_54),
.B2(n_52),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_76),
.B1(n_16),
.B2(n_17),
.Y(n_96)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_83),
.Y(n_100)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_90)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_56),
.B1(n_51),
.B2(n_45),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_87),
.B(n_11),
.C(n_14),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_60),
.B(n_39),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_82),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_2),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_3),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_4),
.Y(n_86)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_5),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_94),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_19),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_100),
.B1(n_91),
.B2(n_96),
.Y(n_104)
);

NOR4xp25_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_100),
.C(n_98),
.D(n_95),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_102),
.B1(n_99),
.B2(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_72),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_88),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_70),
.C(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_25),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_97),
.B(n_27),
.Y(n_114)
);

OAI221xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.C(n_30),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);


endmodule