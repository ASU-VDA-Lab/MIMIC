module fake_netlist_6_4245_n_2039 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2039);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2039;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_128),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_193),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_43),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_70),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_40),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_46),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_72),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_105),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_97),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_3),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_123),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_203),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_156),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_110),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_117),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_152),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_108),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_52),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_161),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_29),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_142),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_66),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_91),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_171),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_153),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_107),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_100),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_112),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_137),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_96),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_175),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_146),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_115),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_169),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_131),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_144),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_160),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_111),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_11),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_165),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_35),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_55),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_0),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_31),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_44),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_162),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_118),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_74),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_126),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_116),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_61),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_36),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_130),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_101),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_40),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_4),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_69),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_31),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_78),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_48),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_87),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_138),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_127),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_170),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_134),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_64),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_192),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_176),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_70),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_84),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_99),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_27),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_125),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_92),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_33),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_172),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_5),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_5),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_179),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_10),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_77),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_24),
.Y(n_297)
);

BUFx10_ASAP7_75t_L g298 ( 
.A(n_158),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_197),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_11),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_38),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_109),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_173),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_196),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_66),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_9),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_37),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_63),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_16),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_51),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_191),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_90),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_95),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_114),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_21),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_143),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_155),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_34),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_181),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_80),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_166),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_189),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_164),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_10),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_27),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_1),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_68),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_102),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_72),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_201),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_88),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_124),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_48),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_121),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_59),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_174),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_185),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_190),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_135),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_81),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_94),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_89),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_187),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_119),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_198),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_43),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_199),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_39),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_30),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_154),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_145),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_33),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_20),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_76),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_25),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_54),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_58),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_36),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_45),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_63),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_53),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_29),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_18),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_44),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_3),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_41),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_57),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_46),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_15),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_64),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_139),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_82),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_86),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_6),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_37),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_17),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_177),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_67),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_93),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_15),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_74),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_13),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_157),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_133),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_13),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_57),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_69),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_14),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_151),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_35),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_45),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_22),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_149),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_106),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_30),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_42),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_188),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_148),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_205),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_51),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_54),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_20),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_184),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_9),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_79),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_19),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_206),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_41),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_34),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_68),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_183),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_168),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_38),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_180),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_186),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_218),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_224),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_218),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_213),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_213),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_257),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_208),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_257),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_220),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_220),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_333),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_221),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_221),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_270),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_234),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_242),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_270),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_327),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_388),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_388),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_384),
.B(n_0),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_234),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_211),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_235),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_210),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_237),
.B(n_1),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_251),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_235),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_333),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_333),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_212),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_333),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_333),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g449 ( 
.A(n_301),
.B(n_2),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_243),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_243),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_267),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_214),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_271),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_244),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_215),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_333),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_219),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_244),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_289),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_354),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_233),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_327),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_345),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_414),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_245),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_273),
.B(n_2),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_245),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_293),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_278),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_324),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_236),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_253),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_209),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_262),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_216),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_217),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_278),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_265),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_279),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_279),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_229),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_280),
.Y(n_483)
);

INVxp33_ASAP7_75t_SL g484 ( 
.A(n_266),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_269),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_280),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_222),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_291),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_223),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_272),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_275),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_232),
.B(n_6),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_324),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_324),
.B(n_7),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_281),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_225),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_291),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_299),
.Y(n_498)
);

NOR2xp67_ASAP7_75t_L g499 ( 
.A(n_349),
.B(n_7),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_378),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_287),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_299),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_297),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_232),
.B(n_8),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_317),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_378),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_306),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_317),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_229),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_307),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_260),
.B(n_8),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_227),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_319),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_319),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_320),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_320),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_228),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_309),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_334),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_260),
.B(n_12),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_444),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_442),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_442),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_442),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_444),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_422),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_422),
.B(n_231),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_442),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_474),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_457),
.B(n_238),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_492),
.B(n_415),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_445),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_445),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g534 ( 
.A(n_440),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_493),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_476),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_447),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_494),
.B(n_378),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_422),
.B(n_231),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_447),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_504),
.B(n_241),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_442),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_494),
.B(n_471),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_448),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_493),
.Y(n_545)
);

OA21x2_ASAP7_75t_L g546 ( 
.A1(n_448),
.A2(n_359),
.B(n_300),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_426),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_426),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_422),
.B(n_250),
.Y(n_549)
);

NOR2x1_ASAP7_75t_L g550 ( 
.A(n_520),
.B(n_250),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_416),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_418),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_424),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_419),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_425),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_511),
.B(n_239),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_427),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_428),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_430),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_437),
.B(n_252),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_419),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_439),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_500),
.B(n_240),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_443),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_506),
.B(n_246),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_450),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_451),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_436),
.A2(n_284),
.B1(n_353),
.B2(n_259),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_SL g569 ( 
.A(n_482),
.B(n_349),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_455),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_459),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_466),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_468),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_441),
.B(n_302),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_470),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_478),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_480),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_481),
.B(n_386),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_483),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_486),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_488),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_497),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_498),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_502),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_505),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_508),
.B(n_386),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_513),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_514),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_420),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_420),
.Y(n_590)
);

OA21x2_ASAP7_75t_L g591 ( 
.A1(n_515),
.A2(n_359),
.B(n_300),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_516),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_519),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_509),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_454),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_484),
.B(n_322),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_469),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_463),
.B(n_256),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_438),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_518),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_499),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_446),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_527),
.A2(n_433),
.B1(n_467),
.B2(n_387),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_596),
.B(n_464),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_535),
.B(n_421),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_555),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_591),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_527),
.A2(n_387),
.B1(n_368),
.B2(n_386),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_547),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_542),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_591),
.Y(n_612)
);

AND3x2_ASAP7_75t_L g613 ( 
.A(n_599),
.B(n_330),
.C(n_252),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_547),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_553),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_548),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_548),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_591),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_543),
.B(n_446),
.Y(n_619)
);

INVx6_ASAP7_75t_L g620 ( 
.A(n_575),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_596),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_525),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_591),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_543),
.B(n_453),
.Y(n_624)
);

OR2x6_ASAP7_75t_L g625 ( 
.A(n_601),
.B(n_334),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_591),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_553),
.Y(n_627)
);

INVxp67_ASAP7_75t_SL g628 ( 
.A(n_530),
.Y(n_628)
);

CKINVDCx6p67_ASAP7_75t_R g629 ( 
.A(n_534),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_591),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_542),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_535),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_546),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_601),
.B(n_518),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_534),
.B(n_477),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_574),
.B(n_453),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_553),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_525),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_526),
.B(n_337),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_574),
.B(n_487),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_546),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_532),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_546),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_555),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_546),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_545),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_542),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_543),
.B(n_456),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_541),
.B(n_489),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_546),
.Y(n_650)
);

INVx11_ASAP7_75t_L g651 ( 
.A(n_599),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_541),
.B(n_496),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_542),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_546),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_579),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_545),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_579),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_601),
.B(n_456),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_542),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_579),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_532),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_529),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_533),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_542),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_579),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_568),
.A2(n_569),
.B1(n_598),
.B2(n_449),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_595),
.B(n_458),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_529),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_530),
.B(n_458),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_526),
.B(n_337),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_533),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_568),
.B(n_550),
.C(n_594),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_563),
.B(n_565),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_579),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_555),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_601),
.B(n_462),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_542),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_601),
.B(n_595),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_531),
.B(n_462),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_553),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_537),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_536),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_569),
.A2(n_374),
.B1(n_390),
.B2(n_355),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_537),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_601),
.B(n_472),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_595),
.B(n_472),
.Y(n_686)
);

INVx8_ASAP7_75t_L g687 ( 
.A(n_527),
.Y(n_687)
);

INVx5_ASAP7_75t_L g688 ( 
.A(n_542),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_595),
.B(n_473),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_555),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_538),
.B(n_578),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_531),
.A2(n_517),
.B1(n_512),
.B2(n_423),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_522),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_540),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_540),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_527),
.A2(n_549),
.B1(n_539),
.B2(n_550),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_544),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_526),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_522),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_601),
.B(n_473),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_553),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_526),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_590),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_556),
.B(n_475),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_553),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_544),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_601),
.B(n_475),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_522),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_536),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_563),
.B(n_479),
.Y(n_710)
);

INVxp33_ASAP7_75t_L g711 ( 
.A(n_598),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_551),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_522),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_551),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_597),
.B(n_600),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_553),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_521),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_538),
.B(n_578),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_556),
.B(n_479),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_521),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_521),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_552),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_552),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_558),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_565),
.B(n_485),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_527),
.B(n_539),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_552),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_552),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_558),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_559),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_602),
.B(n_510),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_598),
.A2(n_602),
.B1(n_594),
.B2(n_600),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_562),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_562),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_553),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_523),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_571),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_571),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_527),
.B(n_485),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_597),
.B(n_490),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_557),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_557),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_597),
.B(n_490),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_572),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_572),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_597),
.B(n_491),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_573),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_573),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_559),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_576),
.Y(n_750)
);

BUFx10_ASAP7_75t_L g751 ( 
.A(n_539),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_597),
.B(n_341),
.Y(n_752)
);

AND2x6_ASAP7_75t_L g753 ( 
.A(n_539),
.B(n_251),
.Y(n_753)
);

OR2x6_ASAP7_75t_L g754 ( 
.A(n_600),
.B(n_341),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_523),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_590),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_L g757 ( 
.A(n_687),
.B(n_600),
.Y(n_757)
);

AO22x1_ASAP7_75t_L g758 ( 
.A1(n_740),
.A2(n_746),
.B1(n_743),
.B2(n_648),
.Y(n_758)
);

INVxp67_ASAP7_75t_SL g759 ( 
.A(n_726),
.Y(n_759)
);

NOR2xp67_ASAP7_75t_L g760 ( 
.A(n_649),
.B(n_603),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_673),
.B(n_539),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_628),
.B(n_539),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_608),
.A2(n_549),
.B1(n_618),
.B2(n_612),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_717),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_751),
.B(n_600),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_711),
.B(n_603),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_667),
.B(n_598),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_712),
.Y(n_768)
);

OAI22xp33_ASAP7_75t_SL g769 ( 
.A1(n_636),
.A2(n_423),
.B1(n_429),
.B2(n_421),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_710),
.B(n_549),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_698),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_725),
.B(n_549),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_629),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_712),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_696),
.B(n_679),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_704),
.B(n_491),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_719),
.B(n_549),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_667),
.B(n_549),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_686),
.B(n_538),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_751),
.B(n_251),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_686),
.B(n_575),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_689),
.B(n_575),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_689),
.B(n_575),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_717),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_751),
.B(n_669),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_678),
.B(n_251),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_SL g787 ( 
.A(n_640),
.B(n_652),
.C(n_666),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_675),
.B(n_575),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_675),
.B(n_557),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_720),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_619),
.B(n_495),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_732),
.B(n_251),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_606),
.B(n_590),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_714),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_690),
.B(n_557),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_714),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_690),
.B(n_557),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_724),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_720),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_691),
.B(n_718),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_724),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_691),
.B(n_557),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_607),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_608),
.A2(n_230),
.B(n_258),
.C(n_255),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_648),
.B(n_554),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_729),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_721),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_715),
.B(n_251),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_687),
.A2(n_524),
.B(n_523),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_718),
.B(n_557),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_698),
.B(n_557),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_624),
.B(n_495),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_739),
.B(n_283),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_729),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_733),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_687),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_687),
.B(n_639),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_733),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_687),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_672),
.B(n_501),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_702),
.B(n_639),
.Y(n_821)
);

BUFx6f_ASAP7_75t_SL g822 ( 
.A(n_632),
.Y(n_822)
);

INVx8_ASAP7_75t_L g823 ( 
.A(n_752),
.Y(n_823)
);

NOR2xp67_ASAP7_75t_L g824 ( 
.A(n_692),
.B(n_554),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_702),
.B(n_564),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_639),
.B(n_283),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_639),
.B(n_670),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_670),
.B(n_564),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_656),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_SL g830 ( 
.A(n_629),
.B(n_561),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_605),
.B(n_501),
.Y(n_831)
);

NOR2xp67_ASAP7_75t_L g832 ( 
.A(n_632),
.B(n_561),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_634),
.A2(n_589),
.B1(n_431),
.B2(n_452),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_753),
.B(n_247),
.Y(n_834)
);

BUFx6f_ASAP7_75t_SL g835 ( 
.A(n_646),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_662),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_670),
.B(n_734),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_670),
.B(n_283),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_734),
.B(n_564),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_736),
.A2(n_524),
.B(n_523),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_737),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_737),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_622),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_738),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_658),
.B(n_503),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_612),
.B(n_283),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_676),
.B(n_503),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_721),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_618),
.B(n_283),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_738),
.B(n_564),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_685),
.A2(n_589),
.B1(n_460),
.B2(n_461),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_722),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_700),
.B(n_507),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_707),
.B(n_507),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_722),
.Y(n_855)
);

NOR3xp33_ASAP7_75t_L g856 ( 
.A(n_606),
.B(n_731),
.C(n_646),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_752),
.A2(n_754),
.B1(n_666),
.B2(n_644),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_621),
.B(n_510),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_744),
.B(n_745),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_623),
.B(n_283),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_623),
.B(n_564),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_703),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_744),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_745),
.B(n_564),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_607),
.Y(n_865)
);

AO22x2_ASAP7_75t_L g866 ( 
.A1(n_633),
.A2(n_383),
.B1(n_343),
.B2(n_351),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_747),
.B(n_748),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_621),
.B(n_429),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_747),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_626),
.A2(n_368),
.B1(n_230),
.B2(n_381),
.Y(n_870)
);

BUFx5_ASAP7_75t_L g871 ( 
.A(n_626),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_621),
.B(n_432),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_703),
.B(n_432),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_748),
.B(n_434),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_750),
.B(n_434),
.Y(n_875)
);

INVxp33_ASAP7_75t_L g876 ( 
.A(n_635),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_630),
.B(n_564),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_750),
.B(n_706),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_622),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_644),
.B(n_578),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_706),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_683),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_752),
.A2(n_417),
.B1(n_465),
.B2(n_435),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_756),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_630),
.B(n_564),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_613),
.B(n_586),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_633),
.B(n_567),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_641),
.B(n_567),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_655),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_641),
.B(n_567),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_643),
.B(n_567),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_723),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_643),
.B(n_567),
.Y(n_893)
);

NOR2x1p5_ASAP7_75t_L g894 ( 
.A(n_756),
.B(n_435),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_645),
.B(n_567),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_620),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_655),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_657),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_645),
.B(n_567),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_604),
.B(n_586),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_651),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_657),
.B(n_567),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_723),
.Y(n_903)
);

NAND2xp33_ASAP7_75t_L g904 ( 
.A(n_753),
.B(n_248),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_660),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_651),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_727),
.Y(n_907)
);

NAND2x1p5_ASAP7_75t_L g908 ( 
.A(n_650),
.B(n_654),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_638),
.B(n_586),
.Y(n_909)
);

CKINVDCx11_ASAP7_75t_R g910 ( 
.A(n_662),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_650),
.B(n_577),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_654),
.B(n_577),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_683),
.B(n_576),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_665),
.B(n_577),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_674),
.B(n_577),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_674),
.B(n_638),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_642),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_752),
.B(n_593),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_642),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_661),
.B(n_577),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_625),
.A2(n_593),
.B(n_592),
.C(n_581),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_659),
.Y(n_922)
);

NOR3xp33_ASAP7_75t_L g923 ( 
.A(n_668),
.B(n_584),
.C(n_581),
.Y(n_923)
);

NAND2xp33_ASAP7_75t_L g924 ( 
.A(n_753),
.B(n_249),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_752),
.A2(n_560),
.B1(n_321),
.B2(n_411),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_661),
.B(n_577),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_803),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_763),
.A2(n_888),
.B(n_887),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_896),
.A2(n_627),
.B(n_615),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_761),
.B(n_754),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_758),
.B(n_759),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_803),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_770),
.B(n_754),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_787),
.B(n_668),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_775),
.A2(n_754),
.B(n_663),
.C(n_681),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_SL g936 ( 
.A(n_836),
.B(n_682),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_896),
.A2(n_627),
.B(n_615),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_763),
.A2(n_754),
.B(n_625),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_772),
.B(n_779),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_800),
.A2(n_778),
.B1(n_820),
.B2(n_900),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_767),
.B(n_625),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_804),
.A2(n_663),
.B(n_681),
.C(n_671),
.Y(n_942)
);

BUFx4f_ASAP7_75t_L g943 ( 
.A(n_901),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_871),
.B(n_671),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_871),
.B(n_684),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_804),
.A2(n_684),
.B(n_695),
.C(n_694),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_762),
.A2(n_627),
.B(n_615),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_773),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_776),
.B(n_682),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_910),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_777),
.B(n_625),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_890),
.A2(n_625),
.B(n_694),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_870),
.A2(n_609),
.B1(n_255),
.B2(n_290),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_781),
.B(n_782),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_760),
.B(n_709),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_783),
.B(n_695),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_870),
.A2(n_258),
.B1(n_292),
.B2(n_290),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_766),
.B(n_709),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_827),
.A2(n_680),
.B(n_637),
.Y(n_959)
);

NAND3xp33_ASAP7_75t_SL g960 ( 
.A(n_776),
.B(n_325),
.C(n_318),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_843),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_871),
.B(n_768),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_871),
.B(n_697),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_922),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_879),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_918),
.A2(n_351),
.B(n_372),
.C(n_343),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_823),
.B(n_906),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_862),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_829),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_791),
.A2(n_620),
.B1(n_753),
.B2(n_697),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_821),
.A2(n_680),
.B(n_637),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_891),
.A2(n_680),
.B(n_637),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_846),
.A2(n_585),
.B(n_592),
.C(n_584),
.Y(n_973)
);

OAI321xp33_ASAP7_75t_L g974 ( 
.A1(n_820),
.A2(n_305),
.A3(n_365),
.B1(n_396),
.B2(n_295),
.C(n_292),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_893),
.A2(n_716),
.B(n_705),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_857),
.A2(n_310),
.B1(n_308),
.B2(n_305),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_879),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_832),
.B(n_585),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_SL g979 ( 
.A1(n_846),
.A2(n_389),
.B(n_393),
.C(n_372),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_823),
.B(n_620),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_880),
.B(n_254),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_895),
.A2(n_728),
.B(n_727),
.Y(n_982)
);

INVx11_ASAP7_75t_L g983 ( 
.A(n_822),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_899),
.A2(n_730),
.B(n_728),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_849),
.A2(n_617),
.B(n_610),
.C(n_614),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_771),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_889),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_911),
.A2(n_716),
.B(n_705),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_897),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_816),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_871),
.B(n_620),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_833),
.B(n_610),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_871),
.B(n_611),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_791),
.B(n_812),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_805),
.B(n_256),
.Y(n_995)
);

AOI21xp33_ASAP7_75t_L g996 ( 
.A1(n_837),
.A2(n_389),
.B(n_383),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_774),
.B(n_611),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_812),
.B(n_326),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_912),
.A2(n_885),
.B(n_757),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_802),
.A2(n_716),
.B(n_705),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_873),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_810),
.A2(n_741),
.B(n_735),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_898),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_905),
.Y(n_1004)
);

BUFx4f_ASAP7_75t_L g1005 ( 
.A(n_886),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_880),
.B(n_845),
.Y(n_1006)
);

NOR2xp67_ASAP7_75t_L g1007 ( 
.A(n_845),
.B(n_614),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_811),
.A2(n_741),
.B(n_735),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_908),
.A2(n_749),
.B(n_730),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_918),
.A2(n_393),
.B(n_412),
.C(n_398),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_794),
.B(n_611),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_849),
.A2(n_617),
.B(n_616),
.C(n_749),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_825),
.A2(n_817),
.B(n_861),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_860),
.A2(n_616),
.B(n_398),
.C(n_407),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_922),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_796),
.B(n_631),
.Y(n_1016)
);

NOR2xp67_ASAP7_75t_L g1017 ( 
.A(n_847),
.B(n_693),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_771),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_798),
.B(n_631),
.Y(n_1019)
);

BUFx8_ASAP7_75t_L g1020 ( 
.A(n_822),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_801),
.B(n_631),
.Y(n_1021)
);

BUFx4f_ASAP7_75t_L g1022 ( 
.A(n_886),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_908),
.A2(n_677),
.B(n_647),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_861),
.A2(n_677),
.B(n_647),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_785),
.A2(n_753),
.B1(n_560),
.B2(n_741),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_806),
.B(n_814),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_884),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_817),
.A2(n_735),
.B(n_664),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_815),
.B(n_647),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_868),
.B(n_329),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_785),
.A2(n_753),
.B1(n_560),
.B2(n_677),
.Y(n_1031)
);

NOR3xp33_ASAP7_75t_L g1032 ( 
.A(n_868),
.B(n_412),
.C(n_407),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_877),
.A2(n_664),
.B(n_659),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_877),
.A2(n_664),
.B(n_659),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_922),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_847),
.A2(n_405),
.B(n_330),
.C(n_336),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_853),
.B(n_261),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_853),
.B(n_263),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_793),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_809),
.A2(n_699),
.B(n_693),
.Y(n_1040)
);

CKINVDCx10_ASAP7_75t_R g1041 ( 
.A(n_882),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_818),
.B(n_753),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_835),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_858),
.B(n_256),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_841),
.B(n_693),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_860),
.A2(n_336),
.B(n_405),
.C(n_559),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_828),
.A2(n_664),
.B(n_659),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_842),
.B(n_699),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_844),
.B(n_699),
.Y(n_1049)
);

NAND2x1_ASAP7_75t_L g1050 ( 
.A(n_819),
.B(n_659),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_863),
.B(n_708),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_854),
.B(n_264),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_764),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_792),
.A2(n_559),
.B(n_570),
.C(n_566),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_909),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_869),
.B(n_708),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_854),
.B(n_268),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_856),
.A2(n_560),
.B1(n_713),
.B2(n_708),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_881),
.B(n_713),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_916),
.A2(n_755),
.B(n_713),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_788),
.A2(n_664),
.B(n_701),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_784),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_874),
.A2(n_560),
.B(n_755),
.C(n_587),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_765),
.A2(n_742),
.B(n_701),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_922),
.Y(n_1065)
);

CKINVDCx10_ASAP7_75t_R g1066 ( 
.A(n_835),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_872),
.B(n_831),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_865),
.Y(n_1068)
);

AOI21x1_ASAP7_75t_L g1069 ( 
.A1(n_902),
.A2(n_528),
.B(n_524),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_878),
.B(n_755),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_872),
.B(n_335),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_831),
.B(n_876),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_790),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_865),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_874),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_859),
.B(n_867),
.Y(n_1076)
);

O2A1O1Ixp5_ASAP7_75t_L g1077 ( 
.A1(n_813),
.A2(n_560),
.B(n_582),
.C(n_588),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_909),
.B(n_701),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_799),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_765),
.A2(n_313),
.B1(n_274),
.B2(n_276),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_913),
.Y(n_1081)
);

O2A1O1Ixp5_ASAP7_75t_L g1082 ( 
.A1(n_813),
.A2(n_583),
.B(n_570),
.C(n_588),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_780),
.A2(n_742),
.B(n_701),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_917),
.B(n_742),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_823),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_919),
.B(n_742),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_780),
.A2(n_742),
.B(n_701),
.Y(n_1087)
);

BUFx4f_ASAP7_75t_L g1088 ( 
.A(n_816),
.Y(n_1088)
);

OAI21xp33_ASAP7_75t_L g1089 ( 
.A1(n_875),
.A2(n_851),
.B(n_923),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_807),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_848),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_883),
.B(n_348),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_824),
.Y(n_1093)
);

OAI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_925),
.A2(n_566),
.B1(n_588),
.B2(n_587),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_875),
.B(n_352),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_819),
.A2(n_653),
.B(n_688),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_808),
.A2(n_311),
.B1(n_340),
.B2(n_339),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_852),
.B(n_566),
.Y(n_1098)
);

AOI21x1_ASAP7_75t_L g1099 ( 
.A1(n_902),
.A2(n_528),
.B(n_524),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_894),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_855),
.B(n_566),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_792),
.A2(n_580),
.B(n_570),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_892),
.B(n_570),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_789),
.A2(n_653),
.B(n_688),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_795),
.A2(n_653),
.B(n_688),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_903),
.B(n_907),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_839),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_850),
.B(n_580),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_864),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_808),
.A2(n_304),
.B1(n_328),
.B2(n_323),
.Y(n_1110)
);

NOR2xp67_ASAP7_75t_L g1111 ( 
.A(n_826),
.B(n_277),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_797),
.A2(n_583),
.B(n_580),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_816),
.A2(n_914),
.B(n_920),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_830),
.B(n_256),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_826),
.A2(n_583),
.B(n_580),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_816),
.A2(n_653),
.B(n_688),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_786),
.A2(n_653),
.B(n_688),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_994),
.A2(n_921),
.B(n_838),
.C(n_786),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_1067),
.B(n_769),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1075),
.A2(n_838),
.B(n_926),
.C(n_915),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_968),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_989),
.Y(n_1122)
);

OR2x6_ASAP7_75t_L g1123 ( 
.A(n_980),
.B(n_866),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_995),
.B(n_866),
.Y(n_1124)
);

OAI21xp33_ASAP7_75t_L g1125 ( 
.A1(n_998),
.A2(n_361),
.B(n_358),
.Y(n_1125)
);

NAND2x1p5_ASAP7_75t_L g1126 ( 
.A(n_1088),
.B(n_926),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_SL g1127 ( 
.A(n_936),
.B(n_226),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_927),
.B(n_915),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_1041),
.Y(n_1129)
);

BUFx8_ASAP7_75t_SL g1130 ( 
.A(n_950),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_991),
.A2(n_904),
.B(n_834),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1076),
.B(n_866),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_949),
.B(n_362),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_969),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_L g1135 ( 
.A(n_1093),
.B(n_282),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_927),
.B(n_582),
.Y(n_1136)
);

NOR2xp67_ASAP7_75t_SL g1137 ( 
.A(n_1085),
.B(n_285),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_961),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_1027),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_939),
.A2(n_924),
.B(n_840),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1081),
.B(n_582),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1072),
.B(n_363),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1076),
.B(n_582),
.Y(n_1143)
);

OAI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_1030),
.A2(n_369),
.B(n_376),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_R g1145 ( 
.A(n_960),
.B(n_286),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1089),
.A2(n_308),
.B(n_396),
.C(n_382),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_990),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_1085),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1001),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1085),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_SL g1151 ( 
.A1(n_1071),
.A2(n_583),
.B(n_588),
.C(n_587),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1039),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1005),
.B(n_288),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_954),
.A2(n_688),
.B(n_653),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_958),
.B(n_364),
.Y(n_1155)
);

OR2x6_ASAP7_75t_L g1156 ( 
.A(n_980),
.B(n_295),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1003),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1005),
.B(n_294),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_934),
.A2(n_406),
.B(n_310),
.C(n_315),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_999),
.A2(n_528),
.B(n_587),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_935),
.A2(n_315),
.B(n_346),
.C(n_356),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_980),
.B(n_346),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1095),
.B(n_366),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_992),
.A2(n_356),
.B(n_357),
.C(n_360),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1069),
.A2(n_528),
.B(n_357),
.Y(n_1165)
);

INVx3_ASAP7_75t_SL g1166 ( 
.A(n_948),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1020),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_940),
.B(n_577),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1020),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1107),
.B(n_577),
.Y(n_1170)
);

NOR3xp33_ASAP7_75t_SL g1171 ( 
.A(n_955),
.B(n_413),
.C(n_410),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1109),
.B(n_296),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_965),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_976),
.A2(n_1032),
.B(n_1006),
.C(n_931),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1022),
.B(n_303),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_976),
.A2(n_409),
.B(n_360),
.C(n_406),
.Y(n_1176)
);

OAI22x1_ASAP7_75t_L g1177 ( 
.A1(n_1114),
.A2(n_380),
.B1(n_408),
.B2(n_404),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1092),
.B(n_367),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_928),
.B(n_312),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1022),
.B(n_314),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_956),
.A2(n_371),
.B(n_403),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1044),
.B(n_1055),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1026),
.B(n_316),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1007),
.B(n_331),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_927),
.B(n_332),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1037),
.A2(n_409),
.B(n_365),
.C(n_370),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1100),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_932),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_928),
.B(n_338),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_1088),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_R g1191 ( 
.A(n_943),
.B(n_342),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_996),
.A2(n_226),
.B1(n_298),
.B2(n_344),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_932),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_932),
.B(n_347),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_SL g1195 ( 
.A1(n_1036),
.A2(n_370),
.B(n_375),
.C(n_382),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_944),
.A2(n_945),
.B(n_947),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1038),
.B(n_385),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1070),
.B(n_350),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_943),
.Y(n_1199)
);

INVxp33_ASAP7_75t_SL g1200 ( 
.A(n_1043),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_967),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1052),
.A2(n_375),
.B(n_381),
.C(n_226),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_990),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_978),
.B(n_391),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_977),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_944),
.A2(n_373),
.B(n_399),
.Y(n_1206)
);

O2A1O1Ixp5_ASAP7_75t_SL g1207 ( 
.A1(n_1057),
.A2(n_996),
.B(n_957),
.C(n_981),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_987),
.Y(n_1208)
);

INVx5_ASAP7_75t_L g1209 ( 
.A(n_964),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_945),
.A2(n_377),
.B(n_397),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1070),
.B(n_394),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_R g1212 ( 
.A(n_1066),
.B(n_379),
.Y(n_1212)
);

NOR3xp33_ASAP7_75t_SL g1213 ( 
.A(n_974),
.B(n_402),
.C(n_401),
.Y(n_1213)
);

OR2x6_ASAP7_75t_SL g1214 ( 
.A(n_953),
.B(n_400),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_930),
.B(n_395),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_951),
.A2(n_140),
.B(n_83),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_962),
.B(n_392),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_938),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1004),
.B(n_17),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_938),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_933),
.B(n_195),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1091),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_966),
.A2(n_298),
.B(n_226),
.C(n_24),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_964),
.Y(n_1224)
);

AND2x4_ASAP7_75t_SL g1225 ( 
.A(n_967),
.B(n_298),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_967),
.Y(n_1226)
);

BUFx8_ASAP7_75t_SL g1227 ( 
.A(n_983),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_986),
.B(n_194),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1053),
.B(n_298),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1090),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1062),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1073),
.Y(n_1232)
);

NOR3xp33_ASAP7_75t_L g1233 ( 
.A(n_957),
.B(n_22),
.C(n_23),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_941),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_952),
.A2(n_970),
.B1(n_953),
.B2(n_963),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1079),
.Y(n_1236)
);

NOR2x1_ASAP7_75t_L g1237 ( 
.A(n_986),
.B(n_182),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1080),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1018),
.B(n_1068),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1074),
.B(n_178),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_952),
.A2(n_26),
.B1(n_28),
.B2(n_32),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_993),
.A2(n_163),
.B(n_159),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1018),
.B(n_1068),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_964),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_SL g1245 ( 
.A1(n_1010),
.A2(n_150),
.B(n_147),
.C(n_141),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1074),
.B(n_28),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1090),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1074),
.B(n_32),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1097),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1078),
.B(n_39),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_929),
.A2(n_136),
.B(n_132),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1106),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_973),
.A2(n_42),
.B(n_47),
.C(n_49),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1013),
.A2(n_946),
.B(n_942),
.C(n_1063),
.Y(n_1254)
);

OAI21xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1023),
.A2(n_47),
.B(n_49),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_SL g1256 ( 
.A(n_1017),
.B(n_129),
.Y(n_1256)
);

BUFx12f_ASAP7_75t_L g1257 ( 
.A(n_1015),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_937),
.A2(n_122),
.B(n_113),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1078),
.B(n_50),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1015),
.Y(n_1260)
);

NOR3xp33_ASAP7_75t_SL g1261 ( 
.A(n_1094),
.B(n_50),
.C(n_52),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1084),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1108),
.B(n_104),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1110),
.B(n_53),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1023),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_R g1266 ( 
.A(n_1015),
.B(n_103),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_979),
.A2(n_56),
.B(n_59),
.C(n_60),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1014),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_1268)
);

AOI222xp33_ASAP7_75t_L g1269 ( 
.A1(n_1111),
.A2(n_62),
.B1(n_65),
.B2(n_67),
.C1(n_71),
.C2(n_73),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1035),
.B(n_75),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_997),
.B(n_65),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_R g1272 ( 
.A(n_1035),
.B(n_85),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1045),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1011),
.B(n_71),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1035),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1016),
.B(n_73),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1084),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1025),
.A2(n_1031),
.B1(n_1009),
.B2(n_1024),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1077),
.A2(n_98),
.B(n_1009),
.C(n_1113),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1065),
.B(n_1042),
.Y(n_1280)
);

NAND3x1_ASAP7_75t_L g1281 ( 
.A(n_1133),
.B(n_1058),
.C(n_1019),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1174),
.A2(n_985),
.B(n_1046),
.C(n_1012),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1254),
.A2(n_1064),
.A3(n_1000),
.B(n_1002),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1134),
.B(n_1029),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1218),
.A2(n_1086),
.B1(n_1021),
.B2(n_1060),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1122),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1121),
.B(n_1086),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1142),
.B(n_1056),
.Y(n_1288)
);

INVx5_ASAP7_75t_L g1289 ( 
.A(n_1257),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1140),
.A2(n_959),
.B(n_971),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1196),
.A2(n_972),
.B(n_975),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1157),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1131),
.A2(n_988),
.B(n_1028),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1201),
.B(n_1065),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1139),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1143),
.A2(n_1008),
.B(n_1061),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1278),
.A2(n_1060),
.B(n_1047),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1161),
.A2(n_1083),
.A3(n_1087),
.B(n_1034),
.Y(n_1298)
);

AO32x2_ASAP7_75t_L g1299 ( 
.A1(n_1218),
.A2(n_1102),
.A3(n_1112),
.B1(n_1082),
.B2(n_1054),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1278),
.A2(n_1033),
.A3(n_1059),
.B(n_1051),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1149),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1182),
.B(n_1115),
.Y(n_1302)
);

NAND3x1_ASAP7_75t_L g1303 ( 
.A(n_1178),
.B(n_1115),
.C(n_1048),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1249),
.A2(n_1065),
.B1(n_1049),
.B2(n_1024),
.Y(n_1304)
);

AO22x2_ASAP7_75t_L g1305 ( 
.A1(n_1220),
.A2(n_1102),
.B1(n_984),
.B2(n_982),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1279),
.A2(n_982),
.B(n_984),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1252),
.B(n_1112),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1222),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1152),
.B(n_1215),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1138),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1235),
.A2(n_1050),
.B(n_1096),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1235),
.A2(n_1116),
.B(n_1098),
.Y(n_1312)
);

INVx5_ASAP7_75t_SL g1313 ( 
.A(n_1148),
.Y(n_1313)
);

INVx3_ASAP7_75t_SL g1314 ( 
.A(n_1166),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1119),
.B(n_1101),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1264),
.B(n_1103),
.C(n_1104),
.Y(n_1316)
);

BUFx5_ASAP7_75t_L g1317 ( 
.A(n_1273),
.Y(n_1317)
);

CKINVDCx6p67_ASAP7_75t_R g1318 ( 
.A(n_1167),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1215),
.B(n_1105),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_SL g1320 ( 
.A1(n_1163),
.A2(n_1117),
.B(n_1099),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1241),
.A2(n_1040),
.A3(n_1220),
.B(n_1265),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1168),
.A2(n_1165),
.B(n_1160),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1217),
.B(n_1262),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_1277),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1125),
.A2(n_1144),
.B(n_1202),
.C(n_1118),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1221),
.A2(n_1263),
.B(n_1256),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_1147),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1170),
.A2(n_1280),
.B(n_1228),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1207),
.A2(n_1189),
.B(n_1179),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1208),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1132),
.A2(n_1238),
.B1(n_1123),
.B2(n_1172),
.Y(n_1331)
);

AOI221xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1241),
.A2(n_1265),
.B1(n_1192),
.B2(n_1177),
.C(n_1159),
.Y(n_1332)
);

AOI21xp33_ASAP7_75t_L g1333 ( 
.A1(n_1197),
.A2(n_1155),
.B(n_1179),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_SL g1334 ( 
.A1(n_1132),
.A2(n_1221),
.B(n_1228),
.C(n_1240),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1263),
.A2(n_1154),
.B(n_1170),
.Y(n_1335)
);

AOI31xp67_ASAP7_75t_L g1336 ( 
.A1(n_1189),
.A2(n_1274),
.A3(n_1270),
.B(n_1198),
.Y(n_1336)
);

AOI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1233),
.A2(n_1124),
.B1(n_1269),
.B2(n_1259),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1188),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1214),
.B(n_1183),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1198),
.A2(n_1211),
.B(n_1184),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1251),
.A2(n_1258),
.B(n_1239),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1255),
.A2(n_1213),
.B(n_1271),
.C(n_1120),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1211),
.A2(n_1243),
.B(n_1172),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1206),
.A2(n_1210),
.B(n_1181),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1239),
.A2(n_1126),
.B(n_1216),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1126),
.A2(n_1242),
.B(n_1237),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1190),
.B(n_1193),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1141),
.B(n_1204),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1209),
.A2(n_1180),
.B(n_1175),
.Y(n_1349)
);

NAND3xp33_ASAP7_75t_L g1350 ( 
.A(n_1127),
.B(n_1261),
.C(n_1146),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1229),
.B(n_1136),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1209),
.A2(n_1158),
.B(n_1153),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1173),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1187),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1250),
.A2(n_1276),
.B(n_1219),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1200),
.B(n_1199),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1209),
.A2(n_1151),
.B(n_1123),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1205),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1234),
.A2(n_1164),
.B(n_1253),
.C(n_1176),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1231),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_SL g1361 ( 
.A(n_1145),
.B(n_1223),
.C(n_1191),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1128),
.B(n_1232),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1128),
.B(n_1236),
.Y(n_1363)
);

OR2x6_ASAP7_75t_L g1364 ( 
.A(n_1156),
.B(n_1162),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1147),
.A2(n_1203),
.B(n_1247),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1136),
.A2(n_1230),
.B(n_1135),
.Y(n_1366)
);

AO31x2_ASAP7_75t_L g1367 ( 
.A1(n_1234),
.A2(n_1246),
.A3(n_1248),
.B(n_1224),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1203),
.A2(n_1185),
.B(n_1194),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1209),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1171),
.B(n_1190),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1186),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1260),
.Y(n_1372)
);

O2A1O1Ixp5_ASAP7_75t_L g1373 ( 
.A1(n_1137),
.A2(n_1226),
.B(n_1224),
.C(n_1245),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1267),
.A2(n_1268),
.B(n_1195),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1156),
.B(n_1162),
.Y(n_1375)
);

BUFx10_ASAP7_75t_L g1376 ( 
.A(n_1129),
.Y(n_1376)
);

A2O1A1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1225),
.A2(n_1148),
.B(n_1150),
.C(n_1275),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1156),
.B(n_1162),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1123),
.A2(n_1272),
.B(n_1266),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1244),
.A2(n_1275),
.B(n_1148),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1227),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1150),
.B(n_1212),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1150),
.B(n_1169),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1130),
.B(n_994),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1133),
.A2(n_994),
.B(n_1067),
.C(n_998),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1133),
.B(n_994),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1207),
.A2(n_994),
.B(n_1067),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1133),
.B(n_994),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1133),
.A2(n_994),
.B(n_1067),
.C(n_998),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1264),
.A2(n_994),
.B1(n_787),
.B2(n_1067),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1142),
.B(n_805),
.Y(n_1391)
);

OAI22x1_ASAP7_75t_L g1392 ( 
.A1(n_1119),
.A2(n_994),
.B1(n_1067),
.B2(n_949),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1207),
.A2(n_994),
.B(n_1067),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1254),
.A2(n_1196),
.B(n_1161),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1207),
.A2(n_994),
.B(n_1067),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1140),
.A2(n_896),
.B(n_757),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1140),
.A2(n_896),
.B(n_757),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1165),
.A2(n_1160),
.B(n_1196),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1257),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1133),
.B(n_994),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1119),
.A2(n_994),
.B(n_787),
.C(n_1067),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1140),
.A2(n_896),
.B(n_757),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1140),
.A2(n_896),
.B(n_757),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1133),
.B(n_994),
.Y(n_1404)
);

NOR2xp67_ASAP7_75t_L g1405 ( 
.A(n_1147),
.B(n_1203),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1165),
.A2(n_1160),
.B(n_1196),
.Y(n_1406)
);

AO31x2_ASAP7_75t_L g1407 ( 
.A1(n_1254),
.A2(n_1161),
.A3(n_1278),
.B(n_1235),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1190),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1207),
.A2(n_994),
.B(n_1067),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1207),
.A2(n_994),
.B(n_1067),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1165),
.A2(n_1160),
.B(n_1196),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1140),
.A2(n_896),
.B(n_757),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1119),
.A2(n_994),
.B(n_787),
.C(n_1067),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1130),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1134),
.B(n_1081),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1207),
.A2(n_994),
.B(n_1067),
.Y(n_1416)
);

NAND3xp33_ASAP7_75t_L g1417 ( 
.A(n_1133),
.B(n_994),
.C(n_1067),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1140),
.A2(n_896),
.B(n_757),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1133),
.A2(n_994),
.B1(n_1067),
.B2(n_949),
.Y(n_1419)
);

AO31x2_ASAP7_75t_L g1420 ( 
.A1(n_1254),
.A2(n_1161),
.A3(n_1278),
.B(n_1235),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1122),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1133),
.B(n_994),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1165),
.A2(n_1160),
.B(n_1196),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1133),
.B(n_994),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1140),
.A2(n_896),
.B(n_757),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1165),
.A2(n_1160),
.B(n_1196),
.Y(n_1426)
);

CKINVDCx11_ASAP7_75t_R g1427 ( 
.A(n_1166),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1119),
.A2(n_994),
.B(n_787),
.C(n_1067),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1121),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1133),
.B(n_994),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1207),
.A2(n_994),
.B(n_1067),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1140),
.A2(n_896),
.B(n_757),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1207),
.A2(n_994),
.B(n_1067),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1134),
.B(n_1081),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_SL g1435 ( 
.A1(n_1278),
.A2(n_816),
.B(n_819),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1190),
.Y(n_1436)
);

AO31x2_ASAP7_75t_L g1437 ( 
.A1(n_1254),
.A2(n_1161),
.A3(n_1278),
.B(n_1235),
.Y(n_1437)
);

AO21x1_ASAP7_75t_L g1438 ( 
.A1(n_1241),
.A2(n_994),
.B(n_1218),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1257),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1140),
.A2(n_896),
.B(n_757),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1133),
.A2(n_994),
.B(n_1067),
.C(n_998),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1119),
.A2(n_994),
.B(n_787),
.C(n_1067),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1264),
.A2(n_994),
.B1(n_787),
.B2(n_1067),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1422),
.A2(n_1430),
.B1(n_1424),
.B2(n_1417),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1386),
.B(n_1388),
.Y(n_1445)
);

OAI22x1_ASAP7_75t_L g1446 ( 
.A1(n_1443),
.A2(n_1390),
.B1(n_1417),
.B2(n_1337),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1295),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1400),
.B(n_1404),
.Y(n_1448)
);

CKINVDCx11_ASAP7_75t_R g1449 ( 
.A(n_1376),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1427),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1314),
.Y(n_1451)
);

INVx6_ASAP7_75t_L g1452 ( 
.A(n_1289),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1390),
.A2(n_1443),
.B1(n_1419),
.B2(n_1337),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1317),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1438),
.A2(n_1333),
.B1(n_1392),
.B2(n_1350),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1385),
.A2(n_1389),
.B1(n_1441),
.B2(n_1339),
.Y(n_1456)
);

BUFx12f_ASAP7_75t_L g1457 ( 
.A(n_1376),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1317),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1286),
.Y(n_1459)
);

INVxp67_ASAP7_75t_SL g1460 ( 
.A(n_1324),
.Y(n_1460)
);

BUFx10_ASAP7_75t_L g1461 ( 
.A(n_1414),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1323),
.B(n_1391),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1361),
.A2(n_1331),
.B1(n_1351),
.B2(n_1384),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1317),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1381),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1292),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1350),
.A2(n_1409),
.B1(n_1410),
.B2(n_1387),
.Y(n_1467)
);

INVx6_ASAP7_75t_L g1468 ( 
.A(n_1289),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1393),
.A2(n_1433),
.B1(n_1431),
.B2(n_1395),
.Y(n_1469)
);

BUFx10_ASAP7_75t_L g1470 ( 
.A(n_1356),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1379),
.A2(n_1355),
.B1(n_1416),
.B2(n_1375),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1415),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1371),
.A2(n_1315),
.B1(n_1288),
.B2(n_1305),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1289),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1305),
.A2(n_1309),
.B1(n_1329),
.B2(n_1348),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1364),
.A2(n_1326),
.B1(n_1302),
.B2(n_1330),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1401),
.A2(n_1442),
.B1(n_1413),
.B2(n_1428),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1284),
.B(n_1434),
.Y(n_1478)
);

CKINVDCx11_ASAP7_75t_R g1479 ( 
.A(n_1318),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1364),
.A2(n_1378),
.B1(n_1370),
.B2(n_1382),
.Y(n_1480)
);

CKINVDCx11_ASAP7_75t_R g1481 ( 
.A(n_1399),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1308),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1372),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1429),
.Y(n_1484)
);

CKINVDCx11_ASAP7_75t_R g1485 ( 
.A(n_1399),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1369),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_1347),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1343),
.B(n_1332),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1325),
.A2(n_1342),
.B1(n_1287),
.B2(n_1362),
.Y(n_1489)
);

BUFx2_ASAP7_75t_SL g1490 ( 
.A(n_1399),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1363),
.A2(n_1281),
.B1(n_1304),
.B2(n_1338),
.Y(n_1491)
);

BUFx8_ASAP7_75t_SL g1492 ( 
.A(n_1439),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1394),
.A2(n_1360),
.B1(n_1353),
.B2(n_1358),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1408),
.A2(n_1436),
.B1(n_1307),
.B2(n_1377),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1310),
.Y(n_1495)
);

CKINVDCx11_ASAP7_75t_R g1496 ( 
.A(n_1439),
.Y(n_1496)
);

CKINVDCx12_ASAP7_75t_R g1497 ( 
.A(n_1285),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1439),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1383),
.Y(n_1499)
);

OAI21xp33_ASAP7_75t_L g1500 ( 
.A1(n_1359),
.A2(n_1319),
.B(n_1366),
.Y(n_1500)
);

BUFx10_ASAP7_75t_L g1501 ( 
.A(n_1383),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1394),
.A2(n_1374),
.B1(n_1297),
.B2(n_1306),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1294),
.Y(n_1503)
);

INVxp67_ASAP7_75t_SL g1504 ( 
.A(n_1405),
.Y(n_1504)
);

INVx4_ASAP7_75t_SL g1505 ( 
.A(n_1367),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_SL g1506 ( 
.A1(n_1285),
.A2(n_1344),
.B1(n_1368),
.B2(n_1313),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1407),
.B(n_1437),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1316),
.A2(n_1327),
.B1(n_1405),
.B2(n_1340),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1316),
.A2(n_1352),
.B1(n_1349),
.B2(n_1312),
.Y(n_1509)
);

CKINVDCx11_ASAP7_75t_R g1510 ( 
.A(n_1313),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_SL g1511 ( 
.A1(n_1346),
.A2(n_1357),
.B1(n_1345),
.B2(n_1341),
.Y(n_1511)
);

CKINVDCx11_ASAP7_75t_R g1512 ( 
.A(n_1336),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1321),
.A2(n_1311),
.B1(n_1437),
.B2(n_1407),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1328),
.A2(n_1335),
.B1(n_1420),
.B2(n_1437),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1380),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1435),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1367),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1303),
.Y(n_1518)
);

BUFx10_ASAP7_75t_L g1519 ( 
.A(n_1320),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1407),
.A2(n_1420),
.B1(n_1322),
.B2(n_1296),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_SL g1521 ( 
.A1(n_1321),
.A2(n_1420),
.B1(n_1365),
.B2(n_1334),
.Y(n_1521)
);

CKINVDCx11_ASAP7_75t_R g1522 ( 
.A(n_1373),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1300),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1322),
.A2(n_1321),
.B1(n_1291),
.B2(n_1290),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1396),
.A2(n_1403),
.B1(n_1432),
.B2(n_1425),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1282),
.A2(n_1402),
.B1(n_1418),
.B2(n_1412),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1300),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1298),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1398),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1283),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1293),
.A2(n_1440),
.B1(n_1397),
.B2(n_1406),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1298),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1283),
.Y(n_1533)
);

BUFx12f_ASAP7_75t_L g1534 ( 
.A(n_1283),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1411),
.Y(n_1535)
);

NAND2x1p5_ASAP7_75t_L g1536 ( 
.A(n_1426),
.B(n_1423),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1299),
.B(n_1422),
.Y(n_1537)
);

BUFx8_ASAP7_75t_SL g1538 ( 
.A(n_1414),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1324),
.Y(n_1539)
);

INVx6_ASAP7_75t_L g1540 ( 
.A(n_1289),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1422),
.A2(n_1430),
.B1(n_1424),
.B2(n_994),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1369),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1422),
.A2(n_1430),
.B1(n_1424),
.B2(n_994),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1544)
);

BUFx10_ASAP7_75t_L g1545 ( 
.A(n_1414),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1421),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1547)
);

BUFx2_ASAP7_75t_SL g1548 ( 
.A(n_1289),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1354),
.Y(n_1549)
);

CKINVDCx16_ASAP7_75t_R g1550 ( 
.A(n_1381),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1421),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1552)
);

BUFx8_ASAP7_75t_SL g1553 ( 
.A(n_1414),
.Y(n_1553)
);

CKINVDCx20_ASAP7_75t_R g1554 ( 
.A(n_1427),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1301),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1391),
.B(n_805),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1422),
.A2(n_1430),
.B1(n_1424),
.B2(n_994),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1427),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1562)
);

BUFx8_ASAP7_75t_L g1563 ( 
.A(n_1399),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_SL g1564 ( 
.A1(n_1422),
.A2(n_1430),
.B1(n_1424),
.B2(n_994),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1421),
.Y(n_1567)
);

OAI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1419),
.A2(n_994),
.B1(n_1424),
.B2(n_1422),
.Y(n_1568)
);

BUFx10_ASAP7_75t_L g1569 ( 
.A(n_1414),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1570)
);

INVx6_ASAP7_75t_L g1571 ( 
.A(n_1289),
.Y(n_1571)
);

BUFx8_ASAP7_75t_L g1572 ( 
.A(n_1399),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1354),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1421),
.Y(n_1575)
);

INVx8_ASAP7_75t_L g1576 ( 
.A(n_1289),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1301),
.Y(n_1577)
);

CKINVDCx11_ASAP7_75t_R g1578 ( 
.A(n_1376),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1369),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1580)
);

BUFx12f_ASAP7_75t_L g1581 ( 
.A(n_1427),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_SL g1582 ( 
.A1(n_1422),
.A2(n_1430),
.B1(n_1424),
.B2(n_994),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1430),
.B2(n_994),
.Y(n_1583)
);

BUFx12f_ASAP7_75t_L g1584 ( 
.A(n_1427),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1475),
.B(n_1467),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1552),
.A2(n_1570),
.B1(n_1566),
.B2(n_1561),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1533),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1517),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1507),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1472),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1536),
.A2(n_1531),
.B(n_1524),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1528),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1475),
.B(n_1537),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1445),
.B(n_1448),
.Y(n_1594)
);

OR2x6_ASAP7_75t_L g1595 ( 
.A(n_1534),
.B(n_1532),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1523),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1467),
.B(n_1469),
.Y(n_1597)
);

CKINVDCx6p67_ASAP7_75t_R g1598 ( 
.A(n_1479),
.Y(n_1598)
);

NOR2x1_ASAP7_75t_SL g1599 ( 
.A(n_1477),
.B(n_1534),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1515),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1456),
.A2(n_1500),
.B(n_1568),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1454),
.B(n_1458),
.Y(n_1602)
);

OAI21x1_ASAP7_75t_L g1603 ( 
.A1(n_1536),
.A2(n_1531),
.B(n_1524),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1505),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1508),
.A2(n_1488),
.B(n_1453),
.Y(n_1605)
);

OAI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1502),
.A2(n_1535),
.B(n_1526),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1473),
.B(n_1469),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1576),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1458),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1464),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1478),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1530),
.Y(n_1612)
);

AOI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1488),
.A2(n_1446),
.B(n_1535),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1527),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1455),
.B(n_1513),
.Y(n_1615)
);

AOI222xp33_ASAP7_75t_L g1616 ( 
.A1(n_1453),
.A2(n_1559),
.B1(n_1565),
.B2(n_1544),
.C1(n_1547),
.C2(n_1574),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1455),
.B(n_1546),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1502),
.A2(n_1520),
.B(n_1509),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1518),
.B(n_1462),
.Y(n_1619)
);

NAND3xp33_ASAP7_75t_L g1620 ( 
.A(n_1543),
.B(n_1557),
.C(n_1564),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1459),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1493),
.B(n_1466),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1493),
.B(n_1520),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1509),
.A2(n_1514),
.B(n_1476),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1582),
.A2(n_1561),
.B1(n_1566),
.B2(n_1580),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1460),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1484),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1541),
.A2(n_1570),
.B1(n_1583),
.B2(n_1580),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1538),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1482),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1514),
.A2(n_1476),
.B(n_1489),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1452),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1552),
.B(n_1560),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1539),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1529),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1483),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1521),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1491),
.A2(n_1494),
.B(n_1511),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1576),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1519),
.B(n_1506),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1551),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1560),
.A2(n_1583),
.B1(n_1444),
.B2(n_1562),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1555),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1463),
.B(n_1471),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1567),
.Y(n_1645)
);

AO21x2_ASAP7_75t_L g1646 ( 
.A1(n_1508),
.A2(n_1525),
.B(n_1512),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1575),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1576),
.Y(n_1648)
);

OR2x6_ASAP7_75t_L g1649 ( 
.A(n_1529),
.B(n_1480),
.Y(n_1649)
);

OA21x2_ASAP7_75t_L g1650 ( 
.A1(n_1495),
.A2(n_1444),
.B(n_1516),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1556),
.B(n_1577),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1452),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1497),
.Y(n_1653)
);

INVx4_ASAP7_75t_SL g1654 ( 
.A(n_1452),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1504),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1522),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1470),
.B(n_1499),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1487),
.B(n_1503),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1553),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1468),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1542),
.A2(n_1579),
.B(n_1540),
.Y(n_1661)
);

INVx4_ASAP7_75t_L g1662 ( 
.A(n_1468),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1447),
.Y(n_1663)
);

BUFx8_ASAP7_75t_SL g1664 ( 
.A(n_1581),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1447),
.B(n_1549),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1540),
.A2(n_1571),
.B(n_1486),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1540),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1501),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1501),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1571),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1510),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1474),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1548),
.Y(n_1673)
);

CKINVDCx11_ASAP7_75t_R g1674 ( 
.A(n_1554),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1573),
.B(n_1451),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1457),
.Y(n_1676)
);

OAI21x1_ASAP7_75t_L g1677 ( 
.A1(n_1490),
.A2(n_1563),
.B(n_1572),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1573),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1451),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1470),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1620),
.A2(n_1586),
.B1(n_1616),
.B2(n_1628),
.Y(n_1681)
);

BUFx3_ASAP7_75t_L g1682 ( 
.A(n_1671),
.Y(n_1682)
);

AO32x2_ASAP7_75t_L g1683 ( 
.A1(n_1679),
.A2(n_1449),
.A3(n_1578),
.B1(n_1563),
.B2(n_1572),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1611),
.B(n_1550),
.Y(n_1684)
);

OA21x2_ASAP7_75t_L g1685 ( 
.A1(n_1618),
.A2(n_1498),
.B(n_1450),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1594),
.B(n_1457),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1621),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1636),
.Y(n_1688)
);

AO32x2_ASAP7_75t_L g1689 ( 
.A1(n_1679),
.A2(n_1496),
.A3(n_1485),
.B1(n_1481),
.B2(n_1584),
.Y(n_1689)
);

AO21x1_ASAP7_75t_L g1690 ( 
.A1(n_1601),
.A2(n_1584),
.B(n_1581),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1620),
.A2(n_1558),
.B1(n_1465),
.B2(n_1492),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1625),
.A2(n_1569),
.B1(n_1461),
.B2(n_1545),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1628),
.A2(n_1569),
.B1(n_1461),
.B2(n_1545),
.Y(n_1693)
);

AO22x2_ASAP7_75t_L g1694 ( 
.A1(n_1644),
.A2(n_1597),
.B1(n_1585),
.B2(n_1607),
.Y(n_1694)
);

A2O1A1Ixp33_ASAP7_75t_L g1695 ( 
.A1(n_1605),
.A2(n_1644),
.B(n_1631),
.C(n_1597),
.Y(n_1695)
);

AOI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1642),
.A2(n_1585),
.B1(n_1633),
.B2(n_1615),
.C(n_1607),
.Y(n_1696)
);

INVxp33_ASAP7_75t_L g1697 ( 
.A(n_1651),
.Y(n_1697)
);

A2O1A1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1631),
.A2(n_1638),
.B(n_1656),
.C(n_1615),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1600),
.B(n_1627),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1626),
.Y(n_1700)
);

A2O1A1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1638),
.A2(n_1656),
.B(n_1624),
.C(n_1640),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1600),
.A2(n_1599),
.B(n_1646),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1590),
.B(n_1634),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1600),
.B(n_1643),
.Y(n_1704)
);

AND2x2_ASAP7_75t_SL g1705 ( 
.A(n_1650),
.B(n_1656),
.Y(n_1705)
);

OA21x2_ASAP7_75t_L g1706 ( 
.A1(n_1618),
.A2(n_1606),
.B(n_1624),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1619),
.A2(n_1593),
.B1(n_1653),
.B2(n_1650),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1653),
.A2(n_1646),
.B1(n_1617),
.B2(n_1619),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1637),
.A2(n_1680),
.B1(n_1622),
.B2(n_1657),
.C(n_1646),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1650),
.A2(n_1637),
.B1(n_1680),
.B2(n_1598),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1623),
.A2(n_1677),
.B(n_1678),
.C(n_1673),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_R g1712 ( 
.A(n_1629),
.B(n_1659),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1613),
.A2(n_1606),
.B(n_1650),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1665),
.B(n_1675),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_SL g1715 ( 
.A1(n_1599),
.A2(n_1649),
.B1(n_1676),
.B2(n_1671),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1655),
.Y(n_1716)
);

NOR2x1_ASAP7_75t_SL g1717 ( 
.A(n_1649),
.B(n_1595),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1658),
.Y(n_1718)
);

O2A1O1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1663),
.A2(n_1673),
.B(n_1675),
.C(n_1672),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1649),
.A2(n_1676),
.B1(n_1672),
.B2(n_1622),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1649),
.A2(n_1676),
.B1(n_1671),
.B2(n_1623),
.Y(n_1721)
);

NOR2x1_ASAP7_75t_SL g1722 ( 
.A(n_1649),
.B(n_1595),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1598),
.A2(n_1658),
.B1(n_1668),
.B2(n_1669),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1654),
.B(n_1602),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1655),
.A2(n_1676),
.B1(n_1671),
.B2(n_1672),
.Y(n_1725)
);

AO32x2_ASAP7_75t_L g1726 ( 
.A1(n_1632),
.A2(n_1662),
.A3(n_1589),
.B1(n_1614),
.B2(n_1612),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1609),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1630),
.B(n_1609),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1671),
.A2(n_1652),
.B1(n_1660),
.B2(n_1670),
.Y(n_1729)
);

NOR2xp67_ASAP7_75t_SL g1730 ( 
.A(n_1608),
.B(n_1639),
.Y(n_1730)
);

NOR2x1_ASAP7_75t_SL g1731 ( 
.A(n_1595),
.B(n_1589),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1645),
.B(n_1647),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1674),
.B(n_1664),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1677),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1588),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1666),
.A2(n_1661),
.B(n_1591),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1735),
.Y(n_1737)
);

AND2x2_ASAP7_75t_SL g1738 ( 
.A(n_1705),
.B(n_1604),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1687),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1700),
.B(n_1718),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1716),
.Y(n_1741)
);

INVxp67_ASAP7_75t_SL g1742 ( 
.A(n_1703),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1706),
.B(n_1603),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1726),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1736),
.B(n_1717),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1686),
.B(n_1670),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1734),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1727),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1706),
.B(n_1592),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1726),
.B(n_1592),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1697),
.B(n_1670),
.Y(n_1751)
);

OR2x2_ASAP7_75t_SL g1752 ( 
.A(n_1685),
.B(n_1647),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1736),
.B(n_1635),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1713),
.B(n_1596),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1708),
.B(n_1596),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1688),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1713),
.B(n_1587),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1732),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1728),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1722),
.B(n_1635),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1708),
.B(n_1587),
.Y(n_1761)
);

NOR2xp67_ASAP7_75t_L g1762 ( 
.A(n_1710),
.B(n_1641),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1681),
.A2(n_1595),
.B1(n_1670),
.B2(n_1667),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1685),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1681),
.A2(n_1694),
.B1(n_1696),
.B2(n_1690),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1719),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1707),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1707),
.Y(n_1768)
);

BUFx2_ASAP7_75t_SL g1769 ( 
.A(n_1682),
.Y(n_1769)
);

INVxp67_ASAP7_75t_SL g1770 ( 
.A(n_1710),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1744),
.B(n_1698),
.Y(n_1771)
);

NOR2x1_ASAP7_75t_L g1772 ( 
.A(n_1766),
.B(n_1702),
.Y(n_1772)
);

OAI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1765),
.A2(n_1695),
.B(n_1701),
.Y(n_1773)
);

INVx1_ASAP7_75t_SL g1774 ( 
.A(n_1756),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1737),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1756),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1770),
.A2(n_1709),
.B1(n_1693),
.B2(n_1691),
.C(n_1692),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1750),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1742),
.B(n_1694),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1737),
.Y(n_1780)
);

NOR3xp33_ASAP7_75t_L g1781 ( 
.A(n_1770),
.B(n_1693),
.C(n_1684),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1744),
.B(n_1731),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1760),
.B(n_1724),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1760),
.B(n_1753),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1747),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_L g1786 ( 
.A(n_1766),
.B(n_1711),
.C(n_1725),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1742),
.B(n_1714),
.Y(n_1787)
);

NAND4xp75_ASAP7_75t_L g1788 ( 
.A(n_1762),
.B(n_1733),
.C(n_1689),
.D(n_1725),
.Y(n_1788)
);

INVxp67_ASAP7_75t_L g1789 ( 
.A(n_1741),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1750),
.B(n_1761),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1737),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1762),
.A2(n_1721),
.B1(n_1720),
.B2(n_1715),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1747),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1739),
.Y(n_1794)
);

INVx5_ASAP7_75t_SL g1795 ( 
.A(n_1745),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1748),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1749),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1747),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1767),
.B(n_1610),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1748),
.Y(n_1800)
);

OAI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1755),
.A2(n_1729),
.B1(n_1723),
.B2(n_1704),
.Y(n_1801)
);

BUFx2_ASAP7_75t_L g1802 ( 
.A(n_1753),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1749),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1801),
.B(n_1738),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1775),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1778),
.B(n_1738),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1780),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1780),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1779),
.B(n_1767),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1778),
.B(n_1738),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1791),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1797),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1797),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1791),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1797),
.B(n_1768),
.Y(n_1815)
);

NAND2xp33_ASAP7_75t_L g1816 ( 
.A(n_1788),
.B(n_1712),
.Y(n_1816)
);

AND2x4_ASAP7_75t_SL g1817 ( 
.A(n_1783),
.B(n_1745),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1802),
.B(n_1768),
.Y(n_1818)
);

INVxp67_ASAP7_75t_SL g1819 ( 
.A(n_1779),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1785),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1802),
.B(n_1745),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1802),
.B(n_1745),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1790),
.B(n_1745),
.Y(n_1823)
);

OR2x6_ASAP7_75t_L g1824 ( 
.A(n_1788),
.B(n_1769),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1790),
.B(n_1754),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1789),
.B(n_1790),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1771),
.B(n_1754),
.Y(n_1827)
);

BUFx2_ASAP7_75t_L g1828 ( 
.A(n_1784),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1771),
.B(n_1754),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1771),
.B(n_1743),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1773),
.A2(n_1763),
.B1(n_1751),
.B2(n_1746),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1782),
.B(n_1743),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1794),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1789),
.B(n_1796),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1782),
.B(n_1753),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1803),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1796),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1782),
.B(n_1753),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1784),
.B(n_1753),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1794),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1800),
.Y(n_1841)
);

AOI221xp5_ASAP7_75t_L g1842 ( 
.A1(n_1773),
.A2(n_1755),
.B1(n_1740),
.B2(n_1758),
.C(n_1757),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1800),
.B(n_1759),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1837),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1820),
.B(n_1823),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1823),
.B(n_1806),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1837),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1820),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1823),
.B(n_1784),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1841),
.Y(n_1850)
);

NAND2xp67_ASAP7_75t_SL g1851 ( 
.A(n_1842),
.B(n_1806),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1809),
.B(n_1799),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1820),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1841),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1843),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1806),
.B(n_1784),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1842),
.B(n_1781),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1811),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1809),
.B(n_1781),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1826),
.B(n_1799),
.Y(n_1860)
);

BUFx2_ASAP7_75t_L g1861 ( 
.A(n_1820),
.Y(n_1861)
);

NAND2x1_ASAP7_75t_L g1862 ( 
.A(n_1810),
.B(n_1784),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1815),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1804),
.B(n_1787),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1810),
.B(n_1795),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1816),
.A2(n_1804),
.B1(n_1824),
.B2(n_1788),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1819),
.B(n_1787),
.Y(n_1867)
);

NAND2xp33_ASAP7_75t_L g1868 ( 
.A(n_1831),
.B(n_1772),
.Y(n_1868)
);

NAND2x1p5_ASAP7_75t_L g1869 ( 
.A(n_1810),
.B(n_1772),
.Y(n_1869)
);

NOR2x1p5_ASAP7_75t_SL g1870 ( 
.A(n_1812),
.B(n_1764),
.Y(n_1870)
);

OAI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1824),
.A2(n_1777),
.B1(n_1786),
.B2(n_1792),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1819),
.B(n_1801),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1843),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1811),
.Y(n_1874)
);

INVx2_ASAP7_75t_SL g1875 ( 
.A(n_1817),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1811),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1814),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1817),
.B(n_1795),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1817),
.B(n_1827),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1826),
.B(n_1799),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1814),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1834),
.Y(n_1882)
);

AND2x4_ASAP7_75t_SL g1883 ( 
.A(n_1824),
.B(n_1783),
.Y(n_1883)
);

OAI21xp33_ASAP7_75t_L g1884 ( 
.A1(n_1824),
.A2(n_1816),
.B(n_1786),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1814),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1833),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1833),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1817),
.B(n_1795),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1827),
.B(n_1795),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1827),
.B(n_1795),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1850),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1883),
.B(n_1829),
.Y(n_1892)
);

AO22x1_ASAP7_75t_L g1893 ( 
.A1(n_1871),
.A2(n_1792),
.B1(n_1824),
.B2(n_1699),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1844),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1883),
.B(n_1829),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_L g1896 ( 
.A(n_1868),
.B(n_1824),
.C(n_1777),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1861),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1889),
.B(n_1829),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1852),
.B(n_1834),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1864),
.B(n_1831),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1859),
.B(n_1830),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1858),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1889),
.B(n_1828),
.Y(n_1903)
);

NAND2x1_ASAP7_75t_L g1904 ( 
.A(n_1890),
.B(n_1824),
.Y(n_1904)
);

INVxp67_ASAP7_75t_L g1905 ( 
.A(n_1868),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1858),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1852),
.B(n_1815),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1890),
.B(n_1828),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1879),
.B(n_1828),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1877),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1884),
.A2(n_1740),
.B(n_1818),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1861),
.B(n_1821),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1879),
.B(n_1865),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1844),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1857),
.B(n_1830),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1865),
.B(n_1821),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1872),
.B(n_1783),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1882),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1846),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1867),
.B(n_1830),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1866),
.B(n_1825),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1855),
.B(n_1825),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_SL g1923 ( 
.A(n_1869),
.B(n_1774),
.Y(n_1923)
);

INVx2_ASAP7_75t_SL g1924 ( 
.A(n_1845),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1869),
.B(n_1795),
.Y(n_1925)
);

OR2x6_ASAP7_75t_L g1926 ( 
.A(n_1869),
.B(n_1608),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1860),
.B(n_1815),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1897),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1905),
.B(n_1846),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1900),
.B(n_1875),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1893),
.A2(n_1896),
.B(n_1923),
.Y(n_1931)
);

NOR3xp33_ASAP7_75t_L g1932 ( 
.A(n_1893),
.B(n_1853),
.C(n_1848),
.Y(n_1932)
);

AOI21xp33_ASAP7_75t_L g1933 ( 
.A1(n_1918),
.A2(n_1891),
.B(n_1914),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1913),
.A2(n_1845),
.B1(n_1888),
.B2(n_1878),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1901),
.B(n_1860),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1924),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1921),
.A2(n_1851),
.B(n_1862),
.Y(n_1937)
);

AOI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1913),
.A2(n_1845),
.B1(n_1888),
.B2(n_1878),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1924),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1902),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1915),
.B(n_1848),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1902),
.Y(n_1942)
);

AOI221xp5_ASAP7_75t_L g1943 ( 
.A1(n_1891),
.A2(n_1851),
.B1(n_1873),
.B2(n_1854),
.C(n_1847),
.Y(n_1943)
);

AOI221x1_ASAP7_75t_L g1944 ( 
.A1(n_1894),
.A2(n_1847),
.B1(n_1853),
.B2(n_1885),
.C(n_1881),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1912),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1906),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1919),
.B(n_1818),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1919),
.B(n_1911),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1916),
.B(n_1856),
.Y(n_1949)
);

OAI32xp33_ASAP7_75t_L g1950 ( 
.A1(n_1917),
.A2(n_1880),
.A3(n_1875),
.B1(n_1774),
.B2(n_1776),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1906),
.Y(n_1951)
);

OAI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1904),
.A2(n_1752),
.B1(n_1776),
.B2(n_1862),
.Y(n_1952)
);

OAI32xp33_ASAP7_75t_L g1953 ( 
.A1(n_1903),
.A2(n_1880),
.A3(n_1821),
.B1(n_1822),
.B2(n_1863),
.Y(n_1953)
);

AOI211xp5_ASAP7_75t_L g1954 ( 
.A1(n_1925),
.A2(n_1895),
.B(n_1892),
.C(n_1916),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1949),
.B(n_1898),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1928),
.B(n_1898),
.Y(n_1956)
);

INVxp67_ASAP7_75t_L g1957 ( 
.A(n_1930),
.Y(n_1957)
);

AOI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1931),
.A2(n_1904),
.B(n_1926),
.Y(n_1958)
);

OAI221xp5_ASAP7_75t_L g1959 ( 
.A1(n_1943),
.A2(n_1932),
.B1(n_1937),
.B2(n_1954),
.C(n_1933),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1940),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1945),
.B(n_1892),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1936),
.B(n_1912),
.Y(n_1962)
);

INVx2_ASAP7_75t_SL g1963 ( 
.A(n_1939),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1929),
.B(n_1912),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1942),
.Y(n_1965)
);

AOI221xp5_ASAP7_75t_SL g1966 ( 
.A1(n_1953),
.A2(n_1950),
.B1(n_1933),
.B2(n_1952),
.C(n_1948),
.Y(n_1966)
);

INVx2_ASAP7_75t_SL g1967 ( 
.A(n_1947),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1946),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1951),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1947),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_1948),
.Y(n_1971)
);

NOR3xp33_ASAP7_75t_L g1972 ( 
.A(n_1941),
.B(n_1899),
.C(n_1920),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1934),
.A2(n_1926),
.B1(n_1895),
.B2(n_1903),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1935),
.B(n_1908),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1938),
.B(n_1899),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1965),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1965),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1959),
.A2(n_1944),
.B(n_1952),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1963),
.Y(n_1979)
);

XNOR2x2_ASAP7_75t_L g1980 ( 
.A(n_1971),
.B(n_1910),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1963),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1961),
.Y(n_1982)
);

OAI211xp5_ASAP7_75t_L g1983 ( 
.A1(n_1966),
.A2(n_1908),
.B(n_1909),
.C(n_1910),
.Y(n_1983)
);

AOI211xp5_ASAP7_75t_L g1984 ( 
.A1(n_1958),
.A2(n_1909),
.B(n_1922),
.C(n_1927),
.Y(n_1984)
);

AOI21xp33_ASAP7_75t_L g1985 ( 
.A1(n_1957),
.A2(n_1975),
.B(n_1973),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1955),
.B(n_1926),
.Y(n_1986)
);

O2A1O1Ixp5_ASAP7_75t_L g1987 ( 
.A1(n_1956),
.A2(n_1927),
.B(n_1907),
.C(n_1863),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1968),
.Y(n_1988)
);

OAI211xp5_ASAP7_75t_L g1989 ( 
.A1(n_1978),
.A2(n_1962),
.B(n_1964),
.C(n_1975),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1980),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1986),
.B(n_1974),
.Y(n_1991)
);

NOR2x1_ASAP7_75t_L g1992 ( 
.A(n_1979),
.B(n_1968),
.Y(n_1992)
);

NAND3xp33_ASAP7_75t_L g1993 ( 
.A(n_1985),
.B(n_1970),
.C(n_1967),
.Y(n_1993)
);

NOR3xp33_ASAP7_75t_L g1994 ( 
.A(n_1982),
.B(n_1960),
.C(n_1969),
.Y(n_1994)
);

NAND3xp33_ASAP7_75t_L g1995 ( 
.A(n_1984),
.B(n_1967),
.C(n_1969),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1979),
.B(n_1961),
.Y(n_1996)
);

NOR3x1_ASAP7_75t_L g1997 ( 
.A(n_1983),
.B(n_1977),
.C(n_1976),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1981),
.B(n_1955),
.Y(n_1998)
);

INVxp67_ASAP7_75t_L g1999 ( 
.A(n_1981),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1986),
.B(n_1972),
.Y(n_2000)
);

AOI22xp33_ASAP7_75t_SL g2001 ( 
.A1(n_1990),
.A2(n_1980),
.B1(n_1988),
.B2(n_1926),
.Y(n_2001)
);

OAI211xp5_ASAP7_75t_L g2002 ( 
.A1(n_1989),
.A2(n_1988),
.B(n_1960),
.C(n_1987),
.Y(n_2002)
);

OAI221xp5_ASAP7_75t_L g2003 ( 
.A1(n_1993),
.A2(n_1907),
.B1(n_1793),
.B2(n_1785),
.C(n_1885),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1998),
.B(n_1856),
.Y(n_2004)
);

OAI211xp5_ASAP7_75t_L g2005 ( 
.A1(n_1995),
.A2(n_1689),
.B(n_1822),
.C(n_1793),
.Y(n_2005)
);

NAND5xp2_ASAP7_75t_L g2006 ( 
.A(n_1996),
.B(n_1689),
.C(n_1822),
.D(n_1683),
.E(n_1849),
.Y(n_2006)
);

NAND3xp33_ASAP7_75t_SL g2007 ( 
.A(n_2000),
.B(n_1793),
.C(n_1785),
.Y(n_2007)
);

AOI222xp33_ASAP7_75t_L g2008 ( 
.A1(n_1999),
.A2(n_1870),
.B1(n_1818),
.B2(n_1881),
.C1(n_1877),
.C2(n_1887),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_2001),
.B(n_1997),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_2002),
.B(n_1991),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_2005),
.A2(n_1994),
.B1(n_1992),
.B2(n_1849),
.Y(n_2011)
);

BUFx4f_ASAP7_75t_L g2012 ( 
.A(n_2007),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_2004),
.Y(n_2013)
);

AOI22xp33_ASAP7_75t_SL g2014 ( 
.A1(n_2003),
.A2(n_1798),
.B1(n_1769),
.B2(n_1839),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_2008),
.B(n_1798),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_2006),
.A2(n_1870),
.B(n_1876),
.C(n_1874),
.Y(n_2016)
);

NOR3xp33_ASAP7_75t_L g2017 ( 
.A(n_2010),
.B(n_1886),
.C(n_1662),
.Y(n_2017)
);

XOR2xp5_ASAP7_75t_L g2018 ( 
.A(n_2013),
.B(n_1639),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2011),
.Y(n_2019)
);

NAND4xp75_ASAP7_75t_L g2020 ( 
.A(n_2009),
.B(n_2015),
.C(n_2012),
.D(n_2014),
.Y(n_2020)
);

AOI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_2016),
.A2(n_1798),
.B1(n_1839),
.B2(n_1838),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2013),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_2022),
.A2(n_2018),
.B(n_2019),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_2020),
.B(n_1833),
.Y(n_2024)
);

AOI221x1_ASAP7_75t_L g2025 ( 
.A1(n_2017),
.A2(n_1840),
.B1(n_1808),
.B2(n_1807),
.C(n_1805),
.Y(n_2025)
);

AOI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_2023),
.A2(n_2021),
.B1(n_1798),
.B2(n_1838),
.C(n_1835),
.Y(n_2026)
);

INVxp67_ASAP7_75t_SL g2027 ( 
.A(n_2026),
.Y(n_2027)
);

XNOR2xp5_ASAP7_75t_L g2028 ( 
.A(n_2027),
.B(n_2024),
.Y(n_2028)
);

OAI22x1_ASAP7_75t_L g2029 ( 
.A1(n_2027),
.A2(n_2025),
.B1(n_1839),
.B2(n_1836),
.Y(n_2029)
);

OAI22x1_ASAP7_75t_L g2030 ( 
.A1(n_2028),
.A2(n_2029),
.B1(n_1839),
.B2(n_1813),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2028),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2030),
.Y(n_2032)
);

OAI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_2031),
.A2(n_1812),
.B1(n_1813),
.B2(n_1836),
.Y(n_2033)
);

OAI21xp5_ASAP7_75t_SL g2034 ( 
.A1(n_2032),
.A2(n_2033),
.B(n_1683),
.Y(n_2034)
);

AO21x2_ASAP7_75t_L g2035 ( 
.A1(n_2032),
.A2(n_1813),
.B(n_1812),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_2034),
.A2(n_1832),
.B1(n_1839),
.B2(n_1838),
.Y(n_2036)
);

XNOR2xp5_ASAP7_75t_L g2037 ( 
.A(n_2036),
.B(n_2035),
.Y(n_2037)
);

OAI221xp5_ASAP7_75t_R g2038 ( 
.A1(n_2037),
.A2(n_1683),
.B1(n_1812),
.B2(n_1836),
.C(n_1813),
.Y(n_2038)
);

AOI211xp5_ASAP7_75t_L g2039 ( 
.A1(n_2038),
.A2(n_1648),
.B(n_1639),
.C(n_1730),
.Y(n_2039)
);


endmodule