module fake_netlist_6_4729_n_1327 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_152, n_92, n_105, n_227, n_132, n_102, n_204, n_261, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_231, n_40, n_240, n_139, n_41, n_134, n_273, n_95, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1327);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_152;
input n_92;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_231;
input n_40;
input n_240;
input n_139;
input n_41;
input n_134;
input n_273;
input n_95;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1327;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_102),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_300),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_201),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_37),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_71),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_280),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_258),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_114),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_92),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_2),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_267),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_101),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_197),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_46),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_261),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_228),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_45),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_66),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_234),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_4),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_251),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_193),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_103),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_284),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_206),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_187),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_100),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_257),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_123),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_252),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_135),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_117),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_265),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_33),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_32),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_3),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_75),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_190),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_12),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_98),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_177),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_1),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_127),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_293),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_286),
.Y(n_352)
);

BUFx2_ASAP7_75t_SL g353 ( 
.A(n_175),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_297),
.Y(n_354)
);

BUFx10_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_242),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_270),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_124),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_137),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_178),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_26),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_167),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_179),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_287),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_171),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_168),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_196),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_11),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_43),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_166),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_115),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_106),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_140),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_285),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_269),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_40),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_80),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_141),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_276),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_172),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_181),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_108),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_63),
.Y(n_383)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_244),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_24),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_184),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_153),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_254),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_202),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_205),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_139),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_83),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_144),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_295),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_263),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_253),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_194),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_176),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_283),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_180),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_215),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_256),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_60),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_274),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_210),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_212),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_200),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_10),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_217),
.Y(n_409)
);

BUFx2_ASAP7_75t_SL g410 ( 
.A(n_240),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_268),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_36),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_305),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_110),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_220),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_216),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_0),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_281),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_162),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_74),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_224),
.Y(n_421)
);

INVxp33_ASAP7_75t_R g422 ( 
.A(n_70),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_105),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_249),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_159),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_243),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_129),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_64),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_271),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_161),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_147),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_68),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_236),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_301),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_5),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_226),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_204),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_7),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_119),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_298),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_42),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_111),
.Y(n_442)
);

HB1xp67_ASAP7_75t_SL g443 ( 
.A(n_90),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_50),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_6),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_288),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_61),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_282),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_62),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_128),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_255),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_14),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_118),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_73),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_109),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_78),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_59),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_302),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_165),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_221),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_227),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_207),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_170),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_86),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_136),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_259),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_65),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_279),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_272),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_7),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_246),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_143),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_88),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_85),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_275),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_28),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_307),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_248),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_121),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_211),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_294),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_93),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_21),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_29),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_182),
.B(n_266),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_8),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_304),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_315),
.B(n_31),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_388),
.B(n_0),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_343),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_384),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_312),
.B(n_337),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_317),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_315),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_355),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_323),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_327),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_411),
.B(n_1),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_315),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_385),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_346),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_315),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_384),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_384),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_416),
.Y(n_505)
);

AND2x2_ASAP7_75t_SL g506 ( 
.A(n_308),
.B(n_363),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_349),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_476),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_452),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_355),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_357),
.B(n_2),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_483),
.Y(n_512)
);

BUFx12f_ASAP7_75t_L g513 ( 
.A(n_361),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_416),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_329),
.A2(n_35),
.B(n_34),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_416),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_416),
.Y(n_517)
);

AOI22x1_ASAP7_75t_SL g518 ( 
.A1(n_435),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_412),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_484),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_486),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_432),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_377),
.B(n_6),
.Y(n_523)
);

OA21x2_ASAP7_75t_L g524 ( 
.A1(n_311),
.A2(n_8),
.B(n_9),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_408),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_432),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_432),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_438),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_384),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_364),
.A2(n_39),
.B(n_38),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_444),
.B(n_9),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_384),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_462),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_318),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_384),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_462),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_445),
.Y(n_538)
);

BUFx8_ASAP7_75t_L g539 ( 
.A(n_417),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_470),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_462),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_368),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_480),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_324),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_372),
.B(n_10),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_309),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_321),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_387),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_487),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_397),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_322),
.Y(n_552)
);

INVx6_ASAP7_75t_L g553 ( 
.A(n_365),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_310),
.Y(n_554)
);

BUFx8_ASAP7_75t_SL g555 ( 
.A(n_332),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_406),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_325),
.Y(n_557)
);

OA21x2_ASAP7_75t_L g558 ( 
.A1(n_326),
.A2(n_11),
.B(n_12),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_415),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_333),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_453),
.B(n_471),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_334),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_330),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_313),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_335),
.B(n_345),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_397),
.B(n_13),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_347),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_340),
.Y(n_568)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_485),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_314),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_443),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_443),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_362),
.A2(n_44),
.B(n_41),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_370),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_344),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_371),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_373),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_353),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_316),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_376),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_380),
.Y(n_581)
);

BUFx12f_ASAP7_75t_L g582 ( 
.A(n_319),
.Y(n_582)
);

BUFx12f_ASAP7_75t_L g583 ( 
.A(n_320),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_400),
.B(n_16),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_401),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_404),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_405),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_555),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_569),
.B(n_351),
.Y(n_589)
);

CKINVDCx16_ASAP7_75t_R g590 ( 
.A(n_496),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_548),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_557),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_547),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_544),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_535),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_569),
.B(n_407),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_494),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_570),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_582),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_583),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_519),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_552),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_494),
.Y(n_604)
);

AO21x2_ASAP7_75t_L g605 ( 
.A1(n_566),
.A2(n_414),
.B(n_413),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_579),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_553),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_549),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_568),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_513),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_554),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_549),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_549),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_511),
.B(n_427),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_578),
.B(n_418),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_R g616 ( 
.A(n_501),
.B(n_328),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_495),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_556),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_564),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_553),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_501),
.Y(n_621)
);

NAND2x1_ASAP7_75t_L g622 ( 
.A(n_488),
.B(n_424),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_578),
.B(n_538),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_494),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_556),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_572),
.B(n_331),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_507),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_556),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_R g629 ( 
.A(n_510),
.B(n_350),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_507),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_559),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_572),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_540),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_559),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_578),
.B(n_425),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_540),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_R g637 ( 
.A(n_506),
.B(n_375),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_493),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_497),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_559),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_572),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_525),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_490),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_528),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_R g645 ( 
.A(n_539),
.B(n_392),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_R g646 ( 
.A(n_550),
.B(n_336),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_539),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_500),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_543),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_R g650 ( 
.A(n_550),
.B(n_398),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_R g651 ( 
.A(n_571),
.B(n_402),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_542),
.Y(n_652)
);

NAND2x1_ASAP7_75t_L g653 ( 
.A(n_488),
.B(n_430),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_492),
.B(n_338),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_551),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_492),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_551),
.Y(n_657)
);

CKINVDCx6p67_ASAP7_75t_R g658 ( 
.A(n_498),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_580),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_576),
.Y(n_660)
);

CKINVDCx8_ASAP7_75t_R g661 ( 
.A(n_531),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_499),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_576),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_581),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_581),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_565),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_508),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_565),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_489),
.B(n_339),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_523),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_499),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_624),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_649),
.Y(n_673)
);

BUFx5_ASAP7_75t_L g674 ( 
.A(n_591),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_655),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_614),
.B(n_531),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_643),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_629),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_614),
.B(n_584),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_669),
.B(n_514),
.Y(n_680)
);

NOR2xp67_ASAP7_75t_L g681 ( 
.A(n_623),
.B(n_514),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_671),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_589),
.B(n_563),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_624),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_605),
.B(n_589),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_648),
.Y(n_686)
);

BUFx6f_ASAP7_75t_SL g687 ( 
.A(n_607),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_667),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_L g689 ( 
.A(n_596),
.B(n_561),
.C(n_546),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_605),
.B(n_514),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_671),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_598),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_604),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_597),
.B(n_516),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_662),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_624),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_603),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_597),
.B(n_611),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_608),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_654),
.A2(n_546),
.B1(n_584),
.B2(n_561),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_624),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_646),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_612),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_613),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_618),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_663),
.B(n_560),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_619),
.B(n_442),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_625),
.B(n_516),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_628),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_661),
.B(n_454),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_631),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_651),
.B(n_341),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_656),
.B(n_342),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_634),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_640),
.B(n_516),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_622),
.B(n_558),
.C(n_524),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_592),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_666),
.B(n_545),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_593),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_660),
.B(n_348),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_602),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_668),
.B(n_545),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_632),
.Y(n_723)
);

INVxp33_ASAP7_75t_L g724 ( 
.A(n_650),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_606),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_615),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_635),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_626),
.B(n_545),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_664),
.B(n_567),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_653),
.B(n_534),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_641),
.B(n_352),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_617),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_658),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_594),
.B(n_534),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_638),
.B(n_586),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_657),
.B(n_499),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_639),
.B(n_502),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_670),
.Y(n_738)
);

INVxp33_ASAP7_75t_SL g739 ( 
.A(n_645),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_642),
.B(n_509),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_644),
.B(n_502),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_607),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_621),
.B(n_354),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_627),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_630),
.B(n_502),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_633),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_636),
.Y(n_747)
);

INVxp33_ASAP7_75t_L g748 ( 
.A(n_637),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_652),
.B(n_520),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_647),
.B(n_599),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_659),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_665),
.B(n_574),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_600),
.B(n_356),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_601),
.B(n_587),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_610),
.B(n_505),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_620),
.B(n_491),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_590),
.B(n_503),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_609),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_595),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_588),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_616),
.B(n_505),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_614),
.A2(n_573),
.B(n_529),
.C(n_533),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_759),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_677),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_686),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_688),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_717),
.Y(n_767)
);

OR2x2_ASAP7_75t_SL g768 ( 
.A(n_733),
.B(n_422),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_676),
.B(n_488),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_673),
.B(n_512),
.Y(n_770)
);

AND2x6_ASAP7_75t_SL g771 ( 
.A(n_758),
.B(n_521),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_721),
.B(n_431),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_739),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_679),
.A2(n_524),
.B1(n_558),
.B2(n_410),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_740),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_734),
.B(n_358),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_687),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_685),
.A2(n_575),
.B1(n_437),
.B2(n_447),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_697),
.Y(n_779)
);

CKINVDCx11_ASAP7_75t_R g780 ( 
.A(n_675),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_719),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_692),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_693),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_675),
.B(n_587),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_695),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_734),
.B(n_359),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_702),
.A2(n_366),
.B1(n_367),
.B2(n_360),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_723),
.Y(n_788)
);

AO22x1_ASAP7_75t_L g789 ( 
.A1(n_761),
.A2(n_449),
.B1(n_451),
.B2(n_433),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_699),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_746),
.Y(n_791)
);

OAI22xp33_ASAP7_75t_L g792 ( 
.A1(n_683),
.A2(n_460),
.B1(n_464),
.B2(n_457),
.Y(n_792)
);

INVx4_ASAP7_75t_L g793 ( 
.A(n_746),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_703),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_746),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_704),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_727),
.B(n_726),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_689),
.B(n_468),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_716),
.A2(n_472),
.B1(n_474),
.B2(n_469),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_698),
.B(n_369),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_SL g801 ( 
.A(n_710),
.B(n_378),
.C(n_374),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_682),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_687),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_742),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_689),
.A2(n_381),
.B1(n_382),
.B2(n_379),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_700),
.B(n_475),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_749),
.B(n_383),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_706),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_729),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_L g810 ( 
.A(n_730),
.B(n_386),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_694),
.B(n_479),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_724),
.B(n_678),
.Y(n_812)
);

BUFx4f_ASAP7_75t_SL g813 ( 
.A(n_725),
.Y(n_813)
);

INVx5_ASAP7_75t_L g814 ( 
.A(n_672),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_674),
.B(n_481),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_R g816 ( 
.A(n_760),
.B(n_389),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_757),
.B(n_390),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_757),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_736),
.B(n_391),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_709),
.B(n_515),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_725),
.Y(n_821)
);

AND2x6_ASAP7_75t_L g822 ( 
.A(n_690),
.B(n_754),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_735),
.B(n_393),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_691),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_674),
.B(n_574),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_674),
.B(n_574),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_674),
.B(n_577),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_672),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_745),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_752),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_711),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_748),
.B(n_577),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_738),
.B(n_577),
.Y(n_833)
);

OR2x6_ASAP7_75t_L g834 ( 
.A(n_751),
.B(n_530),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_674),
.B(n_585),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_756),
.B(n_394),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_705),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_705),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_714),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_737),
.B(n_741),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_718),
.B(n_395),
.Y(n_841)
);

AOI221x1_ASAP7_75t_L g842 ( 
.A1(n_716),
.A2(n_504),
.B1(n_536),
.B2(n_585),
.C(n_541),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_732),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_701),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_672),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_684),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_756),
.Y(n_847)
);

NOR3xp33_ASAP7_75t_L g848 ( 
.A(n_707),
.B(n_399),
.C(n_396),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_680),
.B(n_585),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_762),
.A2(n_409),
.B(n_403),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_744),
.B(n_419),
.Y(n_851)
);

INVx5_ASAP7_75t_L g852 ( 
.A(n_684),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_684),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_712),
.A2(n_459),
.B1(n_421),
.B2(n_423),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_747),
.B(n_420),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_722),
.A2(n_428),
.B(n_426),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_769),
.A2(n_728),
.B(n_713),
.Y(n_857)
);

INVx5_ASAP7_75t_L g858 ( 
.A(n_795),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_795),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_830),
.B(n_743),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_821),
.B(n_720),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_764),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_799),
.A2(n_731),
.B1(n_429),
.B2(n_473),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_765),
.Y(n_864)
);

INVx6_ASAP7_75t_L g865 ( 
.A(n_793),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_840),
.B(n_755),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_766),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_779),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_800),
.A2(n_753),
.B(n_477),
.C(n_467),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_782),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_822),
.A2(n_681),
.B1(n_434),
.B2(n_466),
.Y(n_871)
);

NAND2xp33_ASAP7_75t_L g872 ( 
.A(n_822),
.B(n_696),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_774),
.A2(n_715),
.B(n_708),
.Y(n_873)
);

AOI21x1_ASAP7_75t_L g874 ( 
.A1(n_825),
.A2(n_681),
.B(n_696),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_838),
.A2(n_696),
.B(n_750),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_817),
.B(n_436),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_780),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_785),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_790),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_794),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_796),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_808),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_847),
.B(n_518),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_826),
.A2(n_541),
.B(n_517),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_827),
.A2(n_835),
.B(n_814),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_791),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_831),
.Y(n_887)
);

AO32x2_ASAP7_75t_L g888 ( 
.A1(n_778),
.A2(n_518),
.A3(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_767),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_840),
.B(n_439),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_784),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_806),
.A2(n_465),
.B1(n_441),
.B2(n_446),
.Y(n_892)
);

OA22x2_ASAP7_75t_L g893 ( 
.A1(n_818),
.A2(n_440),
.B1(n_448),
.B2(n_450),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_770),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_792),
.A2(n_455),
.B(n_456),
.C(n_458),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_814),
.A2(n_517),
.B(n_505),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_833),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_SL g898 ( 
.A1(n_850),
.A2(n_461),
.B(n_463),
.C(n_478),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_812),
.B(n_482),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_814),
.A2(n_852),
.B(n_797),
.Y(n_900)
);

XOR2x2_ASAP7_75t_L g901 ( 
.A(n_848),
.B(n_17),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_832),
.B(n_18),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_798),
.A2(n_541),
.B(n_537),
.C(n_532),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_852),
.A2(n_522),
.B(n_517),
.Y(n_904)
);

BUFx8_ASAP7_75t_L g905 ( 
.A(n_763),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_770),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_836),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_829),
.B(n_819),
.Y(n_908)
);

OA22x2_ASAP7_75t_L g909 ( 
.A1(n_809),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_909)
);

CKINVDCx8_ASAP7_75t_R g910 ( 
.A(n_771),
.Y(n_910)
);

NOR2xp67_ASAP7_75t_L g911 ( 
.A(n_773),
.B(n_47),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_788),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_843),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_822),
.A2(n_537),
.B1(n_532),
.B2(n_527),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_775),
.B(n_22),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_798),
.A2(n_537),
.B1(n_532),
.B2(n_527),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_837),
.B(n_522),
.Y(n_917)
);

CKINVDCx6p67_ASAP7_75t_R g918 ( 
.A(n_804),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_783),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_837),
.A2(n_527),
.B1(n_526),
.B2(n_522),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_852),
.A2(n_526),
.B(n_49),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_849),
.B(n_811),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_772),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_802),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_781),
.B(n_526),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_912),
.Y(n_926)
);

AO21x2_ASAP7_75t_L g927 ( 
.A1(n_898),
.A2(n_885),
.B(n_873),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_858),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_891),
.B(n_841),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_879),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_912),
.Y(n_931)
);

BUFx4_ASAP7_75t_SL g932 ( 
.A(n_859),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_902),
.B(n_841),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_858),
.B(n_828),
.Y(n_934)
);

OAI21x1_ASAP7_75t_L g935 ( 
.A1(n_874),
.A2(n_842),
.B(n_844),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_908),
.B(n_815),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_875),
.A2(n_853),
.B(n_846),
.Y(n_937)
);

AO21x2_ASAP7_75t_L g938 ( 
.A1(n_857),
.A2(n_856),
.B(n_823),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_862),
.Y(n_939)
);

OAI21x1_ASAP7_75t_SL g940 ( 
.A1(n_907),
.A2(n_824),
.B(n_839),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_900),
.A2(n_845),
.B(n_786),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_858),
.B(n_772),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_913),
.Y(n_943)
);

BUFx2_ASAP7_75t_SL g944 ( 
.A(n_886),
.Y(n_944)
);

INVx6_ASAP7_75t_L g945 ( 
.A(n_865),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_865),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_886),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_897),
.Y(n_948)
);

AO21x2_ASAP7_75t_L g949 ( 
.A1(n_914),
.A2(n_801),
.B(n_776),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_884),
.A2(n_855),
.B(n_851),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_925),
.A2(n_807),
.B(n_854),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_905),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_864),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_882),
.B(n_816),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_918),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_917),
.A2(n_787),
.B(n_834),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_867),
.Y(n_957)
);

BUFx4f_ASAP7_75t_L g958 ( 
.A(n_894),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_923),
.Y(n_959)
);

NAND2x1p5_ASAP7_75t_L g960 ( 
.A(n_868),
.B(n_828),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_906),
.B(n_828),
.Y(n_961)
);

AO21x2_ASAP7_75t_L g962 ( 
.A1(n_876),
.A2(n_820),
.B(n_810),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_881),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_899),
.B(n_813),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_919),
.A2(n_834),
.B(n_805),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_889),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_870),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_878),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_922),
.A2(n_887),
.B(n_880),
.Y(n_969)
);

BUFx12f_ASAP7_75t_L g970 ( 
.A(n_910),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_866),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_924),
.Y(n_972)
);

AOI22x1_ASAP7_75t_L g973 ( 
.A1(n_921),
.A2(n_820),
.B1(n_803),
.B2(n_777),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_877),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_911),
.B(n_48),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_883),
.B(n_789),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_890),
.A2(n_52),
.B(n_51),
.Y(n_977)
);

AO21x1_ASAP7_75t_L g978 ( 
.A1(n_872),
.A2(n_23),
.B(n_25),
.Y(n_978)
);

BUFx2_ASAP7_75t_SL g979 ( 
.A(n_909),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_861),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_915),
.A2(n_860),
.B(n_895),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_871),
.B(n_53),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_903),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_892),
.B(n_768),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_939),
.Y(n_985)
);

BUFx2_ASAP7_75t_R g986 ( 
.A(n_952),
.Y(n_986)
);

AOI21x1_ASAP7_75t_L g987 ( 
.A1(n_935),
.A2(n_937),
.B(n_956),
.Y(n_987)
);

BUFx8_ASAP7_75t_SL g988 ( 
.A(n_970),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_953),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_982),
.A2(n_901),
.B1(n_893),
.B2(n_863),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_963),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_930),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_966),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_963),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_957),
.Y(n_995)
);

OAI22xp33_ASAP7_75t_L g996 ( 
.A1(n_957),
.A2(n_888),
.B1(n_916),
.B2(n_920),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_966),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_982),
.A2(n_888),
.B1(n_869),
.B2(n_904),
.Y(n_998)
);

AOI21x1_ASAP7_75t_L g999 ( 
.A1(n_965),
.A2(n_896),
.B(n_55),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_932),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_934),
.Y(n_1001)
);

OAI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_971),
.A2(n_888),
.B1(n_26),
.B2(n_27),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_972),
.Y(n_1003)
);

NAND2x1p5_ASAP7_75t_L g1004 ( 
.A(n_958),
.B(n_54),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_967),
.Y(n_1005)
);

NAND2x1p5_ASAP7_75t_L g1006 ( 
.A(n_958),
.B(n_56),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_967),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_926),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_971),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_969),
.Y(n_1010)
);

AO21x2_ASAP7_75t_L g1011 ( 
.A1(n_927),
.A2(n_189),
.B(n_303),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_981),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_968),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_969),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_940),
.Y(n_1015)
);

CKINVDCx14_ASAP7_75t_R g1016 ( 
.A(n_952),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_968),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_960),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_964),
.A2(n_30),
.B1(n_58),
.B2(n_67),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_976),
.B(n_69),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_926),
.Y(n_1021)
);

BUFx12f_ASAP7_75t_L g1022 ( 
.A(n_943),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_960),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_961),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_961),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_945),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_983),
.Y(n_1027)
);

CKINVDCx11_ASAP7_75t_R g1028 ( 
.A(n_955),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_979),
.Y(n_1029)
);

OAI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_936),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_941),
.Y(n_1031)
);

NAND3xp33_ASAP7_75t_SL g1032 ( 
.A(n_981),
.B(n_79),
.C(n_81),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_927),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_933),
.B(n_82),
.Y(n_1034)
);

INVxp67_ASAP7_75t_L g1035 ( 
.A(n_944),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_950),
.A2(n_84),
.B(n_87),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_934),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_936),
.Y(n_1038)
);

AOI21x1_ASAP7_75t_L g1039 ( 
.A1(n_951),
.A2(n_306),
.B(n_91),
.Y(n_1039)
);

CKINVDCx16_ASAP7_75t_R g1040 ( 
.A(n_1016),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_991),
.B(n_980),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1020),
.B(n_929),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_990),
.A2(n_964),
.B1(n_954),
.B2(n_980),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_1008),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_988),
.Y(n_1045)
);

OAI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_1029),
.A2(n_980),
.B1(n_984),
.B2(n_955),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_992),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_990),
.B(n_942),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_992),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1038),
.B(n_946),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_985),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1038),
.B(n_946),
.Y(n_1052)
);

AO31x2_ASAP7_75t_L g1053 ( 
.A1(n_1033),
.A2(n_978),
.A3(n_962),
.B(n_938),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_989),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_1025),
.B(n_947),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_988),
.Y(n_1056)
);

CKINVDCx16_ASAP7_75t_R g1057 ( 
.A(n_1016),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1003),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_995),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_994),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_1026),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1034),
.B(n_942),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1027),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1012),
.A2(n_949),
.B1(n_975),
.B2(n_973),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_R g1065 ( 
.A(n_1000),
.B(n_945),
.Y(n_1065)
);

OR2x6_ASAP7_75t_L g1066 ( 
.A(n_1026),
.B(n_945),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_986),
.Y(n_1067)
);

AOI21xp33_ASAP7_75t_L g1068 ( 
.A1(n_998),
.A2(n_938),
.B(n_949),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_1028),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_998),
.A2(n_948),
.B1(n_959),
.B2(n_928),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1010),
.B(n_959),
.Y(n_1071)
);

AO31x2_ASAP7_75t_L g1072 ( 
.A1(n_1033),
.A2(n_962),
.A3(n_977),
.B(n_975),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_993),
.Y(n_1073)
);

CKINVDCx16_ASAP7_75t_R g1074 ( 
.A(n_1022),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1012),
.A2(n_1014),
.B(n_1032),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1024),
.B(n_959),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1027),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_993),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_1021),
.B(n_947),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_997),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1002),
.A2(n_974),
.B1(n_931),
.B2(n_928),
.Y(n_1081)
);

OR2x6_ASAP7_75t_L g1082 ( 
.A(n_1004),
.B(n_931),
.Y(n_1082)
);

OR2x2_ASAP7_75t_SL g1083 ( 
.A(n_1005),
.B(n_932),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_997),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_1035),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_1028),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_R g1087 ( 
.A(n_1037),
.B(n_89),
.Y(n_1087)
);

AND2x6_ASAP7_75t_L g1088 ( 
.A(n_1037),
.B(n_94),
.Y(n_1088)
);

NOR2x1p5_ASAP7_75t_L g1089 ( 
.A(n_1013),
.B(n_95),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_1001),
.Y(n_1090)
);

NAND2xp33_ASAP7_75t_R g1091 ( 
.A(n_1018),
.B(n_96),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1017),
.A2(n_97),
.B1(n_99),
.B2(n_104),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1007),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_1001),
.Y(n_1094)
);

CKINVDCx16_ASAP7_75t_R g1095 ( 
.A(n_1037),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1002),
.A2(n_107),
.B1(n_112),
.B2(n_113),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_1037),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_996),
.B(n_299),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1015),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1019),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_1053),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1053),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_1066),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_1079),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_1050),
.B(n_1015),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1048),
.B(n_1023),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1047),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1049),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1063),
.B(n_996),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1042),
.B(n_1004),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1062),
.B(n_1006),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_1052),
.B(n_1059),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_1082),
.B(n_1036),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_1082),
.B(n_1011),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1073),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1090),
.B(n_1011),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1078),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1079),
.B(n_999),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1051),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1094),
.B(n_1039),
.Y(n_1120)
);

INVxp33_ASAP7_75t_L g1121 ( 
.A(n_1041),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1084),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_1066),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1077),
.B(n_1031),
.Y(n_1124)
);

NAND2xp33_ASAP7_75t_SL g1125 ( 
.A(n_1087),
.B(n_1009),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1060),
.B(n_987),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1053),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1099),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1054),
.B(n_1006),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1058),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1093),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1080),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1055),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_1072),
.Y(n_1134)
);

INVx6_ASAP7_75t_L g1135 ( 
.A(n_1095),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1097),
.B(n_1031),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1043),
.B(n_1030),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_1065),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_1071),
.B(n_1030),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1076),
.B(n_116),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1070),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_1044),
.B(n_120),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1055),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1068),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1085),
.B(n_122),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1061),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1072),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1098),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1083),
.B(n_125),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_1046),
.B(n_126),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1081),
.B(n_130),
.Y(n_1151)
);

AOI211xp5_ASAP7_75t_SL g1152 ( 
.A1(n_1096),
.A2(n_131),
.B(n_132),
.C(n_133),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1088),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1088),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1075),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1064),
.B(n_134),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1088),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1100),
.B(n_138),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1112),
.B(n_1040),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1126),
.B(n_1089),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1155),
.B(n_1057),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1126),
.B(n_1119),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1130),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_1121),
.B(n_1074),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1131),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1104),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1148),
.B(n_1069),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1105),
.B(n_1086),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1106),
.B(n_1067),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1128),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1109),
.B(n_1092),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1110),
.B(n_142),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1137),
.B(n_1091),
.C(n_1056),
.Y(n_1173)
);

NOR3xp33_ASAP7_75t_L g1174 ( 
.A(n_1125),
.B(n_1045),
.C(n_146),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1143),
.B(n_296),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1111),
.B(n_145),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1114),
.B(n_1157),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1135),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1128),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1114),
.B(n_291),
.Y(n_1180)
);

OAI221xp5_ASAP7_75t_SL g1181 ( 
.A1(n_1137),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.C(n_151),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1132),
.B(n_152),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_1109),
.B(n_154),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1124),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1107),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1125),
.B(n_155),
.C(n_156),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1124),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_L g1188 ( 
.A(n_1120),
.B(n_157),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1108),
.Y(n_1189)
);

NOR2xp67_ASAP7_75t_L g1190 ( 
.A(n_1120),
.B(n_158),
.Y(n_1190)
);

NOR2xp67_ASAP7_75t_L g1191 ( 
.A(n_1118),
.B(n_160),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1115),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1135),
.B(n_290),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1117),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1135),
.B(n_163),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1144),
.B(n_164),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1133),
.B(n_169),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1144),
.B(n_173),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1133),
.B(n_174),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1122),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1141),
.B(n_1139),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1133),
.B(n_289),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1162),
.B(n_1177),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1163),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1165),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1162),
.B(n_1101),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1170),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1201),
.B(n_1116),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1179),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1177),
.B(n_1103),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1189),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1192),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1194),
.B(n_1116),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1184),
.B(n_1101),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1200),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1185),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1187),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1164),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1159),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1160),
.B(n_1118),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1161),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1160),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1178),
.B(n_1153),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1196),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1168),
.B(n_1154),
.Y(n_1225)
);

INVx1_ASAP7_75t_SL g1226 ( 
.A(n_1166),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1171),
.B(n_1129),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1198),
.B(n_1102),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_1169),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1182),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1180),
.B(n_1102),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1183),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1209),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1206),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1204),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1209),
.B(n_1127),
.Y(n_1236)
);

OAI21xp33_ASAP7_75t_L g1237 ( 
.A1(n_1232),
.A2(n_1181),
.B(n_1186),
.Y(n_1237)
);

XOR2x2_ASAP7_75t_L g1238 ( 
.A(n_1226),
.B(n_1173),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1208),
.B(n_1127),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1220),
.B(n_1180),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1214),
.B(n_1134),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1204),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1214),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1232),
.B(n_1171),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1227),
.B(n_1167),
.Y(n_1245)
);

AND2x2_ASAP7_75t_SL g1246 ( 
.A(n_1220),
.B(n_1174),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_1205),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1218),
.B(n_1134),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1217),
.B(n_1147),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1221),
.B(n_1173),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1203),
.B(n_1138),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1203),
.B(n_1172),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1229),
.A2(n_1186),
.B1(n_1151),
.B2(n_1156),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1237),
.A2(n_1220),
.B1(n_1219),
.B2(n_1230),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1246),
.A2(n_1156),
.B(n_1152),
.Y(n_1255)
);

OAI21xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1250),
.A2(n_1244),
.B(n_1247),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1238),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1245),
.A2(n_1158),
.B(n_1152),
.C(n_1230),
.Y(n_1258)
);

AO22x1_ASAP7_75t_L g1259 ( 
.A1(n_1240),
.A2(n_1222),
.B1(n_1224),
.B2(n_1223),
.Y(n_1259)
);

OAI21xp33_ASAP7_75t_L g1260 ( 
.A1(n_1253),
.A2(n_1213),
.B(n_1228),
.Y(n_1260)
);

NOR3xp33_ASAP7_75t_L g1261 ( 
.A(n_1236),
.B(n_1158),
.C(n_1149),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1240),
.A2(n_1222),
.B1(n_1191),
.B2(n_1190),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1251),
.A2(n_1222),
.B1(n_1225),
.B2(n_1210),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1234),
.A2(n_1150),
.B(n_1188),
.C(n_1190),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1254),
.B(n_1239),
.Y(n_1265)
);

AOI211xp5_ASAP7_75t_L g1266 ( 
.A1(n_1257),
.A2(n_1188),
.B(n_1191),
.C(n_1145),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1259),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1260),
.B(n_1234),
.Y(n_1268)
);

AOI321xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1256),
.A2(n_1243),
.A3(n_1233),
.B1(n_1236),
.B2(n_1241),
.C(n_1248),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1261),
.B(n_1263),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1262),
.B(n_1252),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1264),
.B(n_1206),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1258),
.B(n_1242),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1255),
.B(n_1235),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1259),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1254),
.B(n_1231),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1259),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1259),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1270),
.A2(n_1273),
.B(n_1274),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1268),
.A2(n_1249),
.B(n_1215),
.Y(n_1280)
);

NAND3xp33_ASAP7_75t_L g1281 ( 
.A(n_1266),
.B(n_1212),
.C(n_1211),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1266),
.A2(n_1249),
.B(n_1207),
.Y(n_1282)
);

AOI21xp33_ASAP7_75t_L g1283 ( 
.A1(n_1267),
.A2(n_1142),
.B(n_1193),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1265),
.B(n_1275),
.Y(n_1284)
);

NAND3xp33_ASAP7_75t_SL g1285 ( 
.A(n_1269),
.B(n_1278),
.C(n_1277),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1271),
.B(n_1231),
.Y(n_1286)
);

AOI21xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1284),
.A2(n_1269),
.B(n_1272),
.Y(n_1287)
);

O2A1O1Ixp5_ASAP7_75t_L g1288 ( 
.A1(n_1279),
.A2(n_1276),
.B(n_1216),
.C(n_1205),
.Y(n_1288)
);

AOI32xp33_ASAP7_75t_L g1289 ( 
.A1(n_1285),
.A2(n_1195),
.A3(n_1176),
.B1(n_1199),
.B2(n_1197),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1286),
.Y(n_1290)
);

NOR2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1281),
.B(n_1123),
.Y(n_1291)
);

OAI211xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1283),
.A2(n_1280),
.B(n_1282),
.C(n_1146),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1287),
.A2(n_1289),
.B1(n_1291),
.B2(n_1290),
.Y(n_1293)
);

NAND2xp33_ASAP7_75t_R g1294 ( 
.A(n_1288),
.B(n_1202),
.Y(n_1294)
);

AOI211xp5_ASAP7_75t_L g1295 ( 
.A1(n_1292),
.A2(n_1123),
.B(n_1140),
.C(n_1175),
.Y(n_1295)
);

NOR3xp33_ASAP7_75t_L g1296 ( 
.A(n_1287),
.B(n_1113),
.C(n_1136),
.Y(n_1296)
);

INVxp33_ASAP7_75t_SL g1297 ( 
.A(n_1293),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1296),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1294),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1295),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1293),
.B(n_183),
.Y(n_1301)
);

NOR3xp33_ASAP7_75t_L g1302 ( 
.A(n_1301),
.B(n_185),
.C(n_186),
.Y(n_1302)
);

AOI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1297),
.A2(n_188),
.B1(n_191),
.B2(n_192),
.C(n_195),
.Y(n_1303)
);

NAND4xp75_ASAP7_75t_L g1304 ( 
.A(n_1300),
.B(n_198),
.C(n_199),
.D(n_203),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1299),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1305),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1304),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1302),
.Y(n_1308)
);

OAI22x1_ASAP7_75t_L g1309 ( 
.A1(n_1307),
.A2(n_1298),
.B1(n_1303),
.B2(n_213),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1306),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1306),
.B(n_208),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1308),
.Y(n_1312)
);

AOI31xp33_ASAP7_75t_L g1313 ( 
.A1(n_1310),
.A2(n_209),
.A3(n_214),
.B(n_218),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1312),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1311),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1309),
.B(n_225),
.Y(n_1316)
);

NAND2xp33_ASAP7_75t_R g1317 ( 
.A(n_1316),
.B(n_229),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1315),
.B(n_230),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1313),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_SL g1320 ( 
.A1(n_1319),
.A2(n_1314),
.B1(n_237),
.B2(n_238),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1318),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1320),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1321),
.A2(n_1317),
.B(n_239),
.Y(n_1323)
);

AOI222xp33_ASAP7_75t_L g1324 ( 
.A1(n_1322),
.A2(n_235),
.B1(n_241),
.B2(n_245),
.C1(n_247),
.C2(n_250),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1323),
.A2(n_260),
.B1(n_262),
.B2(n_264),
.Y(n_1325)
);

OR2x6_ASAP7_75t_L g1326 ( 
.A(n_1325),
.B(n_273),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1326),
.A2(n_1324),
.B1(n_277),
.B2(n_278),
.Y(n_1327)
);


endmodule