module real_jpeg_6061_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_1),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_1),
.A2(n_58),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_1),
.A2(n_58),
.B1(n_278),
.B2(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_2),
.A2(n_126),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_2),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_2),
.A2(n_137),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_3),
.A2(n_163),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_3),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_4),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_4),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_4),
.A2(n_189),
.B(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_4),
.B(n_247),
.C(n_249),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_L g251 ( 
.A1(n_4),
.A2(n_127),
.B1(n_151),
.B2(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_4),
.B(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_4),
.A2(n_76),
.B1(n_171),
.B2(n_299),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_5),
.A2(n_49),
.B1(n_220),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_5),
.A2(n_49),
.B1(n_127),
.B2(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_5),
.A2(n_49),
.B1(n_288),
.B2(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_6),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_64),
.B1(n_69),
.B2(n_70),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_8),
.A2(n_121),
.B1(n_122),
.B2(n_127),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_8),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_8),
.A2(n_50),
.B1(n_121),
.B2(n_206),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_8),
.A2(n_121),
.B1(n_272),
.B2(n_275),
.Y(n_271)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_10),
.Y(n_197)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_10),
.Y(n_282)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_11),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_11),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_11),
.Y(n_227)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_11),
.Y(n_231)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_13),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_13),
.Y(n_191)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_13),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_13),
.Y(n_225)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_13),
.Y(n_228)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_13),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_14),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_14),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_14),
.A2(n_87),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_15),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_15),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_239),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_237),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_174),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_19),
.B(n_174),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_99),
.C(n_138),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_20),
.A2(n_21),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_60),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_22),
.B(n_61),
.C(n_98),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_47),
.B2(n_57),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_23),
.A2(n_25),
.B1(n_57),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_24),
.A2(n_48),
.B1(n_263),
.B2(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_25),
.Y(n_263)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_26),
.Y(n_216)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_27),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_27),
.Y(n_253)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_29),
.Y(n_157)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_31),
.Y(n_214)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_32),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_32),
.Y(n_146)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_32),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_42),
.B2(n_45),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_37),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_38),
.Y(n_143)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_40),
.Y(n_149)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_43),
.A2(n_55),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_91),
.B2(n_98),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_74),
.B(n_75),
.Y(n_62)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_63),
.Y(n_193)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_73),
.Y(n_278)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_73),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_83),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_76),
.A2(n_161),
.B(n_169),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_76),
.A2(n_193),
.B1(n_194),
.B2(n_198),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_76),
.A2(n_271),
.B(n_279),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_76),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_76),
.A2(n_171),
.B1(n_287),
.B2(n_299),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_82),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_82),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_85),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_93),
.A2(n_218),
.B1(n_223),
.B2(n_232),
.Y(n_217)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_94),
.B(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_97),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_99),
.A2(n_138),
.B1(n_139),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_99),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_119),
.B(n_130),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_100),
.A2(n_134),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_101),
.A2(n_133),
.B1(n_251),
.B2(n_254),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_101),
.A2(n_133),
.B1(n_254),
.B2(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_101),
.A2(n_120),
.B1(n_133),
.B2(n_265),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_112),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_111),
.Y(n_102)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_103),
.Y(n_245)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_110),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_111),
.Y(n_266)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_112)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_132),
.B(n_151),
.Y(n_297)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_133),
.B(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_160),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_140),
.B(n_160),
.Y(n_319)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_144),
.A3(n_147),
.B1(n_150),
.B2(n_155),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_SL g322 ( 
.A1(n_142),
.A2(n_150),
.B(n_151),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_151),
.B(n_306),
.Y(n_305)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_161),
.Y(n_280)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_167),
.Y(n_301)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_168),
.Y(n_274)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_168),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_202),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_201),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_192),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_180),
.A3(n_182),
.B1(n_184),
.B2(n_188),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_199),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_202),
.Y(n_332)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_210),
.CI(n_217),
.CON(n_202),
.SN(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_SL g207 ( 
.A(n_208),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_325),
.B(n_331),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_316),
.B(n_324),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_283),
.B(n_315),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_259),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_243),
.B(n_259),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_250),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_250),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_270),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_269),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_261),
.B(n_269),
.C(n_270),
.Y(n_317)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_264),
.Y(n_269)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_295),
.B(n_314),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_294),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_294),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_302),
.B(n_313),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_297),
.B(n_298),
.Y(n_313)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_309),
.Y(n_304)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_318),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_321),
.C(n_323),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);


endmodule