module fake_jpeg_30317_n_140 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_65),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_21),
.B1(n_39),
.B2(n_38),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_46),
.B1(n_57),
.B2(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_0),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_72),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_58),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_52),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_50),
.B1(n_52),
.B2(n_43),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_43),
.B1(n_54),
.B2(n_51),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_93),
.Y(n_111)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_76),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_97),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_87),
.B(n_91),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_55),
.B1(n_44),
.B2(n_45),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_19),
.C(n_37),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_3),
.C(n_5),
.Y(n_99)
);

OA21x2_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_1),
.B(n_2),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_95),
.B(n_82),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_80),
.B1(n_5),
.B2(n_6),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_100),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_94),
.Y(n_100)
);

NOR2x1_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_7),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_40),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_109),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_106),
.B(n_32),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_12),
.C(n_14),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_16),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_17),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_24),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_26),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_29),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_114),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_30),
.B(n_31),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_120),
.B(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_119),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_33),
.B(n_35),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_108),
.C(n_112),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_114),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_116),
.C(n_120),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_130),
.Y(n_134)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_134),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_135),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_126),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_122),
.C(n_129),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_123),
.Y(n_140)
);


endmodule