module fake_jpeg_13805_n_160 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_7),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_15),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_31),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_40),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_0),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_77),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_58),
.B1(n_59),
.B2(n_54),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_80),
.Y(n_96)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_1),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_19),
.B1(n_47),
.B2(n_44),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_69),
.C(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_48),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_3),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_88),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_87),
.B(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_66),
.Y(n_88)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_95),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_51),
.B(n_49),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_52),
.CI(n_55),
.CON(n_107),
.SN(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_6),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_64),
.B1(n_53),
.B2(n_71),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_110),
.B1(n_113),
.B2(n_12),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_53),
.B1(n_51),
.B2(n_64),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_11),
.B(n_12),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_55),
.B(n_52),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_101),
.C(n_15),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_65),
.C(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_17),
.Y(n_134)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_61),
.B1(n_8),
.B2(n_9),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_14),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_110)
);

AOI32xp33_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_20),
.A3(n_39),
.B1(n_33),
.B2(n_30),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_SL g127 ( 
.A(n_112),
.B(n_21),
.C(n_27),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_85),
.B1(n_93),
.B2(n_86),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_13),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_10),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_116),
.B(n_41),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_125),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_10),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_121),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_11),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_134),
.B1(n_136),
.B2(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_128),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_13),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_130),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_16),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_24),
.C(n_26),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_135),
.C(n_104),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_99),
.C(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_17),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_144),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_124),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.C(n_144),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_135),
.A2(n_28),
.B1(n_103),
.B2(n_123),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_146),
.B1(n_133),
.B2(n_127),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_130),
.B1(n_129),
.B2(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_148),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_149),
.A2(n_151),
.B(n_139),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_125),
.B(n_146),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_138),
.B(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_153),
.B(n_155),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_151),
.C(n_152),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_150),
.C(n_140),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_154),
.Y(n_159)
);

HAxp5_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_143),
.CON(n_160),
.SN(n_160)
);


endmodule