module fake_jpeg_5672_n_326 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_40),
.Y(n_44)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_2),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_56),
.Y(n_73)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_20),
.B(n_2),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_68),
.Y(n_95)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_50),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_19),
.B(n_3),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_63),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_21),
.B(n_3),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_66),
.Y(n_86)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_62),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_67),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_3),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_4),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_36),
.B1(n_29),
.B2(n_32),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_69),
.A2(n_78),
.B1(n_83),
.B2(n_111),
.Y(n_123)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_70),
.B(n_71),
.Y(n_148)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_72),
.B(n_74),
.Y(n_149)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_75),
.B(n_81),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_41),
.B1(n_38),
.B2(n_43),
.Y(n_78)
);

OR2x4_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_39),
.Y(n_79)
);

NOR2x1_ASAP7_75t_SL g147 ( 
.A(n_79),
.B(n_112),
.Y(n_147)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_37),
.B1(n_36),
.B2(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_84),
.B(n_107),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_41),
.B1(n_37),
.B2(n_26),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_69),
.B1(n_79),
.B2(n_31),
.Y(n_126)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_93),
.B(n_101),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_61),
.A2(n_23),
.B1(n_26),
.B2(n_22),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_62),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

BUFx2_ASAP7_75t_R g105 ( 
.A(n_58),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_66),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_34),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_57),
.A2(n_23),
.B1(n_30),
.B2(n_27),
.Y(n_111)
);

NAND2xp33_ASAP7_75t_SL g112 ( 
.A(n_58),
.B(n_27),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_39),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_125),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_121),
.B(n_127),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_73),
.B(n_52),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_104),
.B1(n_98),
.B2(n_70),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_39),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_128),
.B1(n_130),
.B2(n_145),
.Y(n_154)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_87),
.B1(n_78),
.B2(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_58),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_141),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_69),
.A2(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_112),
.A2(n_33),
.B(n_32),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_140),
.C(n_72),
.Y(n_165)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_76),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_82),
.B(n_4),
.Y(n_137)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_46),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_5),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_29),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_140),
.Y(n_158)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_83),
.A2(n_29),
.B1(n_28),
.B2(n_49),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_96),
.Y(n_157)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_159),
.Y(n_188)
);

OAI22x1_ASAP7_75t_SL g155 ( 
.A1(n_147),
.A2(n_109),
.B1(n_102),
.B2(n_96),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_155),
.A2(n_133),
.B1(n_127),
.B2(n_116),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_158),
.Y(n_200)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_161),
.A2(n_166),
.B1(n_139),
.B2(n_15),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_98),
.B1(n_109),
.B2(n_102),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_179),
.B1(n_182),
.B2(n_139),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_140),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_167),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_141),
.B(n_136),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_147),
.A2(n_110),
.B1(n_28),
.B2(n_90),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_119),
.B(n_110),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_28),
.B(n_90),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_175),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_114),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_180),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_123),
.A2(n_114),
.B1(n_115),
.B2(n_125),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_150),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_5),
.C(n_7),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_118),
.C(n_113),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_182)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_12),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_184),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_186),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_195),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_196),
.C(n_203),
.Y(n_224)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_149),
.Y(n_190)
);

BUFx4f_ASAP7_75t_SL g225 ( 
.A(n_190),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_156),
.B(n_135),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_152),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_210),
.B1(n_169),
.B2(n_177),
.Y(n_231)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_120),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_183),
.B(n_214),
.Y(n_223)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_204),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_120),
.B(n_132),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_188),
.C(n_191),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_133),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_208),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_151),
.B(n_116),
.C(n_144),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_155),
.B(n_117),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_173),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_171),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_15),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_182),
.B1(n_154),
.B2(n_181),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_166),
.B(n_158),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_211),
.A2(n_200),
.B(n_196),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_160),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_153),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_154),
.B(n_162),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_211),
.C(n_208),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_175),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_217),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_221),
.A2(n_233),
.B1(n_236),
.B2(n_199),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

AOI221xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_235),
.B1(n_241),
.B2(n_194),
.C(n_197),
.Y(n_247)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_228),
.B(n_216),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_234),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_232),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_185),
.B1(n_172),
.B2(n_174),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_190),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_198),
.A2(n_178),
.B1(n_164),
.B2(n_186),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_192),
.B(n_168),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_168),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_242),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_209),
.C(n_187),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_224),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_203),
.B(n_193),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_195),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_230),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_229),
.A2(n_199),
.B1(n_206),
.B2(n_225),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_245),
.A2(n_258),
.B1(n_235),
.B2(n_229),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_247),
.A2(n_254),
.B(n_246),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_219),
.B(n_205),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_248),
.B(n_264),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_253),
.C(n_261),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_256),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_244),
.C(n_239),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_226),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_228),
.A2(n_217),
.B1(n_218),
.B2(n_205),
.Y(n_256)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_206),
.B1(n_218),
.B2(n_234),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_225),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_221),
.Y(n_276)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_226),
.C(n_227),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_235),
.C(n_249),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_259),
.B(n_220),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_273),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_236),
.Y(n_270)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_280),
.C(n_253),
.Y(n_291)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_260),
.B(n_220),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_231),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_281),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_276),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_277),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_254),
.B1(n_251),
.B2(n_245),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_265),
.Y(n_285)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_267),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_292),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_246),
.B(n_252),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_291),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_290),
.B(n_282),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_278),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_273),
.Y(n_295)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

AOI21x1_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_281),
.B(n_258),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_289),
.B(n_283),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_268),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_280),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_284),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_304),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_284),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_310),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_271),
.Y(n_310)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_312),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_291),
.C(n_272),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_313),
.A2(n_296),
.B(n_272),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_303),
.B1(n_298),
.B2(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

AOI211xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_255),
.B(n_295),
.C(n_306),
.Y(n_317)
);

OAI21x1_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_311),
.B(n_310),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_315),
.B(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_323),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_321),
.B(n_311),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_324),
.Y(n_326)
);


endmodule