module real_jpeg_9962_n_17 (n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_1),
.A2(n_57),
.B1(n_65),
.B2(n_68),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_2),
.A2(n_11),
.B(n_32),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_3),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_3),
.A2(n_65),
.B1(n_68),
.B2(n_92),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_92),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_92),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_4),
.A2(n_65),
.B1(n_68),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_4),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_157),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_157),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_4),
.A2(n_23),
.B1(n_25),
.B2(n_157),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_5),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_10),
.A2(n_65),
.B1(n_68),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_10),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_109),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_109),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_10),
.A2(n_23),
.B1(n_25),
.B2(n_109),
.Y(n_245)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_11),
.A2(n_48),
.B(n_60),
.C(n_89),
.D(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_11),
.B(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_11),
.B(n_46),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_11),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_11),
.A2(n_110),
.B(n_113),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_11),
.A2(n_31),
.B(n_42),
.C(n_145),
.D(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_11),
.B(n_31),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_11),
.B(n_35),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_126),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_13),
.A2(n_23),
.B1(n_25),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_55),
.B1(n_65),
.B2(n_68),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_14),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_14),
.A2(n_22),
.B1(n_65),
.B2(n_68),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_14),
.A2(n_22),
.B1(n_47),
.B2(n_48),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_15),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_15),
.A2(n_34),
.B1(n_65),
.B2(n_68),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_16),
.A2(n_47),
.B1(n_48),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_16),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_16),
.A2(n_65),
.B1(n_68),
.B2(n_104),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_104),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_16),
.A2(n_23),
.B1(n_25),
.B2(n_104),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_78),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_76),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_20),
.B(n_36),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_21),
.A2(n_26),
.B1(n_35),
.B2(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_23),
.A2(n_28),
.B(n_126),
.C(n_188),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_26),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_26),
.B(n_208),
.Y(n_217)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_27),
.A2(n_30),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_27),
.A2(n_30),
.B1(n_216),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_27),
.A2(n_207),
.B(n_245),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_27),
.A2(n_30),
.B1(n_54),
.B2(n_289),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_30),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_30),
.A2(n_217),
.B(n_289),
.Y(n_288)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_35),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_71),
.C(n_73),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_37),
.A2(n_38),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_52),
.C(n_58),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_39),
.A2(n_40),
.B1(n_58),
.B2(n_314),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_41),
.A2(n_50),
.B1(n_166),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_41),
.A2(n_202),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_46),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_42),
.B(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_42),
.A2(n_46),
.B1(n_242),
.B2(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_42),
.A2(n_46),
.B1(n_261),
.B2(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_43),
.B(n_48),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_45),
.A2(n_47),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_61),
.B(n_63),
.C(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_50),
.B(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_50),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_50),
.A2(n_167),
.B(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_52),
.A2(n_53),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_58),
.A2(n_312),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_58),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_69),
.B(n_70),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_59),
.A2(n_69),
.B1(n_103),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_59),
.A2(n_143),
.B(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_59),
.A2(n_69),
.B1(n_199),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_59),
.A2(n_69),
.B1(n_227),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_59),
.A2(n_69),
.B1(n_236),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_60),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_60),
.A2(n_64),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_68),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_61),
.B(n_68),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_65),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_68),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_68),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_69),
.B(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_69),
.A2(n_105),
.B(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_70),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_71),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_332),
.B(n_338),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_305),
.A3(n_325),
.B1(n_330),
.B2(n_331),
.C(n_340),
.Y(n_79)
);

AOI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_253),
.A3(n_293),
.B1(n_299),
.B2(n_304),
.C(n_341),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_210),
.C(n_249),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_181),
.B(n_209),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_160),
.B(n_180),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_137),
.B(n_159),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_115),
.B(n_136),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_87),
.B(n_97),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_93),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_88),
.A2(n_93),
.B1(n_94),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_90),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_102),
.C(n_107),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_110),
.B(n_113),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_110),
.A2(n_128),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_110),
.A2(n_128),
.B1(n_192),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_110),
.A2(n_128),
.B1(n_225),
.B2(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_110),
.A2(n_128),
.B(n_234),
.Y(n_266)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_111),
.A2(n_112),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_114),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_111),
.A2(n_112),
.B1(n_156),
.B2(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_112),
.B(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_112),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_123),
.B(n_135),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_121),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_130),
.B(n_134),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_127),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_128),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_129),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_138),
.B(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_150),
.B2(n_158),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_142),
.Y(n_149)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_149),
.C(n_158),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_145),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_146),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_150),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_154),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_161),
.B(n_162),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_174),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_176),
.C(n_178),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_169),
.B2(n_173),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_170),
.C(n_171),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_175),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_176),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_182),
.B(n_183),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_196),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_185),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_185),
.B(n_195),
.C(n_196),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_190),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_204),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_198),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_203),
.C(n_204),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_211),
.A2(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_229),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_212),
.B(n_229),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_223),
.C(n_228),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_218),
.B1(n_219),
.B2(n_221),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_215),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_228),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_226),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_247),
.B2(n_248),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_237),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_232),
.B(n_237),
.C(n_248),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_235),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_243),
.C(n_246),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_243),
.B1(n_244),
.B2(n_246),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_240),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_247),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_250),
.B(n_251),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_271),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_254),
.B(n_271),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_264),
.C(n_270),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_255),
.A2(n_256),
.B1(n_264),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_260),
.C(n_262),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_264),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_265),
.A2(n_266),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_265),
.A2(n_284),
.B(n_288),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_267),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_267),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_268),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_291),
.B2(n_292),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_282),
.B2(n_283),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_283),
.C(n_292),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_279),
.B(n_281),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_279),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_280),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_281),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_281),
.A2(n_307),
.B1(n_316),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_290),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_286),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_294),
.A2(n_300),
.B(n_303),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_295),
.B(n_296),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_318),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_318),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_316),
.C(n_317),
.Y(n_306)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_308),
.A2(n_309),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_314),
.C(n_315),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_320),
.C(n_324),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_312),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_324),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_337),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_337),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_334),
.Y(n_336)
);


endmodule