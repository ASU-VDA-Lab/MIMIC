module fake_jpeg_15708_n_136 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_63),
.Y(n_71)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_51),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_2),
.B(n_3),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_46),
.B1(n_49),
.B2(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_48),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_44),
.B1(n_49),
.B2(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_0),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_42),
.B1(n_55),
.B2(n_43),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_56),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_0),
.Y(n_70)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_55),
.B1(n_50),
.B2(n_45),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_76),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_21),
.B1(n_39),
.B2(n_38),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_2),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_84),
.B1(n_90),
.B2(n_96),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_1),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_1),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_91),
.Y(n_107)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_5),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_94),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_6),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_6),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_7),
.B(n_8),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_9),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_106),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_11),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_80),
.B(n_104),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_116),
.B(n_117),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

OAI211xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_98),
.B(n_99),
.C(n_97),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_120),
.A2(n_110),
.B1(n_92),
.B2(n_101),
.Y(n_122)
);

CKINVDCx6p67_ASAP7_75t_R g121 ( 
.A(n_120),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_122),
.A2(n_115),
.B1(n_118),
.B2(n_17),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_125),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_126),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_20),
.B(n_23),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_24),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_25),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_27),
.B(n_29),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_133),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_134),
.A2(n_35),
.B(n_36),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_37),
.Y(n_136)
);


endmodule