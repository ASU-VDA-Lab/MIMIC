module fake_jpeg_30468_n_528 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_528);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_528;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_53),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_21),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_54),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_106),
.Y(n_119)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_9),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_83),
.Y(n_120)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_30),
.A2(n_9),
.B(n_16),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_25),
.C(n_34),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_74),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_34),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_85),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_18),
.B(n_8),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_104),
.Y(n_136)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_101),
.Y(n_138)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_105),
.Y(n_158)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_108),
.Y(n_123)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_22),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_112),
.B(n_148),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_59),
.A2(n_48),
.B1(n_52),
.B2(n_24),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_116),
.A2(n_126),
.B1(n_153),
.B2(n_11),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_57),
.A2(n_52),
.B1(n_49),
.B2(n_51),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_121),
.A2(n_173),
.B1(n_109),
.B2(n_104),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_83),
.A2(n_23),
.B1(n_40),
.B2(n_38),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_108),
.A2(n_52),
.B1(n_50),
.B2(n_47),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_137),
.A2(n_82),
.B1(n_53),
.B2(n_42),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_93),
.B(n_23),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_142),
.B(n_150),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_54),
.B(n_20),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_60),
.A2(n_40),
.B1(n_20),
.B2(n_27),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_76),
.B(n_27),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_172),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_88),
.B(n_29),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_157),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_80),
.B(n_38),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_62),
.B(n_29),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_68),
.A2(n_52),
.B1(n_51),
.B2(n_50),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_176),
.B(n_189),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g242 ( 
.A(n_177),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_119),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_178),
.B(n_181),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_84),
.B1(n_75),
.B2(n_72),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_179),
.A2(n_207),
.B1(n_220),
.B2(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_180),
.Y(n_259)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_182),
.Y(n_257)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_183),
.B(n_185),
.Y(n_268)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_186),
.Y(n_261)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_116),
.A2(n_45),
.B1(n_24),
.B2(n_44),
.Y(n_189)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_120),
.B(n_22),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_194),
.B(n_199),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_113),
.A2(n_86),
.B1(n_101),
.B2(n_96),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_196),
.A2(n_197),
.B1(n_213),
.B2(n_215),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_113),
.A2(n_33),
.B1(n_47),
.B2(n_45),
.Y(n_197)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_198),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_22),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_202),
.Y(n_269)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_203),
.Y(n_273)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_204),
.Y(n_256)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_205),
.Y(n_279)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_122),
.B(n_85),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_206),
.B(n_217),
.C(n_225),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_173),
.A2(n_70),
.B1(n_69),
.B2(n_73),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_128),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_133),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_209),
.B(n_221),
.Y(n_243)
);

INVx3_ASAP7_75t_SL g211 ( 
.A(n_170),
.Y(n_211)
);

INVx6_ASAP7_75t_SL g251 ( 
.A(n_211),
.Y(n_251)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_222),
.Y(n_249)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_123),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_135),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_22),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_163),
.A2(n_33),
.B1(n_42),
.B2(n_44),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_218),
.A2(n_219),
.B1(n_224),
.B2(n_230),
.Y(n_265)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_115),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_137),
.A2(n_37),
.B1(n_73),
.B2(n_71),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_115),
.A2(n_94),
.B1(n_71),
.B2(n_69),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_37),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_110),
.A2(n_37),
.B1(n_94),
.B2(n_9),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_226),
.A2(n_231),
.B1(n_145),
.B2(n_164),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_160),
.B(n_37),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_227),
.A2(n_229),
.B(n_161),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_110),
.A2(n_8),
.B1(n_15),
.B2(n_12),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_228),
.A2(n_158),
.B1(n_164),
.B2(n_131),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_111),
.B(n_0),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_146),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_130),
.A2(n_7),
.B1(n_15),
.B2(n_11),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_121),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_232),
.B(n_125),
.Y(n_241)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_128),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_233),
.A2(n_161),
.B1(n_132),
.B2(n_169),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_236),
.A2(n_241),
.B1(n_275),
.B2(n_276),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_200),
.B(n_168),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_255),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_L g245 ( 
.A(n_191),
.B(n_144),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_191),
.B(n_194),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_266),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_254),
.A2(n_274),
.B1(n_202),
.B2(n_175),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g262 ( 
.A(n_190),
.B(n_194),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_201),
.C(n_162),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_217),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_190),
.B(n_125),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_232),
.A2(n_146),
.B1(n_169),
.B2(n_131),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_222),
.A2(n_151),
.B1(n_145),
.B2(n_139),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_189),
.A2(n_151),
.B1(n_139),
.B2(n_152),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_190),
.B(n_152),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_278),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_132),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_249),
.A2(n_176),
.B1(n_216),
.B2(n_206),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_282),
.A2(n_286),
.B1(n_292),
.B2(n_313),
.Y(n_343)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_242),
.Y(n_287)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_287),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_250),
.B(n_210),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_293),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_249),
.A2(n_206),
.B1(n_207),
.B2(n_229),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_203),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_294),
.B(n_302),
.Y(n_340)
);

OAI32xp33_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_193),
.A3(n_192),
.B1(n_186),
.B2(n_182),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_300),
.Y(n_324)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_243),
.B(n_205),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_298),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_262),
.B(n_199),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_242),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_299),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_262),
.B(n_199),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_303),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_252),
.A2(n_217),
.B1(n_225),
.B2(n_227),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_262),
.B(n_225),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_252),
.A2(n_227),
.B1(n_204),
.B2(n_188),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_305),
.A2(n_273),
.B1(n_258),
.B2(n_247),
.Y(n_329)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_239),
.Y(n_306)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_306),
.Y(n_345)
);

OAI32xp33_ASAP7_75t_L g307 ( 
.A1(n_278),
.A2(n_219),
.A3(n_215),
.B1(n_213),
.B2(n_230),
.Y(n_307)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_255),
.B(n_198),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_309),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_249),
.B(n_212),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_310),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_235),
.B(n_211),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_311),
.B(n_235),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_244),
.B(n_177),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_312),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_246),
.A2(n_184),
.B1(n_187),
.B2(n_143),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_316),
.Y(n_321)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_237),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_271),
.B(n_177),
.C(n_214),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_280),
.A2(n_290),
.B1(n_252),
.B2(n_246),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_318),
.A2(n_329),
.B1(n_335),
.B2(n_341),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_271),
.C(n_264),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_338),
.C(n_314),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_322),
.B(n_297),
.Y(n_370)
);

OA22x2_ASAP7_75t_L g323 ( 
.A1(n_290),
.A2(n_241),
.B1(n_276),
.B2(n_275),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_327),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_291),
.A2(n_271),
.B1(n_248),
.B2(n_265),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_309),
.A2(n_264),
.B(n_273),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_328),
.A2(n_346),
.B(n_238),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_284),
.A2(n_236),
.B1(n_259),
.B2(n_267),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_281),
.B(n_268),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_296),
.A2(n_251),
.B1(n_259),
.B2(n_253),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_282),
.A2(n_251),
.B1(n_267),
.B2(n_240),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_344),
.A2(n_305),
.B1(n_308),
.B2(n_293),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_284),
.A2(n_268),
.B(n_260),
.Y(n_346)
);

OAI32xp33_ASAP7_75t_L g347 ( 
.A1(n_288),
.A2(n_258),
.A3(n_247),
.B1(n_256),
.B2(n_279),
.Y(n_347)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_347),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_349),
.A2(n_371),
.B1(n_373),
.B2(n_375),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_333),
.B(n_289),
.Y(n_350)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_350),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_348),
.A2(n_313),
.B1(n_294),
.B2(n_292),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_351),
.B(n_372),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_328),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_353),
.B(n_363),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_346),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_354),
.Y(n_400)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_339),
.Y(n_355)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_355),
.Y(n_387)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_320),
.Y(n_357)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_320),
.Y(n_358)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_333),
.B(n_288),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_366),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_342),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_360),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

BUFx8_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_322),
.B(n_311),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_319),
.Y(n_386)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_325),
.Y(n_365)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_365),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_329),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_301),
.C(n_298),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_374),
.C(n_340),
.Y(n_390)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_347),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_370),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_343),
.A2(n_302),
.B1(n_303),
.B2(n_295),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_348),
.A2(n_294),
.B1(n_286),
.B2(n_316),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_343),
.A2(n_307),
.B1(n_316),
.B2(n_283),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_321),
.B(n_285),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_324),
.A2(n_315),
.B1(n_310),
.B2(n_306),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_376),
.B(n_336),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_377),
.A2(n_340),
.B(n_326),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_256),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_337),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_362),
.A2(n_372),
.B(n_369),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_379),
.A2(n_383),
.B(n_270),
.Y(n_426)
);

AO21x2_ASAP7_75t_SL g381 ( 
.A1(n_352),
.A2(n_318),
.B(n_323),
.Y(n_381)
);

AO21x2_ASAP7_75t_L g422 ( 
.A1(n_381),
.A2(n_384),
.B(n_382),
.Y(n_422)
);

OAI22x1_ASAP7_75t_SL g382 ( 
.A1(n_362),
.A2(n_323),
.B1(n_324),
.B2(n_327),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_382),
.A2(n_399),
.B1(n_371),
.B2(n_367),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_362),
.A2(n_332),
.B(n_334),
.Y(n_383)
);

AO22x1_ASAP7_75t_L g384 ( 
.A1(n_352),
.A2(n_323),
.B1(n_344),
.B2(n_335),
.Y(n_384)
);

AO22x1_ASAP7_75t_L g418 ( 
.A1(n_384),
.A2(n_365),
.B1(n_361),
.B2(n_355),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_386),
.B(n_389),
.C(n_390),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_388),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_374),
.B(n_338),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_361),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_375),
.A2(n_323),
.B1(n_340),
.B2(n_317),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_356),
.A2(n_317),
.B1(n_332),
.B2(n_334),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_401),
.A2(n_349),
.B1(n_360),
.B2(n_359),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_373),
.A2(n_331),
.B(n_345),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_403),
.A2(n_261),
.B(n_257),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_364),
.B(n_345),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_239),
.C(n_299),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_405),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_354),
.A2(n_330),
.B1(n_339),
.B2(n_234),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_406),
.A2(n_287),
.B1(n_253),
.B2(n_234),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_409),
.A2(n_418),
.B1(n_421),
.B2(n_422),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_408),
.B(n_378),
.Y(n_410)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

OAI32xp33_ASAP7_75t_L g411 ( 
.A1(n_393),
.A2(n_370),
.A3(n_351),
.B1(n_350),
.B2(n_356),
.Y(n_411)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_411),
.Y(n_445)
);

AOI21xp33_ASAP7_75t_L g412 ( 
.A1(n_397),
.A2(n_377),
.B(n_357),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_412),
.A2(n_403),
.B(n_402),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_413),
.A2(n_402),
.B1(n_384),
.B2(n_401),
.Y(n_443)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_414),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_330),
.Y(n_415)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_415),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_368),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_417),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_392),
.B(n_358),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_393),
.B(n_279),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_419),
.B(n_425),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_432),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_380),
.B(n_304),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_426),
.B(n_428),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_270),
.C(n_261),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_431),
.C(n_390),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_394),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_429),
.B(n_430),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_391),
.B(n_267),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_233),
.C(n_208),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_391),
.B(n_407),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_380),
.B(n_240),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_433),
.B(n_399),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_418),
.Y(n_437)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_437),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_438),
.B(n_455),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_411),
.Y(n_471)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_442),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_443),
.A2(n_453),
.B1(n_426),
.B2(n_419),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_418),
.A2(n_385),
.B1(n_379),
.B2(n_381),
.Y(n_446)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_446),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_423),
.B(n_389),
.C(n_402),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_448),
.B(n_452),
.C(n_454),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_385),
.C(n_388),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_414),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_420),
.B(n_383),
.C(n_387),
.Y(n_454)
);

MAJx2_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_424),
.C(n_410),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_413),
.B(n_381),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_456),
.B(n_428),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_458),
.B(n_465),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_462),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_445),
.A2(n_434),
.B(n_453),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_443),
.A2(n_409),
.B1(n_422),
.B2(n_424),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_464),
.A2(n_472),
.B1(n_446),
.B2(n_422),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_435),
.B(n_415),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_431),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_469),
.C(n_444),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_449),
.A2(n_422),
.B(n_416),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_467),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_433),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_441),
.B(n_425),
.C(n_417),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_470),
.B(n_471),
.C(n_473),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_440),
.A2(n_422),
.B1(n_452),
.B2(n_456),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_439),
.B(n_387),
.C(n_432),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_SL g474 ( 
.A1(n_468),
.A2(n_450),
.B1(n_422),
.B2(n_429),
.Y(n_474)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_474),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_472),
.A2(n_468),
.B1(n_459),
.B2(n_440),
.Y(n_477)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_477),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_460),
.A2(n_451),
.B(n_455),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_479),
.A2(n_480),
.B(n_482),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_460),
.A2(n_447),
.B(n_436),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_481),
.B(n_484),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_439),
.C(n_442),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_458),
.A2(n_464),
.B1(n_457),
.B2(n_463),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_483),
.B(n_463),
.C(n_461),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_394),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_486),
.B(n_487),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_444),
.C(n_430),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_473),
.B(n_407),
.C(n_396),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_488),
.B(n_469),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_478),
.C(n_482),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_492),
.B(n_493),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_394),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_462),
.C(n_467),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_495),
.B(n_499),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_474),
.A2(n_381),
.B(n_395),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_496),
.A2(n_234),
.B(n_195),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_396),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_395),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_500),
.B(n_487),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_494),
.A2(n_489),
.B(n_493),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_501),
.A2(n_509),
.B(n_510),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_504),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_475),
.C(n_240),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_505),
.B(n_508),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_17),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_490),
.A2(n_7),
.B1(n_15),
.B2(n_10),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_5),
.C(n_10),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_498),
.B(n_496),
.C(n_7),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_513),
.B(n_515),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_507),
.B(n_5),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_507),
.A2(n_7),
.B(n_10),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_516),
.A2(n_4),
.B(n_9),
.Y(n_519)
);

MAJx2_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_502),
.C(n_4),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_518),
.B(n_511),
.Y(n_521)
);

OAI321xp33_ASAP7_75t_L g522 ( 
.A1(n_519),
.A2(n_520),
.A3(n_17),
.B1(n_4),
.B2(n_2),
.C(n_1),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_514),
.B(n_4),
.Y(n_520)
);

AO21x1_ASAP7_75t_L g523 ( 
.A1(n_521),
.A2(n_522),
.B(n_517),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_0),
.B(n_1),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_0),
.C(n_1),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_0),
.C(n_1),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_2),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_2),
.B(n_507),
.Y(n_528)
);


endmodule