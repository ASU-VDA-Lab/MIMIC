module fake_jpeg_3914_n_312 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx2_ASAP7_75t_SL g95 ( 
.A(n_36),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_22),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_38),
.B(n_46),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_39),
.B(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_13),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_0),
.Y(n_46)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_47),
.B(n_25),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_33),
.B1(n_16),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_50),
.A2(n_54),
.B1(n_64),
.B2(n_69),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_29),
.B1(n_22),
.B2(n_34),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_51),
.A2(n_34),
.A3(n_21),
.B1(n_19),
.B2(n_24),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_33),
.B1(n_16),
.B2(n_26),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_89),
.B1(n_96),
.B2(n_49),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_16),
.B1(n_31),
.B2(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_17),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_59),
.B(n_62),
.Y(n_118)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_63),
.B(n_68),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_32),
.C(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_28),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_23),
.B1(n_20),
.B2(n_30),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_37),
.A2(n_23),
.B1(n_20),
.B2(n_30),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_70),
.A2(n_74),
.B1(n_93),
.B2(n_0),
.Y(n_119)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_75),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_32),
.Y(n_73)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_37),
.A2(n_21),
.B1(n_18),
.B2(n_19),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_11),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_11),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_87),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_11),
.B(n_12),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_97),
.B(n_99),
.C(n_51),
.Y(n_115)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_85),
.Y(n_100)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_86),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_10),
.Y(n_87)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_90),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_35),
.A2(n_21),
.B1(n_18),
.B2(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_39),
.B(n_22),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_39),
.B(n_24),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_94),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_34),
.B1(n_21),
.B2(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_9),
.Y(n_94)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_44),
.A2(n_19),
.B(n_25),
.C(n_9),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_102),
.A2(n_107),
.B1(n_81),
.B2(n_84),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_93),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_19),
.B(n_24),
.C(n_3),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_117),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_10),
.B(n_2),
.C(n_5),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_80),
.B(n_92),
.C(n_5),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_129),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_127),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_95),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_131),
.B(n_139),
.Y(n_170)
);

NAND2x1_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_98),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_132),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_64),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_140),
.Y(n_176)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_138),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_113),
.B1(n_102),
.B2(n_50),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_136),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_99),
.B1(n_54),
.B2(n_74),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_142),
.B1(n_108),
.B2(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_70),
.B(n_82),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_66),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_59),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_141),
.B(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_63),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_96),
.B1(n_49),
.B2(n_60),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_145),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_60),
.B1(n_81),
.B2(n_77),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_78),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_149),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_53),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_157),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_76),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_162),
.B(n_163),
.Y(n_187)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_155),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_123),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_156),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_106),
.B(n_65),
.Y(n_154)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_109),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_72),
.B(n_71),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_0),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_0),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_161),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_111),
.A2(n_85),
.B1(n_72),
.B2(n_6),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_2),
.B(n_5),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_103),
.A2(n_114),
.B(n_110),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_185),
.B1(n_186),
.B2(n_151),
.Y(n_214)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_180),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_110),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_191),
.B(n_162),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_174),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_129),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_148),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_131),
.B(n_100),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_139),
.Y(n_207)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_188),
.Y(n_219)
);

AO22x1_ASAP7_75t_SL g185 ( 
.A1(n_131),
.A2(n_125),
.B1(n_114),
.B2(n_112),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_112),
.B1(n_126),
.B2(n_120),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_133),
.B(n_120),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_151),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_126),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_197),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_137),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_193),
.B(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_100),
.Y(n_197)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_199),
.B(n_161),
.Y(n_223)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_204),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_136),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_221),
.C(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_207),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_192),
.B(n_138),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_128),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_185),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_177),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_216),
.B1(n_225),
.B2(n_179),
.Y(n_229)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_170),
.A2(n_156),
.B(n_135),
.C(n_132),
.D(n_151),
.Y(n_215)
);

OAI22x1_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_147),
.B1(n_160),
.B2(n_144),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_222),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_190),
.B(n_135),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_182),
.A2(n_130),
.B(n_149),
.Y(n_222)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_170),
.A2(n_146),
.B(n_141),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_229),
.B(n_175),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_187),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_239),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_176),
.C(n_171),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_243),
.C(n_206),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_214),
.A2(n_172),
.B1(n_175),
.B2(n_184),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_172),
.B1(n_173),
.B2(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_174),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_245),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_195),
.C(n_193),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

OAI321xp33_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_221),
.A3(n_213),
.B1(n_222),
.B2(n_215),
.C(n_209),
.Y(n_246)
);

OAI321xp33_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_173),
.A3(n_195),
.B1(n_220),
.B2(n_202),
.C(n_207),
.Y(n_249)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_201),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_250),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_218),
.B(n_217),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_235),
.A2(n_218),
.B(n_217),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_253),
.A2(n_245),
.B1(n_234),
.B2(n_165),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_226),
.Y(n_255)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

XOR2x2_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_187),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_227),
.C(n_230),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_262),
.Y(n_271)
);

BUFx12f_ASAP7_75t_SL g259 ( 
.A(n_248),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_260),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_228),
.A2(n_191),
.B1(n_169),
.B2(n_203),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_186),
.B1(n_142),
.B2(n_210),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_181),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_243),
.C(n_238),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_264),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_266),
.B(n_232),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_255),
.C(n_262),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_265),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_237),
.C(n_227),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_276),
.C(n_277),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_261),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_236),
.C(n_196),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_236),
.C(n_164),
.Y(n_277)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_272),
.A2(n_256),
.B1(n_247),
.B2(n_205),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_285),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_274),
.A2(n_250),
.B(n_251),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_280),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_283),
.C(n_286),
.Y(n_296)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_253),
.C(n_263),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_233),
.C(n_244),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_165),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_273),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_292),
.Y(n_301)
);

OAI221xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_273),
.B1(n_277),
.B2(n_266),
.C(n_269),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_142),
.B1(n_268),
.B2(n_231),
.Y(n_294)
);

NAND4xp25_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_130),
.C(n_178),
.D(n_160),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_285),
.A2(n_231),
.B1(n_281),
.B2(n_204),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_180),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_298),
.A2(n_167),
.B(n_158),
.Y(n_303)
);

XNOR2x1_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_281),
.Y(n_299)
);

AOI221xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_302),
.B1(n_304),
.B2(n_291),
.C(n_293),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_294),
.B1(n_167),
.B2(n_290),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_296),
.C(n_199),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_208),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.C(n_307),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_296),
.B1(n_282),
.B2(n_252),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_308),
.B(n_301),
.C(n_168),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_308),
.B1(n_100),
.B2(n_134),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_309),
.Y(n_312)
);


endmodule