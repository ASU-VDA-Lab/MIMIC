module real_aes_15489_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g852 ( .A(n_0), .B(n_853), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_1), .A2(n_4), .B1(n_265), .B2(n_266), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_2), .A2(n_42), .B1(n_122), .B2(n_192), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_3), .A2(n_23), .B1(n_192), .B2(n_201), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_5), .A2(n_15), .B1(n_499), .B2(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_6), .A2(n_61), .B1(n_150), .B2(n_151), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_7), .A2(n_16), .B1(n_122), .B2(n_124), .Y(n_121) );
INVx1_ASAP7_75t_L g853 ( .A(n_8), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_9), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_10), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_11), .A2(n_17), .B1(n_500), .B2(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g802 ( .A(n_12), .B(n_38), .Y(n_802) );
BUFx2_ASAP7_75t_L g848 ( .A(n_12), .Y(n_848) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_13), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_14), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_18), .A2(n_102), .B1(n_266), .B2(n_499), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_19), .A2(n_37), .B1(n_158), .B2(n_516), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_20), .B(n_157), .Y(n_513) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_21), .A2(n_58), .B(n_135), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_22), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_24), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_25), .B(n_127), .Y(n_221) );
INVx4_ASAP7_75t_R g174 ( .A(n_26), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_27), .A2(n_54), .B1(n_819), .B2(n_820), .Y(n_818) );
CKINVDCx5p33_ASAP7_75t_R g819 ( .A(n_27), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_28), .A2(n_46), .B1(n_129), .B2(n_263), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_29), .A2(n_53), .B1(n_129), .B2(n_499), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_30), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_31), .B(n_516), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_32), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_33), .B(n_192), .Y(n_227) );
INVx1_ASAP7_75t_L g270 ( .A(n_34), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_SL g198 ( .A1(n_35), .A2(n_122), .B(n_126), .C(n_199), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_36), .A2(n_55), .B1(n_122), .B2(n_129), .Y(n_210) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_38), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_39), .A2(n_87), .B1(n_122), .B2(n_489), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_40), .A2(n_80), .B1(n_787), .B2(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_40), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_41), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_43), .A2(n_45), .B1(n_122), .B2(n_124), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_44), .A2(n_59), .B1(n_499), .B2(n_551), .Y(n_567) );
INVx1_ASAP7_75t_L g224 ( .A(n_47), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_48), .B(n_122), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g831 ( .A1(n_49), .A2(n_832), .B(n_839), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_50), .Y(n_243) );
INVx2_ASAP7_75t_L g797 ( .A(n_51), .Y(n_797) );
BUFx3_ASAP7_75t_L g800 ( .A(n_52), .Y(n_800) );
INVx1_ASAP7_75t_L g815 ( .A(n_52), .Y(n_815) );
INVx1_ASAP7_75t_L g820 ( .A(n_54), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_56), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_57), .A2(n_88), .B1(n_122), .B2(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g784 ( .A1(n_60), .A2(n_785), .B1(n_786), .B2(n_789), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_60), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_62), .A2(n_75), .B1(n_263), .B2(n_551), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_63), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_64), .A2(n_78), .B1(n_122), .B2(n_124), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_65), .A2(n_100), .B1(n_499), .B2(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g135 ( .A(n_66), .Y(n_135) );
AND2x4_ASAP7_75t_L g137 ( .A(n_67), .B(n_138), .Y(n_137) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_68), .A2(n_105), .B1(n_842), .B2(n_854), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_69), .A2(n_90), .B1(n_129), .B2(n_263), .Y(n_262) );
AO22x1_ASAP7_75t_L g155 ( .A1(n_70), .A2(n_76), .B1(n_156), .B2(n_158), .Y(n_155) );
INVx1_ASAP7_75t_L g138 ( .A(n_71), .Y(n_138) );
AND2x2_ASAP7_75t_L g202 ( .A(n_72), .B(n_203), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_73), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_74), .B(n_150), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_77), .B(n_192), .Y(n_244) );
INVx2_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
INVx1_ASAP7_75t_L g788 ( .A(n_80), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_81), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_82), .B(n_203), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_83), .A2(n_99), .B1(n_129), .B2(n_150), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_84), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_85), .B(n_133), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_86), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_89), .B(n_203), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_91), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_92), .B(n_203), .Y(n_240) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_92), .Y(n_823) );
INVx1_ASAP7_75t_L g477 ( .A(n_93), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_93), .B(n_829), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_94), .A2(n_783), .B1(n_790), .B2(n_791), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_94), .Y(n_790) );
NAND2xp33_ASAP7_75t_L g517 ( .A(n_95), .B(n_157), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_96), .A2(n_131), .B(n_150), .C(n_170), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g840 ( .A(n_97), .Y(n_840) );
AND2x2_ASAP7_75t_L g179 ( .A(n_98), .B(n_180), .Y(n_179) );
AOI22xp33_ASAP7_75t_SL g822 ( .A1(n_101), .A2(n_823), .B1(n_824), .B2(n_825), .Y(n_822) );
INVxp67_ASAP7_75t_SL g824 ( .A(n_101), .Y(n_824) );
NAND2xp33_ASAP7_75t_L g248 ( .A(n_103), .B(n_175), .Y(n_248) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_803), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_793), .Y(n_106) );
AOI22xp33_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_781), .B1(n_782), .B2(n_792), .Y(n_107) );
INVx2_ASAP7_75t_L g792 ( .A(n_108), .Y(n_792) );
AO22x2_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_473), .B1(n_474), .B2(n_478), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
NOR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_387), .Y(n_110) );
NAND4xp75_ASAP7_75t_L g111 ( .A(n_112), .B(n_292), .C(n_334), .D(n_358), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OAI211xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_181), .B(n_229), .C(n_271), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g378 ( .A(n_116), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g472 ( .A(n_116), .B(n_409), .Y(n_472) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_142), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g287 ( .A(n_118), .B(n_239), .Y(n_287) );
AND2x2_ASAP7_75t_L g328 ( .A(n_118), .B(n_289), .Y(n_328) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g235 ( .A(n_119), .B(n_164), .Y(n_235) );
OR2x2_ASAP7_75t_L g253 ( .A(n_119), .B(n_164), .Y(n_253) );
INVx2_ASAP7_75t_L g279 ( .A(n_119), .Y(n_279) );
AND2x2_ASAP7_75t_L g309 ( .A(n_119), .B(n_239), .Y(n_309) );
AND2x2_ASAP7_75t_L g338 ( .A(n_119), .B(n_163), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_119), .B(n_290), .Y(n_374) );
AO31x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_132), .A3(n_136), .B(n_139), .Y(n_119) );
OAI22x1_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_125), .B1(n_128), .B2(n_130), .Y(n_120) );
INVx4_ASAP7_75t_L g124 ( .A(n_122), .Y(n_124) );
INVx1_ASAP7_75t_L g500 ( .A(n_122), .Y(n_500) );
INVx1_ASAP7_75t_L g551 ( .A(n_122), .Y(n_551) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_123), .Y(n_129) );
INVx1_ASAP7_75t_L g150 ( .A(n_123), .Y(n_150) );
INVx1_ASAP7_75t_L g152 ( .A(n_123), .Y(n_152) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_123), .Y(n_157) );
INVx1_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_123), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_123), .Y(n_176) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_123), .Y(n_192) );
INVx1_ASAP7_75t_L g194 ( .A(n_123), .Y(n_194) );
INVx2_ASAP7_75t_L g201 ( .A(n_123), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_124), .A2(n_243), .B(n_244), .C(n_245), .Y(n_242) );
O2A1O1Ixp5_ASAP7_75t_L g511 ( .A1(n_124), .A2(n_126), .B(n_512), .C(n_513), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_125), .A2(n_146), .B1(n_209), .B2(n_210), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_125), .A2(n_130), .B1(n_262), .B2(n_264), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_125), .A2(n_130), .B1(n_488), .B2(n_490), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_125), .A2(n_498), .B1(n_501), .B2(n_502), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_125), .A2(n_515), .B(n_517), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_125), .A2(n_523), .B1(n_524), .B2(n_525), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_125), .A2(n_502), .B1(n_534), .B2(n_536), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_125), .A2(n_524), .B1(n_543), .B2(n_544), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_125), .A2(n_524), .B1(n_550), .B2(n_552), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_125), .A2(n_524), .B1(n_566), .B2(n_567), .Y(n_565) );
INVx6_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_126), .B(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_126), .A2(n_248), .B(n_249), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_126), .A2(n_145), .B(n_155), .C(n_161), .Y(n_291) );
BUFx8_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g131 ( .A(n_127), .Y(n_131) );
INVx2_ASAP7_75t_L g148 ( .A(n_127), .Y(n_148) );
INVx1_ASAP7_75t_L g197 ( .A(n_127), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_129), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g265 ( .A(n_129), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_130), .B(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_SL g502 ( .A(n_131), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_132), .B(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_132), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g141 ( .A(n_133), .Y(n_141) );
OAI21xp33_ASAP7_75t_L g161 ( .A1(n_133), .A2(n_153), .B(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_134), .Y(n_204) );
INVx2_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
AO31x2_ASAP7_75t_L g521 ( .A1(n_136), .A2(n_211), .A3(n_522), .B(n_526), .Y(n_521) );
AO31x2_ASAP7_75t_L g532 ( .A1(n_136), .A2(n_187), .A3(n_533), .B(n_537), .Y(n_532) );
AO31x2_ASAP7_75t_L g541 ( .A1(n_136), .A2(n_486), .A3(n_542), .B(n_546), .Y(n_541) );
BUFx10_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g162 ( .A(n_137), .Y(n_162) );
BUFx10_ASAP7_75t_L g212 ( .A(n_137), .Y(n_212) );
INVx1_ASAP7_75t_L g268 ( .A(n_137), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
INVx2_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
BUFx2_ASAP7_75t_L g187 ( .A(n_141), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_141), .B(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_141), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g351 ( .A(n_142), .B(n_280), .Y(n_351) );
INVx2_ASAP7_75t_L g446 ( .A(n_142), .Y(n_446) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_163), .Y(n_142) );
INVx2_ASAP7_75t_L g234 ( .A(n_143), .Y(n_234) );
AND2x4_ASAP7_75t_L g277 ( .A(n_143), .B(n_164), .Y(n_277) );
AOI21x1_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_154), .B(n_160), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_149), .B(n_153), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_146), .A2(n_226), .B(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g524 ( .A(n_147), .Y(n_524) );
BUFx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g246 ( .A(n_148), .Y(n_246) );
INVx1_ASAP7_75t_L g535 ( .A(n_151), .Y(n_535) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_152), .B(n_171), .Y(n_170) );
INVxp67_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g499 ( .A(n_157), .Y(n_499) );
OAI21xp33_ASAP7_75t_SL g220 ( .A1(n_158), .A2(n_221), .B(n_222), .Y(n_220) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_162), .A2(n_189), .B(n_198), .Y(n_188) );
AND2x2_ASAP7_75t_L g436 ( .A(n_163), .B(n_234), .Y(n_436) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g300 ( .A(n_164), .Y(n_300) );
AND2x2_ASAP7_75t_L g357 ( .A(n_164), .B(n_239), .Y(n_357) );
AND2x2_ASAP7_75t_L g372 ( .A(n_164), .B(n_280), .Y(n_372) );
AND2x2_ASAP7_75t_L g394 ( .A(n_164), .B(n_234), .Y(n_394) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B(n_179), .Y(n_164) );
AO31x2_ASAP7_75t_L g548 ( .A1(n_165), .A2(n_267), .A3(n_549), .B(n_553), .Y(n_548) );
AO31x2_ASAP7_75t_L g564 ( .A1(n_165), .A2(n_503), .A3(n_565), .B(n_568), .Y(n_564) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_167), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_SL g537 ( .A(n_167), .B(n_538), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_178), .Y(n_168) );
OAI22xp33_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B1(n_176), .B2(n_177), .Y(n_173) );
INVx2_ASAP7_75t_L g263 ( .A(n_175), .Y(n_263) );
INVx1_ASAP7_75t_L g516 ( .A(n_175), .Y(n_516) );
INVx1_ASAP7_75t_L g545 ( .A(n_176), .Y(n_545) );
INVx1_ASAP7_75t_L g503 ( .A(n_178), .Y(n_503) );
OAI211xp5_ASAP7_75t_SL g441 ( .A1(n_181), .A2(n_442), .B(n_444), .C(n_451), .Y(n_441) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_215), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_L g428 ( .A(n_184), .B(n_364), .Y(n_428) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_205), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_185), .B(n_217), .Y(n_327) );
INVxp67_ASAP7_75t_L g341 ( .A(n_185), .Y(n_341) );
AND2x2_ASAP7_75t_L g361 ( .A(n_185), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_185), .B(n_274), .Y(n_368) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g257 ( .A(n_186), .Y(n_257) );
AOI21x1_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_202), .Y(n_186) );
AO31x2_ASAP7_75t_L g260 ( .A1(n_187), .A2(n_261), .A3(n_267), .B(n_269), .Y(n_260) );
AO31x2_ASAP7_75t_L g496 ( .A1(n_187), .A2(n_497), .A3(n_503), .B(n_504), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_193), .B(n_196), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx2_ASAP7_75t_L g266 ( .A(n_194), .Y(n_266) );
BUFx4f_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_197), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx2_ASAP7_75t_SL g489 ( .A(n_201), .Y(n_489) );
INVx2_ASAP7_75t_L g211 ( .A(n_203), .Y(n_211) );
NOR2x1_ASAP7_75t_L g250 ( .A(n_203), .B(n_251), .Y(n_250) );
INVx4_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g228 ( .A(n_204), .B(n_212), .Y(n_228) );
BUFx3_ASAP7_75t_L g486 ( .A(n_204), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_204), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g509 ( .A(n_204), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_204), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_204), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g302 ( .A(n_205), .B(n_284), .Y(n_302) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g350 ( .A(n_206), .B(n_257), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_206), .B(n_260), .Y(n_356) );
INVx2_ASAP7_75t_SL g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g256 ( .A(n_207), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g325 ( .A(n_207), .B(n_260), .Y(n_325) );
BUFx2_ASAP7_75t_L g332 ( .A(n_207), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_207), .B(n_260), .Y(n_412) );
AO31x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_211), .A3(n_212), .B(n_213), .Y(n_207) );
INVx1_ASAP7_75t_L g251 ( .A(n_212), .Y(n_251) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x4_ASAP7_75t_L g342 ( .A(n_216), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g471 ( .A(n_216), .B(n_256), .Y(n_471) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx3_ASAP7_75t_L g274 ( .A(n_217), .Y(n_274) );
AND2x2_ASAP7_75t_L g285 ( .A(n_217), .B(n_260), .Y(n_285) );
AND2x2_ASAP7_75t_L g331 ( .A(n_217), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g364 ( .A(n_217), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_217), .B(n_275), .Y(n_381) );
AND2x2_ASAP7_75t_L g420 ( .A(n_217), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_225), .B(n_228), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_236), .B(n_254), .Y(n_229) );
INVx2_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_231), .A2(n_399), .B1(n_400), .B2(n_402), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_235), .Y(n_231) );
AND2x2_ASAP7_75t_L g396 ( .A(n_232), .B(n_287), .Y(n_396) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g311 ( .A(n_233), .Y(n_311) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g460 ( .A(n_234), .B(n_280), .Y(n_460) );
AND2x2_ASAP7_75t_L g424 ( .A(n_235), .B(n_319), .Y(n_424) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_252), .Y(n_236) );
OR2x2_ASAP7_75t_L g321 ( .A(n_237), .B(n_298), .Y(n_321) );
OR2x2_ASAP7_75t_L g433 ( .A(n_237), .B(n_253), .Y(n_433) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g296 ( .A(n_238), .Y(n_296) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g280 ( .A(n_239), .Y(n_280) );
BUFx3_ASAP7_75t_L g362 ( .A(n_239), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_247), .B(n_250), .Y(n_241) );
INVx2_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g430 ( .A(n_253), .B(n_289), .Y(n_430) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
AND2x2_ASAP7_75t_L g272 ( .A(n_256), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g313 ( .A(n_256), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g450 ( .A(n_256), .Y(n_450) );
INVx1_ASAP7_75t_L g469 ( .A(n_256), .Y(n_469) );
INVx2_ASAP7_75t_L g284 ( .A(n_257), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_257), .B(n_260), .Y(n_333) );
INVx1_ASAP7_75t_L g397 ( .A(n_258), .Y(n_397) );
BUFx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g458 ( .A(n_259), .Y(n_458) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g275 ( .A(n_260), .Y(n_275) );
INVx1_ASAP7_75t_L g365 ( .A(n_260), .Y(n_365) );
AO31x2_ASAP7_75t_L g485 ( .A1(n_267), .A2(n_486), .A3(n_487), .B(n_491), .Y(n_485) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_SL g518 ( .A(n_268), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_276), .B1(n_281), .B2(n_286), .Y(n_271) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g314 ( .A(n_274), .Y(n_314) );
AND2x2_ASAP7_75t_L g316 ( .A(n_274), .B(n_301), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_274), .B(n_284), .Y(n_376) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx3_ASAP7_75t_L g307 ( .A(n_277), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_277), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g401 ( .A(n_277), .B(n_385), .Y(n_401) );
INVx1_ASAP7_75t_L g305 ( .A(n_278), .Y(n_305) );
AOI222xp33_ASAP7_75t_L g315 ( .A1(n_278), .A2(n_316), .B1(n_317), .B2(n_322), .C1(n_328), .C2(n_329), .Y(n_315) );
OAI21xp33_ASAP7_75t_SL g345 ( .A1(n_278), .A2(n_346), .B(n_347), .Y(n_345) );
AND2x2_ASAP7_75t_L g369 ( .A(n_278), .B(n_288), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_278), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
OR2x2_ASAP7_75t_L g298 ( .A(n_279), .B(n_290), .Y(n_298) );
INVx1_ASAP7_75t_L g386 ( .A(n_279), .Y(n_386) );
BUFx2_ASAP7_75t_L g320 ( .A(n_280), .Y(n_320) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_283), .B(n_324), .Y(n_353) );
OR2x2_ASAP7_75t_L g465 ( .A(n_283), .B(n_325), .Y(n_465) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g348 ( .A(n_285), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g463 ( .A(n_285), .Y(n_463) );
OAI31xp33_ASAP7_75t_L g444 ( .A1(n_286), .A2(n_445), .A3(n_447), .B(n_448), .Y(n_444) );
AND2x4_ASAP7_75t_SL g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_287), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_315), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_301), .B(n_303), .Y(n_293) );
NOR2x1_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x6_ASAP7_75t_L g414 ( .A(n_296), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g346 ( .A(n_299), .Y(n_346) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g437 ( .A(n_300), .B(n_374), .Y(n_437) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_302), .A2(n_391), .B1(n_393), .B2(n_395), .Y(n_390) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_302), .A2(n_363), .B(n_425), .C(n_452), .Y(n_451) );
AOI21xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_308), .B(n_312), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_307), .B(n_405), .C(n_406), .D(n_408), .Y(n_404) );
NAND2x1_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_309), .B(n_311), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_309), .B(n_394), .Y(n_417) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g383 ( .A(n_314), .B(n_343), .Y(n_383) );
NAND2xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_321), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_321), .A2(n_465), .B1(n_466), .B2(n_468), .Y(n_464) );
AOI221x1_ASAP7_75t_L g403 ( .A1(n_322), .A2(n_404), .B1(n_410), .B2(n_413), .C(n_416), .Y(n_403) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g343 ( .A(n_325), .Y(n_343) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g355 ( .A(n_327), .B(n_356), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g418 ( .A(n_328), .B(n_409), .Y(n_418) );
O2A1O1Ixp5_ASAP7_75t_L g431 ( .A1(n_329), .A2(n_413), .B(n_432), .C(n_434), .Y(n_431) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx2_ASAP7_75t_L g380 ( .A(n_332), .Y(n_380) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_344), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_336), .A2(n_354), .B1(n_424), .B2(n_425), .C(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g360 ( .A(n_338), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_338), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g459 ( .A(n_338), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
NAND2x1_ASAP7_75t_L g438 ( .A(n_341), .B(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g462 ( .A(n_341), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g402 ( .A(n_342), .Y(n_402) );
AOI222xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_348), .B1(n_351), .B2(n_352), .C1(n_354), .C2(n_357), .Y(n_344) );
INVx1_ASAP7_75t_L g429 ( .A(n_348), .Y(n_429) );
INVx1_ASAP7_75t_L g392 ( .A(n_349), .Y(n_392) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g426 ( .A(n_350), .Y(n_426) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g367 ( .A(n_356), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g421 ( .A(n_356), .Y(n_421) );
AND2x2_ASAP7_75t_L g384 ( .A(n_357), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_377), .Y(n_358) );
AOI222xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .B1(n_366), .B2(n_369), .C1(n_370), .C2(n_375), .Y(n_359) );
INVx3_ASAP7_75t_L g409 ( .A(n_362), .Y(n_409) );
BUFx2_ASAP7_75t_L g467 ( .A(n_362), .Y(n_467) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g439 ( .A(n_364), .Y(n_439) );
OR2x2_ASAP7_75t_L g449 ( .A(n_364), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx2_ASAP7_75t_SL g407 ( .A(n_372), .Y(n_407) );
AND2x2_ASAP7_75t_L g452 ( .A(n_373), .B(n_409), .Y(n_452) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_374), .Y(n_405) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g411 ( .A(n_376), .B(n_412), .Y(n_411) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_378), .B(n_382), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
OR2x2_ASAP7_75t_L g468 ( .A(n_381), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g399 ( .A(n_383), .Y(n_399) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g406 ( .A(n_386), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g456 ( .A(n_386), .Y(n_456) );
NAND4xp75_ASAP7_75t_L g387 ( .A(n_388), .B(n_422), .C(n_440), .D(n_453), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_403), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_397), .B(n_398), .Y(n_389) );
INVxp33_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_392), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g415 ( .A(n_394), .Y(n_415) );
AND2x2_ASAP7_75t_L g455 ( .A(n_394), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g425 ( .A(n_397), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g443 ( .A(n_408), .Y(n_443) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI22xp33_ASAP7_75t_SL g434 ( .A1(n_411), .A2(n_435), .B1(n_437), .B2(n_438), .Y(n_434) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI21xp33_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_418), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g447 ( .A(n_418), .Y(n_447) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_431), .Y(n_422) );
AOI21xp5_ASAP7_75t_SL g427 ( .A1(n_428), .A2(n_429), .B(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_470), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_457), .B1(n_459), .B2(n_461), .C(n_464), .Y(n_454) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx12f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g837 ( .A(n_476), .B(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g816 ( .A(n_477), .Y(n_816) );
NAND4xp75_ASAP7_75t_L g478 ( .A(n_479), .B(n_621), .C(n_697), .D(n_749), .Y(n_478) );
NAND4xp25_ASAP7_75t_L g821 ( .A(n_479), .B(n_621), .C(n_697), .D(n_749), .Y(n_821) );
AND3x1_ASAP7_75t_L g479 ( .A(n_480), .B(n_594), .C(n_607), .Y(n_479) );
AOI221x1_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_528), .B1(n_555), .B2(n_559), .C(n_571), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_481), .A2(n_595), .B(n_597), .C(n_598), .Y(n_594) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_493), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g558 ( .A(n_485), .Y(n_558) );
BUFx2_ASAP7_75t_L g576 ( .A(n_485), .Y(n_576) );
OR2x2_ASAP7_75t_L g618 ( .A(n_485), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g625 ( .A(n_485), .B(n_496), .Y(n_625) );
AND2x4_ASAP7_75t_L g660 ( .A(n_485), .B(n_495), .Y(n_660) );
OR2x2_ASAP7_75t_L g703 ( .A(n_485), .B(n_521), .Y(n_703) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_506), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_495), .B(n_574), .Y(n_573) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_495), .Y(n_590) );
INVx2_ASAP7_75t_L g617 ( .A(n_495), .Y(n_617) );
INVx3_ASAP7_75t_L g630 ( .A(n_495), .Y(n_630) );
AND2x2_ASAP7_75t_L g748 ( .A(n_495), .B(n_577), .Y(n_748) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g557 ( .A(n_496), .B(n_558), .Y(n_557) );
BUFx2_ASAP7_75t_L g613 ( .A(n_496), .Y(n_613) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g633 ( .A(n_507), .Y(n_633) );
INVx1_ASAP7_75t_L g760 ( .A(n_507), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_520), .Y(n_507) );
AND2x2_ASAP7_75t_L g556 ( .A(n_508), .B(n_521), .Y(n_556) );
INVx1_ASAP7_75t_L g619 ( .A(n_508), .Y(n_619) );
OAI21x1_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_519), .Y(n_508) );
OAI21x1_ASAP7_75t_L g578 ( .A1(n_509), .A2(n_510), .B(n_519), .Y(n_578) );
OAI21x1_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_514), .B(n_518), .Y(n_510) );
INVx2_ASAP7_75t_L g574 ( .A(n_520), .Y(n_574) );
AND2x2_ASAP7_75t_L g626 ( .A(n_520), .B(n_577), .Y(n_626) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g588 ( .A(n_521), .Y(n_588) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_521), .Y(n_648) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_530), .A2(n_620), .B1(n_624), .B2(n_627), .Y(n_623) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_539), .Y(n_530) );
INVx1_ASAP7_75t_L g641 ( .A(n_531), .Y(n_641) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g561 ( .A(n_532), .B(n_541), .Y(n_561) );
AND2x2_ASAP7_75t_L g592 ( .A(n_532), .B(n_548), .Y(n_592) );
INVx4_ASAP7_75t_SL g603 ( .A(n_532), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_532), .B(n_637), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_532), .B(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g674 ( .A(n_540), .B(n_652), .Y(n_674) );
OR2x2_ASAP7_75t_L g707 ( .A(n_540), .B(n_689), .Y(n_707) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_548), .Y(n_540) );
INVx2_ASAP7_75t_L g581 ( .A(n_541), .Y(n_581) );
INVx1_ASAP7_75t_L g586 ( .A(n_541), .Y(n_586) );
AND2x2_ASAP7_75t_L g593 ( .A(n_541), .B(n_563), .Y(n_593) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_541), .Y(n_609) );
INVx1_ASAP7_75t_L g637 ( .A(n_541), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_541), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g570 ( .A(n_548), .Y(n_570) );
AND2x4_ASAP7_75t_L g580 ( .A(n_548), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g606 ( .A(n_548), .Y(n_606) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_548), .Y(n_683) );
INVx1_ASAP7_75t_L g776 ( .A(n_548), .Y(n_776) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_556), .B(n_629), .Y(n_696) );
AND2x2_ASAP7_75t_L g709 ( .A(n_556), .B(n_625), .Y(n_709) );
AND2x2_ASAP7_75t_L g779 ( .A(n_556), .B(n_630), .Y(n_779) );
AND2x4_ASAP7_75t_L g614 ( .A(n_558), .B(n_577), .Y(n_614) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AND2x2_ASAP7_75t_L g681 ( .A(n_561), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g695 ( .A(n_561), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_561), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g597 ( .A(n_562), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_562), .B(n_635), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g691 ( .A1(n_562), .A2(n_692), .B(n_695), .C(n_696), .Y(n_691) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_570), .Y(n_562) );
AND2x2_ASAP7_75t_L g662 ( .A(n_563), .B(n_603), .Y(n_662) );
INVx3_ASAP7_75t_L g689 ( .A(n_563), .Y(n_689) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g584 ( .A(n_564), .Y(n_584) );
AND2x4_ASAP7_75t_L g610 ( .A(n_564), .B(n_570), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_570), .B(n_603), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_579), .B1(n_587), .B2(n_591), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
INVx1_ASAP7_75t_L g728 ( .A(n_573), .Y(n_728) );
AND2x4_ASAP7_75t_L g639 ( .A(n_574), .B(n_619), .Y(n_639) );
INVx1_ASAP7_75t_L g659 ( .A(n_574), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_576), .A2(n_632), .B1(n_642), .B2(n_644), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_576), .B(n_633), .Y(n_690) );
NAND2x1_ASAP7_75t_L g747 ( .A(n_576), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g762 ( .A(n_576), .Y(n_762) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx2_ASAP7_75t_L g701 ( .A(n_578), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
AND2x2_ASAP7_75t_L g620 ( .A(n_580), .B(n_602), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_580), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g661 ( .A(n_580), .B(n_662), .Y(n_661) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_580), .Y(n_735) );
NAND2x1p5_ASAP7_75t_L g742 ( .A(n_580), .B(n_643), .Y(n_742) );
AND2x4_ASAP7_75t_L g765 ( .A(n_580), .B(n_693), .Y(n_765) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx3_ASAP7_75t_L g643 ( .A(n_583), .Y(n_643) );
AND2x2_ASAP7_75t_L g655 ( .A(n_583), .B(n_648), .Y(n_655) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g605 ( .A(n_584), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g653 ( .A(n_584), .Y(n_653) );
INVx1_ASAP7_75t_L g596 ( .A(n_585), .Y(n_596) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g753 ( .A(n_586), .B(n_603), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
AND2x2_ASAP7_75t_L g679 ( .A(n_588), .B(n_660), .Y(n_679) );
INVx2_ASAP7_75t_L g720 ( .A(n_588), .Y(n_720) );
AND2x4_ASAP7_75t_L g721 ( .A(n_588), .B(n_614), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_589), .B(n_639), .Y(n_769) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_592), .B(n_652), .Y(n_651) );
AND2x4_ASAP7_75t_L g664 ( .A(n_592), .B(n_609), .Y(n_664) );
INVx1_ASAP7_75t_L g756 ( .A(n_592), .Y(n_756) );
AND2x2_ASAP7_75t_L g755 ( .A(n_593), .B(n_682), .Y(n_755) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g726 ( .A1(n_597), .A2(n_727), .B1(n_729), .B2(n_731), .Y(n_726) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g635 ( .A(n_603), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g671 ( .A(n_603), .Y(n_671) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_603), .Y(n_677) );
INVx2_ASAP7_75t_L g694 ( .A(n_603), .Y(n_694) );
OR2x2_ASAP7_75t_L g715 ( .A(n_603), .B(n_678), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_603), .B(n_673), .Y(n_725) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g692 ( .A(n_605), .B(n_693), .Y(n_692) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_605), .Y(n_746) );
INVx1_ASAP7_75t_L g673 ( .A(n_606), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_611), .B(n_615), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_610), .B(n_641), .Y(n_640) );
INVx3_ASAP7_75t_L g678 ( .A(n_610), .Y(n_678) );
AND2x2_ASAP7_75t_L g752 ( .A(n_610), .B(n_753), .Y(n_752) );
AOI211x1_ASAP7_75t_SL g680 ( .A1(n_611), .A2(n_681), .B(n_684), .C(n_691), .Y(n_680) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_L g737 ( .A(n_613), .B(n_614), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_614), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_614), .Y(n_730) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_620), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g645 ( .A(n_617), .Y(n_645) );
NOR2x1p5_ASAP7_75t_L g702 ( .A(n_617), .B(n_703), .Y(n_702) );
NOR2x1_ASAP7_75t_L g646 ( .A(n_618), .B(n_647), .Y(n_646) );
NOR2xp67_ASAP7_75t_SL g719 ( .A(n_618), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g780 ( .A(n_620), .B(n_688), .Y(n_780) );
NOR2x1_ASAP7_75t_L g621 ( .A(n_622), .B(n_665), .Y(n_621) );
NAND3xp33_ASAP7_75t_SL g622 ( .A(n_623), .B(n_631), .C(n_649), .Y(n_622) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_625), .Y(n_656) );
AND2x2_ASAP7_75t_L g663 ( .A(n_625), .B(n_659), .Y(n_663) );
AND2x4_ASAP7_75t_SL g777 ( .A(n_625), .B(n_639), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_626), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_628), .A2(n_670), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x4_ASAP7_75t_L g759 ( .A(n_630), .B(n_760), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_638), .B2(n_640), .Y(n_632) );
NAND2x1_ASAP7_75t_L g708 ( .A(n_635), .B(n_688), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_635), .B(n_682), .Y(n_718) );
INVx1_ASAP7_75t_L g745 ( .A(n_635), .Y(n_745) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_638), .A2(n_764), .B(n_767), .Y(n_763) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_639), .A2(n_651), .B(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g724 ( .A(n_643), .Y(n_724) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g668 ( .A(n_646), .Y(n_668) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI222xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_656), .B1(n_657), .B2(n_661), .C1(n_663), .C2(n_664), .Y(n_649) );
AOI21xp33_ASAP7_75t_L g684 ( .A1(n_651), .A2(n_685), .B(n_690), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_652), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g766 ( .A(n_652), .Y(n_766) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_653), .Y(n_772) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
AND2x2_ASAP7_75t_L g736 ( .A(n_658), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g729 ( .A(n_659), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_680), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B1(n_675), .B2(n_679), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_674), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx1_ASAP7_75t_L g686 ( .A(n_672), .Y(n_686) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx4_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g714 ( .A(n_689), .B(n_706), .Y(n_714) );
OR2x2_ASAP7_75t_L g774 ( .A(n_689), .B(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND5xp2_ASAP7_75t_L g750 ( .A(n_695), .B(n_742), .C(n_751), .D(n_754), .E(n_756), .Y(n_750) );
NOR2x1_ASAP7_75t_L g697 ( .A(n_698), .B(n_733), .Y(n_697) );
NAND2xp67_ASAP7_75t_SL g698 ( .A(n_699), .B(n_716), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_704), .B1(n_709), .B2(n_710), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
NAND3xp33_ASAP7_75t_SL g704 ( .A(n_705), .B(n_707), .C(n_708), .Y(n_704) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g739 ( .A(n_708), .Y(n_739) );
NAND3xp33_ASAP7_75t_SL g710 ( .A(n_711), .B(n_714), .C(n_715), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g732 ( .A(n_713), .Y(n_732) );
O2A1O1Ixp33_ASAP7_75t_SL g744 ( .A1(n_714), .A2(n_745), .B(n_746), .C(n_747), .Y(n_744) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_719), .B1(n_721), .B2(n_722), .C(n_726), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_723), .B(n_771), .Y(n_770) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g740 ( .A(n_727), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_738), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g743 ( .A(n_737), .Y(n_743) );
AOI211xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B(n_741), .C(n_744), .Y(n_738) );
AOI211x1_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_757), .B(n_763), .C(n_778), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2x1p5_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2x1_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_770), .B1(n_773), .B2(n_777), .Y(n_767) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AND2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
CKINVDCx6p67_ASAP7_75t_R g791 ( .A(n_783), .Y(n_791) );
BUFx3_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
BUFx6f_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
AND2x6_ASAP7_75t_SL g795 ( .A(n_796), .B(n_798), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx3_ASAP7_75t_L g808 ( .A(n_797), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_797), .B(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_801), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NOR2x1_ASAP7_75t_L g838 ( .A(n_800), .B(n_802), .Y(n_838) );
AND3x2_ASAP7_75t_L g813 ( .A(n_801), .B(n_814), .C(n_816), .Y(n_813) );
AND2x6_ASAP7_75t_SL g827 ( .A(n_801), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OAI21x1_ASAP7_75t_SL g803 ( .A1(n_804), .A2(n_809), .B(n_831), .Y(n_803) );
INVx4_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
BUFx6f_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AOI22x1_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_822), .B1(n_826), .B2(n_830), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_817), .Y(n_810) );
BUFx2_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
INVx4_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g841 ( .A(n_813), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_814), .B(n_850), .Y(n_849) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g829 ( .A(n_815), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_816), .B(n_852), .Y(n_851) );
INVxp67_ASAP7_75t_SL g830 ( .A(n_817), .Y(n_830) );
XNOR2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_821), .Y(n_817) );
NOR2xp33_ASAP7_75t_R g826 ( .A(n_822), .B(n_827), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_823), .Y(n_825) );
INVx3_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx6_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
BUFx10_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NOR2xp33_ASAP7_75t_SL g839 ( .A(n_840), .B(n_841), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_843), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_844), .Y(n_843) );
CKINVDCx11_ASAP7_75t_R g856 ( .A(n_844), .Y(n_856) );
BUFx12f_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NOR2x1p5_ASAP7_75t_L g845 ( .A(n_846), .B(n_849), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_855), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g855 ( .A(n_856), .Y(n_855) );
endmodule