module fake_jpeg_20010_n_95 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_41),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_40),
.B1(n_45),
.B2(n_43),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_39),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_36),
.B(n_34),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_38),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_67)
);

OAI32xp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_73),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_3),
.Y(n_77)
);

NAND2x1_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_1),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_4),
.B1(n_69),
.B2(n_74),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_14),
.B1(n_29),
.B2(n_28),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_12),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_7),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_8),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_71),
.C(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_85),
.B(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_82),
.C(n_86),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_83),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_13),
.C(n_19),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_20),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_22),
.C(n_23),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_24),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_25),
.Y(n_95)
);


endmodule