module real_aes_10805_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_1404;
wire n_602;
wire n_402;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1699;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1691;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1369;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVxp67_ASAP7_75t_L g381 ( .A(n_0), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_0), .A2(n_7), .B1(n_484), .B2(n_488), .Y(n_483) );
XNOR2x2_ASAP7_75t_L g322 ( .A(n_1), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1), .Y(n_1469) );
AOI21xp33_ASAP7_75t_L g1209 ( .A1(n_2), .A2(n_485), .B(n_957), .Y(n_1209) );
INVx1_ASAP7_75t_L g1230 ( .A(n_2), .Y(n_1230) );
INVxp67_ASAP7_75t_L g384 ( .A(n_3), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_3), .A2(n_83), .B1(n_446), .B2(n_475), .C(n_480), .Y(n_474) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_4), .Y(n_311) );
AND2x2_ASAP7_75t_L g335 ( .A(n_4), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_4), .B(n_223), .Y(n_367) );
INVx1_ASAP7_75t_L g415 ( .A(n_4), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g1346 ( .A1(n_5), .A2(n_155), .B1(n_1347), .B2(n_1348), .Y(n_1346) );
INVx1_ASAP7_75t_L g1366 ( .A(n_5), .Y(n_1366) );
INVxp67_ASAP7_75t_L g549 ( .A(n_6), .Y(n_549) );
OAI222xp33_ASAP7_75t_L g570 ( .A1(n_6), .A2(n_49), .B1(n_281), .B2(n_571), .C1(n_573), .C2(n_575), .Y(n_570) );
INVxp67_ASAP7_75t_L g398 ( .A(n_7), .Y(n_398) );
INVx1_ASAP7_75t_L g1373 ( .A(n_8), .Y(n_1373) );
OAI221xp5_ASAP7_75t_L g1659 ( .A1(n_9), .A2(n_667), .B1(n_854), .B2(n_1660), .C(n_1664), .Y(n_1659) );
INVx1_ASAP7_75t_L g1678 ( .A(n_9), .Y(n_1678) );
XNOR2x2_ASAP7_75t_L g832 ( .A(n_10), .B(n_833), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_11), .A2(n_235), .B1(n_896), .B2(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g1006 ( .A(n_11), .Y(n_1006) );
INVxp33_ASAP7_75t_L g925 ( .A(n_12), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g959 ( .A1(n_12), .A2(n_25), .B1(n_960), .B2(n_961), .C(n_962), .Y(n_959) );
CKINVDCx5p33_ASAP7_75t_R g735 ( .A(n_13), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_14), .A2(n_196), .B1(n_779), .B2(n_1101), .C(n_1102), .Y(n_1100) );
INVx1_ASAP7_75t_L g1120 ( .A(n_14), .Y(n_1120) );
OAI221xp5_ASAP7_75t_L g325 ( .A1(n_15), .A2(n_280), .B1(n_326), .B2(n_337), .C(n_344), .Y(n_325) );
INVx1_ASAP7_75t_L g461 ( .A(n_15), .Y(n_461) );
INVx1_ASAP7_75t_L g1376 ( .A(n_16), .Y(n_1376) );
INVx1_ASAP7_75t_L g941 ( .A(n_17), .Y(n_941) );
INVx1_ASAP7_75t_L g1653 ( .A(n_18), .Y(n_1653) );
AOI22xp33_ASAP7_75t_L g1680 ( .A1(n_18), .A2(n_67), .B1(n_421), .B2(n_780), .Y(n_1680) );
AO22x2_ASAP7_75t_L g1284 ( .A1(n_19), .A2(n_1285), .B1(n_1335), .B2(n_1336), .Y(n_1284) );
CKINVDCx14_ASAP7_75t_R g1335 ( .A(n_19), .Y(n_1335) );
INVxp33_ASAP7_75t_SL g715 ( .A(n_20), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g740 ( .A1(n_20), .A2(n_113), .B1(n_619), .B2(n_741), .C(n_743), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_21), .A2(n_95), .B1(n_477), .B2(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_21), .A2(n_39), .B1(n_650), .B2(n_668), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_22), .A2(n_268), .B1(n_589), .B2(n_625), .Y(n_1109) );
INVx1_ASAP7_75t_L g1128 ( .A(n_22), .Y(n_1128) );
INVx1_ASAP7_75t_L g1528 ( .A(n_23), .Y(n_1528) );
AOI221xp5_ASAP7_75t_L g1657 ( .A1(n_24), .A2(n_66), .B1(n_340), .B2(n_680), .C(n_1003), .Y(n_1657) );
INVx1_ASAP7_75t_L g1683 ( .A(n_24), .Y(n_1683) );
INVxp67_ASAP7_75t_L g928 ( .A(n_25), .Y(n_928) );
AOI221xp5_ASAP7_75t_L g777 ( .A1(n_26), .A2(n_279), .B1(n_594), .B2(n_596), .C(n_756), .Y(n_777) );
INVx1_ASAP7_75t_L g801 ( .A(n_26), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_27), .A2(n_137), .B1(n_619), .B2(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g1017 ( .A(n_27), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g1188 ( .A1(n_28), .A2(n_1143), .B1(n_1189), .B2(n_1194), .C(n_1199), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_28), .A2(n_197), .B1(n_678), .B2(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1423 ( .A(n_29), .Y(n_1423) );
AO221x2_ASAP7_75t_L g1433 ( .A1(n_30), .A2(n_69), .B1(n_1404), .B2(n_1412), .C(n_1434), .Y(n_1433) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_31), .A2(n_163), .B1(n_676), .B2(n_678), .C(n_680), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_31), .A2(n_247), .B1(n_697), .B2(n_698), .Y(n_696) );
OR2x2_ASAP7_75t_L g426 ( .A(n_32), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g434 ( .A(n_32), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g1261 ( .A1(n_33), .A2(n_210), .B1(n_728), .B2(n_841), .C(n_1262), .Y(n_1261) );
INVx1_ASAP7_75t_L g1269 ( .A(n_33), .Y(n_1269) );
INVx1_ASAP7_75t_L g1435 ( .A(n_34), .Y(n_1435) );
AO22x1_ASAP7_75t_L g1648 ( .A1(n_34), .A2(n_1435), .B1(n_1649), .B2(n_1685), .Y(n_1648) );
AOI22xp33_ASAP7_75t_L g1690 ( .A1(n_34), .A2(n_1691), .B1(n_1695), .B2(n_1700), .Y(n_1690) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_35), .A2(n_76), .B1(n_619), .B2(n_621), .Y(n_618) );
INVx1_ASAP7_75t_L g666 ( .A(n_35), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g1048 ( .A1(n_36), .A2(n_114), .B1(n_359), .B2(n_369), .C(n_1049), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_36), .A2(n_114), .B1(n_564), .B2(n_785), .Y(n_1075) );
INVx1_ASAP7_75t_L g551 ( .A(n_37), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g1154 ( .A1(n_38), .A2(n_262), .B1(n_785), .B2(n_1155), .Y(n_1154) );
OAI221xp5_ASAP7_75t_L g1167 ( .A1(n_38), .A2(n_262), .B1(n_359), .B2(n_369), .C(n_806), .Y(n_1167) );
OAI222xp33_ASAP7_75t_L g691 ( .A1(n_39), .A2(n_163), .B1(n_169), .B2(n_512), .C1(n_692), .C2(n_695), .Y(n_691) );
INVx1_ASAP7_75t_L g334 ( .A(n_40), .Y(n_334) );
OR2x2_ASAP7_75t_L g366 ( .A(n_40), .B(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g379 ( .A(n_40), .Y(n_379) );
BUFx2_ASAP7_75t_L g514 ( .A(n_40), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_41), .Y(n_405) );
INVx1_ASAP7_75t_L g1526 ( .A(n_42), .Y(n_1526) );
INVx1_ASAP7_75t_L g1000 ( .A(n_43), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_43), .A2(n_273), .B1(n_698), .B2(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1288 ( .A(n_44), .Y(n_1288) );
AOI21xp33_ASAP7_75t_L g1326 ( .A1(n_44), .A2(n_421), .B(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1248 ( .A(n_45), .Y(n_1248) );
CKINVDCx5p33_ASAP7_75t_R g1300 ( .A(n_46), .Y(n_1300) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_47), .A2(n_150), .B1(n_421), .B2(n_780), .Y(n_1208) );
INVx1_ASAP7_75t_L g1231 ( .A(n_47), .Y(n_1231) );
INVx1_ASAP7_75t_L g530 ( .A(n_48), .Y(n_530) );
INVxp67_ASAP7_75t_L g547 ( .A(n_49), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_50), .A2(n_229), .B1(n_625), .B2(n_1147), .Y(n_1146) );
INVx1_ASAP7_75t_L g1172 ( .A(n_50), .Y(n_1172) );
OAI221xp5_ASAP7_75t_L g358 ( .A1(n_51), .A2(n_86), .B1(n_359), .B2(n_368), .C(n_373), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_51), .A2(n_86), .B1(n_429), .B2(n_440), .Y(n_428) );
INVx1_ASAP7_75t_L g935 ( .A(n_52), .Y(n_935) );
INVx1_ASAP7_75t_L g988 ( .A(n_53), .Y(n_988) );
OAI221xp5_ASAP7_75t_L g1011 ( .A1(n_53), .A2(n_854), .B1(n_866), .B2(n_1012), .C(n_1016), .Y(n_1011) );
OAI221xp5_ASAP7_75t_L g1328 ( .A1(n_54), .A2(n_242), .B1(n_440), .B2(n_1329), .C(n_1330), .Y(n_1328) );
INVx1_ASAP7_75t_L g1333 ( .A(n_54), .Y(n_1333) );
CKINVDCx16_ASAP7_75t_R g1413 ( .A(n_55), .Y(n_1413) );
INVx1_ASAP7_75t_L g1522 ( .A(n_56), .Y(n_1522) );
INVx1_ASAP7_75t_L g1663 ( .A(n_57), .Y(n_1663) );
AOI22xp33_ASAP7_75t_L g1674 ( .A1(n_57), .A2(n_160), .B1(n_780), .B2(n_951), .Y(n_1674) );
INVx1_ASAP7_75t_L g1254 ( .A(n_58), .Y(n_1254) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_59), .A2(n_63), .B1(n_839), .B2(n_841), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_59), .A2(n_79), .B1(n_697), .B2(n_698), .Y(n_905) );
OAI22xp5_ASAP7_75t_L g1658 ( .A1(n_60), .A2(n_173), .B1(n_685), .B2(n_687), .Y(n_1658) );
OAI22xp5_ASAP7_75t_SL g1671 ( .A1(n_60), .A2(n_173), .B1(n_633), .B2(n_639), .Y(n_1671) );
CKINVDCx5p33_ASAP7_75t_R g1358 ( .A(n_61), .Y(n_1358) );
INVx1_ASAP7_75t_L g641 ( .A(n_62), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_62), .A2(n_96), .B1(n_685), .B2(n_687), .C(n_688), .Y(n_684) );
INVxp67_ASAP7_75t_SL g902 ( .A(n_63), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g1210 ( .A1(n_64), .A2(n_197), .B1(n_499), .B2(n_501), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_64), .A2(n_289), .B1(n_1219), .B2(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g861 ( .A(n_65), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g1684 ( .A1(n_66), .A2(n_123), .B1(n_698), .B2(n_1027), .Y(n_1684) );
INVx1_ASAP7_75t_L g1654 ( .A(n_67), .Y(n_1654) );
CKINVDCx5p33_ASAP7_75t_R g1104 ( .A(n_68), .Y(n_1104) );
INVx1_ASAP7_75t_L g1069 ( .A(n_70), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_71), .A2(n_293), .B1(n_484), .B2(n_1350), .Y(n_1352) );
OAI22xp33_ASAP7_75t_L g1384 ( .A1(n_71), .A2(n_221), .B1(n_854), .B2(n_1385), .Y(n_1384) );
AOI221xp5_ASAP7_75t_L g1145 ( .A1(n_72), .A2(n_81), .B1(n_580), .B2(n_582), .C(n_756), .Y(n_1145) );
INVxp67_ASAP7_75t_SL g1173 ( .A(n_72), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_73), .A2(n_221), .B1(n_1354), .B2(n_1355), .Y(n_1353) );
OAI22xp33_ASAP7_75t_L g1362 ( .A1(n_73), .A2(n_293), .B1(n_836), .B2(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1446 ( .A(n_74), .Y(n_1446) );
CKINVDCx16_ASAP7_75t_R g1451 ( .A(n_75), .Y(n_1451) );
INVx1_ASAP7_75t_L g664 ( .A(n_76), .Y(n_664) );
INVxp67_ASAP7_75t_L g931 ( .A(n_77), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_77), .A2(n_222), .B1(n_621), .B2(n_964), .Y(n_963) );
CKINVDCx5p33_ASAP7_75t_R g1360 ( .A(n_78), .Y(n_1360) );
AOI221xp5_ASAP7_75t_L g843 ( .A1(n_79), .A2(n_208), .B1(n_680), .B2(n_844), .C(n_846), .Y(n_843) );
INVxp33_ASAP7_75t_SL g1054 ( .A(n_80), .Y(n_1054) );
AOI221xp5_ASAP7_75t_L g1081 ( .A1(n_80), .A2(n_106), .B1(n_753), .B2(n_1082), .C(n_1084), .Y(n_1081) );
INVxp67_ASAP7_75t_SL g1176 ( .A(n_81), .Y(n_1176) );
AOI221xp5_ASAP7_75t_L g1250 ( .A1(n_82), .A2(n_142), .B1(n_672), .B2(n_1061), .C(n_1251), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1272 ( .A1(n_82), .A2(n_101), .B1(n_1086), .B2(n_1088), .Y(n_1272) );
INVxp67_ASAP7_75t_L g392 ( .A(n_83), .Y(n_392) );
INVx1_ASAP7_75t_L g1470 ( .A(n_84), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_85), .A2(n_259), .B1(n_572), .B2(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g802 ( .A(n_85), .Y(n_802) );
INVx1_ASAP7_75t_L g1253 ( .A(n_87), .Y(n_1253) );
AOI221xp5_ASAP7_75t_L g1271 ( .A1(n_87), .A2(n_142), .B1(n_1077), .B2(n_1082), .C(n_1084), .Y(n_1271) );
INVxp33_ASAP7_75t_L g1043 ( .A(n_88), .Y(n_1043) );
AOI221xp5_ASAP7_75t_L g1076 ( .A1(n_88), .A2(n_296), .B1(n_779), .B2(n_1077), .C(n_1078), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_89), .A2(n_157), .B1(n_592), .B2(n_594), .C(n_596), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g600 ( .A1(n_89), .A2(n_176), .B1(n_601), .B2(n_602), .C(n_604), .Y(n_600) );
CKINVDCx16_ASAP7_75t_R g1454 ( .A(n_90), .Y(n_1454) );
AOI22xp5_ASAP7_75t_L g1426 ( .A1(n_91), .A2(n_147), .B1(n_1427), .B2(n_1430), .Y(n_1426) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_92), .A2(n_244), .B1(n_723), .B2(n_729), .Y(n_731) );
INVxp33_ASAP7_75t_L g765 ( .A(n_92), .Y(n_765) );
INVx1_ASAP7_75t_L g427 ( .A(n_93), .Y(n_427) );
INVx1_ASAP7_75t_L g466 ( .A(n_93), .Y(n_466) );
INVx1_ASAP7_75t_L g1140 ( .A(n_94), .Y(n_1140) );
INVx1_ASAP7_75t_L g683 ( .A(n_95), .Y(n_683) );
INVx1_ASAP7_75t_L g637 ( .A(n_96), .Y(n_637) );
AOI22xp33_ASAP7_75t_SL g1696 ( .A1(n_97), .A2(n_1697), .B1(n_1698), .B2(n_1699), .Y(n_1696) );
CKINVDCx5p33_ASAP7_75t_R g1697 ( .A(n_97), .Y(n_1697) );
INVx1_ASAP7_75t_L g1263 ( .A(n_98), .Y(n_1263) );
OAI221xp5_ASAP7_75t_L g1267 ( .A1(n_98), .A2(n_210), .B1(n_573), .B2(n_881), .C(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1195 ( .A(n_99), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_99), .A2(n_172), .B1(n_678), .B2(n_1217), .Y(n_1216) );
INVxp33_ASAP7_75t_L g916 ( .A(n_100), .Y(n_916) );
AOI221xp5_ASAP7_75t_L g948 ( .A1(n_100), .A2(n_194), .B1(n_949), .B2(n_952), .C(n_953), .Y(n_948) );
INVxp67_ASAP7_75t_SL g1252 ( .A(n_101), .Y(n_1252) );
INVx1_ASAP7_75t_L g712 ( .A(n_102), .Y(n_712) );
INVx1_ASAP7_75t_L g1259 ( .A(n_103), .Y(n_1259) );
AOI221xp5_ASAP7_75t_L g1274 ( .A1(n_103), .A2(n_154), .B1(n_879), .B2(n_1275), .C(n_1276), .Y(n_1274) );
INVx1_ASAP7_75t_L g864 ( .A(n_104), .Y(n_864) );
AOI221xp5_ASAP7_75t_L g875 ( .A1(n_104), .A2(n_285), .B1(n_876), .B2(n_878), .C(n_880), .Y(n_875) );
XNOR2xp5_ASAP7_75t_L g519 ( .A(n_105), .B(n_520), .Y(n_519) );
INVxp67_ASAP7_75t_SL g1058 ( .A(n_106), .Y(n_1058) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_107), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_108), .A2(n_1185), .B1(n_1235), .B2(n_1236), .Y(n_1184) );
INVxp67_ASAP7_75t_SL g1235 ( .A(n_108), .Y(n_1235) );
INVxp67_ASAP7_75t_L g528 ( .A(n_109), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_109), .A2(n_179), .B1(n_580), .B2(n_581), .C(n_582), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_110), .A2(n_175), .B1(n_594), .B2(n_623), .Y(n_622) );
AOI21xp33_ASAP7_75t_L g660 ( .A1(n_110), .A2(n_377), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g714 ( .A(n_111), .Y(n_714) );
OAI21xp33_ASAP7_75t_L g1244 ( .A1(n_112), .A2(n_1245), .B(n_1265), .Y(n_1244) );
INVx1_ASAP7_75t_L g1282 ( .A(n_112), .Y(n_1282) );
INVx1_ASAP7_75t_L g1420 ( .A(n_112), .Y(n_1420) );
INVxp33_ASAP7_75t_L g711 ( .A(n_113), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_115), .A2(n_243), .B1(n_481), .B2(n_753), .C(n_756), .Y(n_787) );
INVx1_ASAP7_75t_L g818 ( .A(n_115), .Y(n_818) );
AOI22xp33_ASAP7_75t_SL g722 ( .A1(n_116), .A2(n_263), .B1(n_723), .B2(n_724), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_116), .A2(n_263), .B1(n_761), .B2(n_763), .Y(n_760) );
INVx1_ASAP7_75t_L g1264 ( .A(n_117), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_118), .A2(n_254), .B1(n_1152), .B2(n_1153), .Y(n_1151) );
INVx1_ASAP7_75t_L g1166 ( .A(n_118), .Y(n_1166) );
AO221x2_ASAP7_75t_L g1467 ( .A1(n_119), .A2(n_200), .B1(n_1412), .B2(n_1453), .C(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g345 ( .A(n_120), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_121), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g1462 ( .A1(n_122), .A2(n_231), .B1(n_1453), .B2(n_1463), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g1656 ( .A1(n_123), .A2(n_135), .B1(n_673), .B2(n_728), .Y(n_1656) );
AOI221xp5_ASAP7_75t_L g1150 ( .A1(n_124), .A2(n_236), .B1(n_485), .B2(n_756), .C(n_957), .Y(n_1150) );
INVx1_ASAP7_75t_L g1165 ( .A(n_124), .Y(n_1165) );
INVx1_ASAP7_75t_L g969 ( .A(n_125), .Y(n_969) );
INVx1_ASAP7_75t_L g303 ( .A(n_126), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g1111 ( .A(n_127), .Y(n_1111) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_128), .Y(n_793) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_129), .A2(n_177), .B1(n_724), .B2(n_727), .Y(n_730) );
INVxp33_ASAP7_75t_L g766 ( .A(n_129), .Y(n_766) );
OA22x2_ASAP7_75t_L g771 ( .A1(n_130), .A2(n_772), .B1(n_828), .B2(n_829), .Y(n_771) );
INVx1_ASAP7_75t_L g829 ( .A(n_130), .Y(n_829) );
INVx1_ASAP7_75t_L g913 ( .A(n_131), .Y(n_913) );
CKINVDCx5p33_ASAP7_75t_R g966 ( .A(n_132), .Y(n_966) );
CKINVDCx5p33_ASAP7_75t_R g1297 ( .A(n_133), .Y(n_1297) );
OAI221xp5_ASAP7_75t_SL g1257 ( .A1(n_134), .A2(n_260), .B1(n_663), .B2(n_860), .C(n_1258), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_134), .A2(n_260), .B1(n_951), .B2(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1682 ( .A(n_135), .Y(n_1682) );
AOI22xp5_ASAP7_75t_L g1432 ( .A1(n_136), .A2(n_193), .B1(n_1404), .B2(n_1412), .Y(n_1432) );
INVx1_ASAP7_75t_L g1020 ( .A(n_137), .Y(n_1020) );
INVx1_ASAP7_75t_L g907 ( .A(n_138), .Y(n_907) );
INVx1_ASAP7_75t_L g869 ( .A(n_139), .Y(n_869) );
OAI222xp33_ASAP7_75t_L g522 ( .A1(n_140), .A2(n_180), .B1(n_286), .B2(n_511), .C1(n_523), .C2(n_525), .Y(n_522) );
INVx1_ASAP7_75t_L g562 ( .A(n_140), .Y(n_562) );
INVx1_ASAP7_75t_L g1070 ( .A(n_141), .Y(n_1070) );
INVx1_ASAP7_75t_L g1436 ( .A(n_143), .Y(n_1436) );
CKINVDCx5p33_ASAP7_75t_R g1665 ( .A(n_144), .Y(n_1665) );
CKINVDCx5p33_ASAP7_75t_R g1302 ( .A(n_145), .Y(n_1302) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_146), .Y(n_792) );
XNOR2xp5_ASAP7_75t_L g610 ( .A(n_147), .B(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_SL g726 ( .A1(n_148), .A2(n_151), .B1(n_727), .B2(n_729), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_148), .A2(n_151), .B1(n_753), .B2(n_754), .C(n_757), .Y(n_752) );
CKINVDCx5p33_ASAP7_75t_R g1204 ( .A(n_149), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g1232 ( .A1(n_150), .A2(n_275), .B1(n_1233), .B2(n_1234), .Y(n_1232) );
INVx1_ASAP7_75t_L g1064 ( .A(n_152), .Y(n_1064) );
AOI221xp5_ASAP7_75t_L g1107 ( .A1(n_153), .A2(n_288), .B1(n_580), .B2(n_1084), .C(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1127 ( .A(n_153), .Y(n_1127) );
INVx1_ASAP7_75t_L g1260 ( .A(n_154), .Y(n_1260) );
INVx1_ASAP7_75t_L g1367 ( .A(n_155), .Y(n_1367) );
INVx1_ASAP7_75t_L g999 ( .A(n_156), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_156), .A2(n_264), .B1(n_692), .B2(n_695), .Y(n_1028) );
OAI332xp33_ASAP7_75t_L g526 ( .A1(n_157), .A2(n_376), .A3(n_527), .B1(n_533), .B2(n_540), .B3(n_548), .C1(n_552), .C2(n_554), .Y(n_526) );
INVx1_ASAP7_75t_L g1290 ( .A(n_158), .Y(n_1290) );
AOI22xp33_ASAP7_75t_SL g1324 ( .A1(n_158), .A2(n_217), .B1(n_780), .B2(n_1325), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g1308 ( .A1(n_159), .A2(n_207), .B1(n_554), .B2(n_1309), .Y(n_1308) );
INVx1_ASAP7_75t_L g1318 ( .A(n_159), .Y(n_1318) );
INVx1_ASAP7_75t_L g1661 ( .A(n_160), .Y(n_1661) );
CKINVDCx5p33_ASAP7_75t_R g1097 ( .A(n_161), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_162), .A2(n_188), .B1(n_685), .B2(n_687), .Y(n_849) );
OAI221xp5_ASAP7_75t_L g893 ( .A1(n_162), .A2(n_188), .B1(n_894), .B2(n_896), .C(n_897), .Y(n_893) );
INVxp67_ASAP7_75t_SL g705 ( .A(n_164), .Y(n_705) );
OAI22xp33_ASAP7_75t_L g739 ( .A1(n_164), .A2(n_274), .B1(n_429), .B2(n_440), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g1310 ( .A1(n_165), .A2(n_239), .B1(n_511), .B2(n_1233), .Y(n_1310) );
AOI22xp33_ASAP7_75t_SL g1319 ( .A1(n_165), .A2(n_207), .B1(n_421), .B2(n_780), .Y(n_1319) );
INVx1_ASAP7_75t_L g1144 ( .A(n_166), .Y(n_1144) );
XNOR2xp5_ASAP7_75t_L g1092 ( .A(n_167), .B(n_1093), .Y(n_1092) );
AOI22xp5_ASAP7_75t_L g1461 ( .A1(n_167), .A2(n_212), .B1(n_1427), .B2(n_1430), .Y(n_1461) );
CKINVDCx5p33_ASAP7_75t_R g1377 ( .A(n_168), .Y(n_1377) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_169), .A2(n_247), .B1(n_672), .B2(n_673), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_170), .A2(n_294), .B1(n_447), .B2(n_628), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g1021 ( .A1(n_170), .A2(n_294), .B1(n_1022), .B2(n_1023), .Y(n_1021) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_171), .Y(n_402) );
INVx1_ASAP7_75t_L g1191 ( .A(n_172), .Y(n_1191) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_174), .A2(n_182), .B1(n_448), .B2(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g653 ( .A(n_174), .Y(n_653) );
INVx1_ASAP7_75t_L g659 ( .A(n_175), .Y(n_659) );
INVx1_ASAP7_75t_L g590 ( .A(n_176), .Y(n_590) );
INVxp67_ASAP7_75t_SL g738 ( .A(n_177), .Y(n_738) );
INVx1_ASAP7_75t_L g942 ( .A(n_178), .Y(n_942) );
INVx1_ASAP7_75t_L g534 ( .A(n_179), .Y(n_534) );
INVx1_ASAP7_75t_L g587 ( .A(n_180), .Y(n_587) );
INVxp33_ASAP7_75t_L g1052 ( .A(n_181), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_181), .A2(n_216), .B1(n_1086), .B2(n_1088), .Y(n_1085) );
INVx1_ASAP7_75t_L g655 ( .A(n_182), .Y(n_655) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_183), .Y(n_305) );
AND3x2_ASAP7_75t_L g1405 ( .A(n_183), .B(n_303), .C(n_1406), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1417 ( .A(n_183), .B(n_303), .Y(n_1417) );
INVx1_ASAP7_75t_L g1090 ( .A(n_184), .Y(n_1090) );
OAI22xp33_ASAP7_75t_SL g1098 ( .A1(n_185), .A2(n_203), .B1(n_564), .B2(n_1099), .Y(n_1098) );
OAI221xp5_ASAP7_75t_L g1121 ( .A1(n_185), .A2(n_203), .B1(n_359), .B2(n_369), .C(n_1049), .Y(n_1121) );
AOI21xp33_ASAP7_75t_L g1198 ( .A1(n_186), .A2(n_481), .B(n_951), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1218 ( .A1(n_186), .A2(n_272), .B1(n_1219), .B2(n_1221), .Y(n_1218) );
OAI221xp5_ASAP7_75t_L g918 ( .A1(n_187), .A2(n_225), .B1(n_525), .B2(n_806), .C(n_919), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_187), .A2(n_225), .B1(n_440), .B2(n_947), .Y(n_946) );
CKINVDCx5p33_ASAP7_75t_R g972 ( .A(n_189), .Y(n_972) );
CKINVDCx5p33_ASAP7_75t_R g1298 ( .A(n_190), .Y(n_1298) );
INVx2_ASAP7_75t_L g316 ( .A(n_191), .Y(n_316) );
INVx1_ASAP7_75t_L g1157 ( .A(n_192), .Y(n_1157) );
INVxp33_ASAP7_75t_L g912 ( .A(n_194), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_195), .A2(n_269), .B1(n_449), .B2(n_594), .Y(n_788) );
INVx1_ASAP7_75t_L g812 ( .A(n_195), .Y(n_812) );
INVx1_ASAP7_75t_L g1117 ( .A(n_196), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_198), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g1457 ( .A1(n_199), .A2(n_209), .B1(n_1404), .B2(n_1412), .Y(n_1457) );
OAI211xp5_ASAP7_75t_L g1651 ( .A1(n_201), .A2(n_836), .B(n_1652), .C(n_1655), .Y(n_1651) );
INVx1_ASAP7_75t_L g1679 ( .A(n_201), .Y(n_1679) );
INVx1_ASAP7_75t_L g1247 ( .A(n_202), .Y(n_1247) );
CKINVDCx5p33_ASAP7_75t_R g1203 ( .A(n_204), .Y(n_1203) );
INVx1_ASAP7_75t_L g859 ( .A(n_205), .Y(n_859) );
INVx1_ASAP7_75t_L g1406 ( .A(n_206), .Y(n_1406) );
INVxp67_ASAP7_75t_SL g904 ( .A(n_208), .Y(n_904) );
CKINVDCx16_ASAP7_75t_R g1410 ( .A(n_211), .Y(n_1410) );
INVx1_ASAP7_75t_L g1524 ( .A(n_213), .Y(n_1524) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_214), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g982 ( .A(n_215), .Y(n_982) );
INVxp67_ASAP7_75t_SL g1059 ( .A(n_216), .Y(n_1059) );
INVx1_ASAP7_75t_L g1294 ( .A(n_217), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g1349 ( .A1(n_218), .A2(n_265), .B1(n_484), .B2(n_1350), .Y(n_1349) );
INVx1_ASAP7_75t_L g1371 ( .A(n_218), .Y(n_1371) );
OAI211xp5_ASAP7_75t_L g835 ( .A1(n_219), .A2(n_836), .B(n_837), .C(n_850), .Y(n_835) );
AOI221xp5_ASAP7_75t_L g884 ( .A1(n_219), .A2(n_227), .B1(n_484), .B2(n_885), .C(n_887), .Y(n_884) );
INVx1_ASAP7_75t_L g915 ( .A(n_220), .Y(n_915) );
INVxp33_ASAP7_75t_L g924 ( .A(n_222), .Y(n_924) );
INVx1_ASAP7_75t_L g318 ( .A(n_223), .Y(n_318) );
INVx2_ASAP7_75t_L g336 ( .A(n_223), .Y(n_336) );
INVx1_ASAP7_75t_L g851 ( .A(n_224), .Y(n_851) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_226), .B(n_510), .Y(n_1186) );
OAI221xp5_ASAP7_75t_L g853 ( .A1(n_227), .A2(n_854), .B1(n_856), .B2(n_862), .C(n_866), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g978 ( .A(n_228), .Y(n_978) );
INVx1_ASAP7_75t_L g1177 ( .A(n_229), .Y(n_1177) );
AOI22xp5_ASAP7_75t_L g1456 ( .A1(n_230), .A2(n_267), .B1(n_1427), .B2(n_1430), .Y(n_1456) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_232), .A2(n_1135), .B1(n_1182), .B2(n_1183), .Y(n_1134) );
INVx1_ASAP7_75t_L g1183 ( .A(n_232), .Y(n_1183) );
INVx1_ASAP7_75t_L g1669 ( .A(n_233), .Y(n_1669) );
INVx1_ASAP7_75t_L g1067 ( .A(n_234), .Y(n_1067) );
INVx1_ASAP7_75t_L g1009 ( .A(n_235), .Y(n_1009) );
INVx1_ASAP7_75t_L g1163 ( .A(n_236), .Y(n_1163) );
CKINVDCx5p33_ASAP7_75t_R g1106 ( .A(n_237), .Y(n_1106) );
INVx1_ASAP7_75t_L g1046 ( .A(n_238), .Y(n_1046) );
INVx1_ASAP7_75t_L g1331 ( .A(n_239), .Y(n_1331) );
INVx1_ASAP7_75t_L g1381 ( .A(n_240), .Y(n_1381) );
INVx1_ASAP7_75t_L g1038 ( .A(n_241), .Y(n_1038) );
INVx1_ASAP7_75t_L g1334 ( .A(n_242), .Y(n_1334) );
INVx1_ASAP7_75t_L g813 ( .A(n_243), .Y(n_813) );
INVxp67_ASAP7_75t_L g751 ( .A(n_244), .Y(n_751) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_245), .Y(n_782) );
INVx1_ASAP7_75t_L g1374 ( .A(n_246), .Y(n_1374) );
CKINVDCx5p33_ASAP7_75t_R g1112 ( .A(n_248), .Y(n_1112) );
XOR2xp5_ASAP7_75t_L g1341 ( .A(n_249), .B(n_1342), .Y(n_1341) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_250), .A2(n_257), .B1(n_784), .B2(n_785), .Y(n_783) );
OAI221xp5_ASAP7_75t_L g804 ( .A1(n_250), .A2(n_257), .B1(n_369), .B2(n_805), .C(n_806), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_251), .Y(n_403) );
INVx1_ASAP7_75t_L g1447 ( .A(n_252), .Y(n_1447) );
OA332x1_ASAP7_75t_L g1286 ( .A1(n_253), .A2(n_376), .A3(n_1287), .B1(n_1293), .B2(n_1296), .B3(n_1299), .C1(n_1304), .C2(n_1305), .Y(n_1286) );
AOI21xp5_ASAP7_75t_L g1320 ( .A1(n_253), .A2(n_957), .B(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1161 ( .A(n_254), .Y(n_1161) );
INVx1_ASAP7_75t_L g1409 ( .A(n_255), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_255), .B(n_1419), .Y(n_1422) );
INVx1_ASAP7_75t_L g566 ( .A(n_256), .Y(n_566) );
INVx1_ASAP7_75t_L g1149 ( .A(n_258), .Y(n_1149) );
INVx1_ASAP7_75t_L g798 ( .A(n_259), .Y(n_798) );
INVx1_ASAP7_75t_L g537 ( .A(n_261), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g1001 ( .A1(n_264), .A2(n_273), .B1(n_1002), .B2(n_1003), .C(n_1004), .Y(n_1001) );
INVx1_ASAP7_75t_L g1369 ( .A(n_265), .Y(n_1369) );
CKINVDCx5p33_ASAP7_75t_R g1103 ( .A(n_266), .Y(n_1103) );
INVx1_ASAP7_75t_L g1124 ( .A(n_268), .Y(n_1124) );
INVx1_ASAP7_75t_L g820 ( .A(n_269), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g1666 ( .A(n_270), .Y(n_1666) );
INVx2_ASAP7_75t_L g315 ( .A(n_271), .Y(n_315) );
INVx1_ASAP7_75t_L g1193 ( .A(n_272), .Y(n_1193) );
INVxp67_ASAP7_75t_SL g709 ( .A(n_274), .Y(n_709) );
INVx1_ASAP7_75t_L g1206 ( .A(n_275), .Y(n_1206) );
INVxp33_ASAP7_75t_SL g351 ( .A(n_276), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_276), .A2(n_280), .B1(n_446), .B2(n_449), .C(n_455), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g1295 ( .A(n_277), .Y(n_1295) );
INVx1_ASAP7_75t_L g852 ( .A(n_278), .Y(n_852) );
INVx1_ASAP7_75t_L g799 ( .A(n_279), .Y(n_799) );
INVxp67_ASAP7_75t_L g541 ( .A(n_281), .Y(n_541) );
INVx1_ASAP7_75t_L g991 ( .A(n_282), .Y(n_991) );
OAI211xp5_ASAP7_75t_L g996 ( .A1(n_282), .A2(n_836), .B(n_997), .C(n_1005), .Y(n_996) );
INVx1_ASAP7_75t_L g1044 ( .A(n_283), .Y(n_1044) );
INVx1_ASAP7_75t_L g1113 ( .A(n_284), .Y(n_1113) );
AOI21xp33_ASAP7_75t_L g865 ( .A1(n_285), .A2(n_377), .B(n_844), .Y(n_865) );
INVx1_ASAP7_75t_L g568 ( .A(n_286), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_287), .Y(n_767) );
INVx1_ASAP7_75t_L g1125 ( .A(n_288), .Y(n_1125) );
OAI211xp5_ASAP7_75t_SL g1200 ( .A1(n_289), .A2(n_1201), .B(n_1202), .C(n_1205), .Y(n_1200) );
BUFx3_ASAP7_75t_L g424 ( .A(n_290), .Y(n_424) );
INVx1_ASAP7_75t_L g454 ( .A(n_290), .Y(n_454) );
INVx1_ASAP7_75t_L g423 ( .A(n_291), .Y(n_423) );
BUFx3_ASAP7_75t_L g439 ( .A(n_291), .Y(n_439) );
INVx1_ASAP7_75t_L g1139 ( .A(n_292), .Y(n_1139) );
INVx1_ASAP7_75t_L g939 ( .A(n_295), .Y(n_939) );
INVxp33_ASAP7_75t_L g1047 ( .A(n_296), .Y(n_1047) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_319), .B(n_1394), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_306), .Y(n_300) );
AND2x4_ASAP7_75t_L g1689 ( .A(n_301), .B(n_307), .Y(n_1689) );
NOR2xp33_ASAP7_75t_SL g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_SL g1694 ( .A(n_302), .Y(n_1694) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_302), .B(n_304), .Y(n_1702) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_304), .B(n_1694), .Y(n_1693) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_312), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g721 ( .A(n_310), .B(n_318), .Y(n_721) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g377 ( .A(n_311), .B(n_378), .Y(n_377) );
OR2x6_ASAP7_75t_L g312 ( .A(n_313), .B(n_317), .Y(n_312) );
INVx1_ASAP7_75t_L g383 ( .A(n_313), .Y(n_383) );
OR2x2_ASAP7_75t_L g511 ( .A(n_313), .B(n_366), .Y(n_511) );
INVx2_ASAP7_75t_SL g539 ( .A(n_313), .Y(n_539) );
BUFx2_ASAP7_75t_L g811 ( .A(n_313), .Y(n_811) );
BUFx6f_ASAP7_75t_L g1132 ( .A(n_313), .Y(n_1132) );
INVx2_ASAP7_75t_SL g1171 ( .A(n_313), .Y(n_1171) );
OAI22xp33_ASAP7_75t_L g1251 ( .A1(n_313), .A2(n_387), .B1(n_1252), .B2(n_1253), .Y(n_1251) );
OAI22xp33_ASAP7_75t_L g1262 ( .A1(n_313), .A2(n_387), .B1(n_1263), .B2(n_1264), .Y(n_1262) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g330 ( .A(n_315), .Y(n_330) );
INVx1_ASAP7_75t_L g342 ( .A(n_315), .Y(n_342) );
AND2x2_ASAP7_75t_L g350 ( .A(n_315), .B(n_316), .Y(n_350) );
AND2x4_ASAP7_75t_L g357 ( .A(n_315), .B(n_343), .Y(n_357) );
INVx1_ASAP7_75t_L g390 ( .A(n_315), .Y(n_390) );
INVx1_ASAP7_75t_L g332 ( .A(n_316), .Y(n_332) );
INVx2_ASAP7_75t_L g343 ( .A(n_316), .Y(n_343) );
INVx1_ASAP7_75t_L g364 ( .A(n_316), .Y(n_364) );
INVx1_ASAP7_75t_L g389 ( .A(n_316), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_316), .B(n_330), .Y(n_397) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_1031), .B1(n_1032), .B2(n_1393), .Y(n_319) );
INVx1_ASAP7_75t_L g1393 ( .A(n_320), .Y(n_1393) );
AO22x2_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_769), .B1(n_1029), .B2(n_1030), .Y(n_320) );
INVx1_ASAP7_75t_L g1029 ( .A(n_321), .Y(n_1029) );
XNOR2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_516), .Y(n_321) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_416), .Y(n_323) );
NOR3xp33_ASAP7_75t_SL g324 ( .A(n_325), .B(n_358), .C(n_374), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_327), .A2(n_338), .B1(n_711), .B2(n_712), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_327), .A2(n_347), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_333), .Y(n_327) );
AND2x2_ASAP7_75t_L g524 ( .A(n_328), .B(n_333), .Y(n_524) );
AND2x2_ASAP7_75t_L g803 ( .A(n_328), .B(n_333), .Y(n_803) );
AND2x2_ASAP7_75t_L g917 ( .A(n_328), .B(n_333), .Y(n_917) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g654 ( .A(n_329), .B(n_335), .Y(n_654) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_329), .Y(n_672) );
BUFx6f_ASAP7_75t_L g728 ( .A(n_329), .Y(n_728) );
INVx1_ASAP7_75t_L g840 ( .A(n_329), .Y(n_840) );
INVx1_ASAP7_75t_L g1220 ( .A(n_329), .Y(n_1220) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g372 ( .A(n_330), .Y(n_372) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x6_ASAP7_75t_L g339 ( .A(n_333), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g347 ( .A(n_333), .B(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g354 ( .A(n_333), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g555 ( .A(n_333), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_333), .B(n_546), .Y(n_1162) );
AOI22xp5_ASAP7_75t_L g1256 ( .A1(n_333), .A2(n_1227), .B1(n_1257), .B2(n_1261), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_333), .B(n_661), .Y(n_1306) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g412 ( .A(n_334), .Y(n_412) );
OR2x2_ASAP7_75t_L g694 ( .A(n_334), .B(n_426), .Y(n_694) );
INVx2_ASAP7_75t_L g650 ( .A(n_335), .Y(n_650) );
AND2x4_ASAP7_75t_L g855 ( .A(n_335), .B(n_677), .Y(n_855) );
INVx1_ASAP7_75t_L g378 ( .A(n_336), .Y(n_378) );
INVx1_ASAP7_75t_L g414 ( .A(n_336), .Y(n_414) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_339), .A2(n_354), .B1(n_798), .B2(n_799), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_339), .A2(n_353), .B1(n_912), .B2(n_913), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_339), .A2(n_716), .B1(n_1043), .B2(n_1044), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_339), .A2(n_1103), .B1(n_1117), .B2(n_1118), .Y(n_1116) );
NAND2x1p5_ASAP7_75t_L g373 ( .A(n_340), .B(n_365), .Y(n_373) );
BUFx2_ASAP7_75t_L g1002 ( .A(n_340), .Y(n_1002) );
BUFx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_341), .Y(n_556) );
BUFx2_ASAP7_75t_L g608 ( .A(n_341), .Y(n_608) );
BUFx3_ASAP7_75t_L g679 ( .A(n_341), .Y(n_679) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_341), .Y(n_848) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B1(n_351), .B2(n_352), .Y(n_344) );
OAI221xp5_ASAP7_75t_L g455 ( .A1(n_345), .A2(n_456), .B1(n_461), .B2(n_462), .C(n_465), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_346), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_713) );
BUFx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g601 ( .A(n_347), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_347), .A2(n_801), .B1(n_802), .B2(n_803), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_347), .A2(n_915), .B1(n_916), .B2(n_917), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_347), .A2(n_803), .B1(n_1104), .B2(n_1120), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_347), .A2(n_524), .B1(n_1165), .B2(n_1166), .Y(n_1164) );
AOI221xp5_ASAP7_75t_L g1229 ( .A1(n_347), .A2(n_917), .B1(n_1230), .B2(n_1231), .C(n_1232), .Y(n_1229) );
INVx1_ASAP7_75t_L g845 ( .A(n_348), .Y(n_845) );
BUFx2_ASAP7_75t_L g1217 ( .A(n_348), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_348), .A2(n_608), .B1(n_1259), .B2(n_1260), .Y(n_1258) );
INVx2_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_SL g661 ( .A(n_349), .Y(n_661) );
INVx2_ASAP7_75t_L g690 ( .A(n_349), .Y(n_690) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_350), .Y(n_677) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g603 ( .A(n_354), .Y(n_603) );
BUFx2_ASAP7_75t_L g716 ( .A(n_354), .Y(n_716) );
BUFx2_ASAP7_75t_L g1118 ( .A(n_354), .Y(n_1118) );
BUFx3_ASAP7_75t_L g400 ( .A(n_355), .Y(n_400) );
INVx2_ASAP7_75t_L g860 ( .A(n_355), .Y(n_860) );
INVx1_ASAP7_75t_L g1662 ( .A(n_355), .Y(n_1662) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx3_ASAP7_75t_L g546 ( .A(n_356), .Y(n_546) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_356), .Y(n_674) );
INVx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_357), .Y(n_532) );
INVx1_ASAP7_75t_L g652 ( .A(n_357), .Y(n_652) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_SL g919 ( .A(n_360), .Y(n_919) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_361), .Y(n_805) );
NAND2x1_ASAP7_75t_SL g361 ( .A(n_362), .B(n_365), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g685 ( .A(n_362), .B(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_362), .A2(n_371), .B1(n_1358), .B2(n_1360), .Y(n_1383) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_364), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_365), .B(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g605 ( .A(n_365), .B(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g607 ( .A(n_365), .B(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g706 ( .A(n_365), .B(n_707), .Y(n_706) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g669 ( .A(n_367), .Y(n_669) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx4f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx4f_ASAP7_75t_L g525 ( .A(n_370), .Y(n_525) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x6_ASAP7_75t_L g687 ( .A(n_372), .B(n_668), .Y(n_687) );
BUFx3_ASAP7_75t_L g806 ( .A(n_373), .Y(n_806) );
BUFx2_ASAP7_75t_L g1049 ( .A(n_373), .Y(n_1049) );
OAI33xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_380), .A3(n_391), .B1(n_401), .B2(n_404), .B3(n_409), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI33xp33_ASAP7_75t_L g807 ( .A1(n_376), .A2(n_409), .A3(n_808), .B1(n_814), .B2(n_821), .B3(n_825), .Y(n_807) );
INVx1_ASAP7_75t_L g922 ( .A(n_376), .Y(n_922) );
OAI33xp33_ASAP7_75t_L g1050 ( .A1(n_376), .A2(n_409), .A3(n_1051), .B1(n_1057), .B2(n_1062), .B3(n_1068), .Y(n_1050) );
OAI33xp33_ASAP7_75t_L g1122 ( .A1(n_376), .A2(n_409), .A3(n_1123), .B1(n_1126), .B2(n_1129), .B3(n_1131), .Y(n_1122) );
OAI33xp33_ASAP7_75t_L g1168 ( .A1(n_376), .A2(n_552), .A3(n_1169), .B1(n_1174), .B2(n_1178), .B3(n_1181), .Y(n_1168) );
OR2x6_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
BUFx2_ASAP7_75t_L g505 ( .A(n_379), .Y(n_505) );
INVx2_ASAP7_75t_L g616 ( .A(n_379), .Y(n_616) );
OAI22xp5_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_382), .B1(n_384), .B2(n_385), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_382), .A2(n_393), .B1(n_402), .B2(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g550 ( .A(n_383), .Y(n_550) );
OAI22xp5_ASAP7_75t_SL g548 ( .A1(n_385), .A2(n_549), .B1(n_550), .B2(n_551), .Y(n_548) );
OAI22xp33_ASAP7_75t_L g1068 ( .A1(n_385), .A2(n_1053), .B1(n_1069), .B2(n_1070), .Y(n_1068) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g1013 ( .A(n_386), .Y(n_1013) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g407 ( .A(n_387), .Y(n_407) );
BUFx3_ASAP7_75t_L g926 ( .A(n_387), .Y(n_926) );
OAI22xp33_ASAP7_75t_L g1296 ( .A1(n_387), .A2(n_1132), .B1(n_1297), .B2(n_1298), .Y(n_1296) );
OAI221xp5_ASAP7_75t_L g1375 ( .A1(n_387), .A2(n_550), .B1(n_1376), .B2(n_1377), .C(n_1378), .Y(n_1375) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
AND2x2_ASAP7_75t_L g536 ( .A(n_389), .B(n_390), .Y(n_536) );
INVx1_ASAP7_75t_L g708 ( .A(n_390), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_398), .B2(n_399), .Y(n_391) );
BUFx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g1372 ( .A1(n_394), .A2(n_1060), .B1(n_1373), .B2(n_1374), .Y(n_1372) );
INVx2_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g529 ( .A(n_395), .Y(n_529) );
INVx2_ASAP7_75t_L g1175 ( .A(n_395), .Y(n_1175) );
BUFx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g663 ( .A(n_396), .Y(n_663) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx2_ASAP7_75t_L g544 ( .A(n_397), .Y(n_544) );
INVx1_ASAP7_75t_L g817 ( .A(n_397), .Y(n_817) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_399), .A2(n_405), .B1(n_406), .B2(n_408), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_399), .A2(n_935), .B1(n_936), .B2(n_939), .Y(n_934) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_400), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_402), .A2(n_405), .B1(n_498), .B2(n_500), .Y(n_497) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_403), .A2(n_419), .B(n_428), .C(n_445), .Y(n_418) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g808 ( .A1(n_407), .A2(n_809), .B1(n_812), .B2(n_813), .Y(n_808) );
OAI22xp33_ASAP7_75t_L g1123 ( .A1(n_407), .A2(n_1053), .B1(n_1124), .B2(n_1125), .Y(n_1123) );
OAI22xp33_ASAP7_75t_L g1293 ( .A1(n_407), .A2(n_538), .B1(n_1294), .B2(n_1295), .Y(n_1293) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_408), .A2(n_468), .B1(n_474), .B2(n_483), .C(n_491), .Y(n_467) );
INVx1_ASAP7_75t_L g732 ( .A(n_409), .Y(n_732) );
OAI33xp33_ASAP7_75t_L g920 ( .A1(n_409), .A2(n_921), .A3(n_923), .B1(n_927), .B2(n_934), .B3(n_940), .Y(n_920) );
CKINVDCx8_ASAP7_75t_R g409 ( .A(n_410), .Y(n_409) );
INVx5_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx6_ASAP7_75t_L g553 ( .A(n_411), .Y(n_553) );
OR2x6_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_412), .B(n_431), .Y(n_636) );
INVx2_ASAP7_75t_L g681 ( .A(n_413), .Y(n_681) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_502), .B1(n_506), .B2(n_507), .Y(n_416) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_467), .C(n_497), .Y(n_417) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI211xp5_ASAP7_75t_L g737 ( .A1(n_420), .A2(n_738), .B(n_739), .C(n_740), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_420), .A2(n_498), .B1(n_935), .B2(n_941), .Y(n_965) );
AOI211xp5_ASAP7_75t_SL g1074 ( .A1(n_420), .A2(n_1064), .B(n_1075), .C(n_1076), .Y(n_1074) );
AOI211xp5_ASAP7_75t_SL g1096 ( .A1(n_420), .A2(n_1097), .B(n_1098), .C(n_1100), .Y(n_1096) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_425), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx3_ASAP7_75t_L g448 ( .A(n_422), .Y(n_448) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_422), .Y(n_572) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_422), .Y(n_580) );
INVx2_ASAP7_75t_SL g620 ( .A(n_422), .Y(n_620) );
BUFx2_ASAP7_75t_L g753 ( .A(n_422), .Y(n_753) );
BUFx6f_ASAP7_75t_L g951 ( .A(n_422), .Y(n_951) );
BUFx2_ASAP7_75t_L g960 ( .A(n_422), .Y(n_960) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_422), .Y(n_1101) );
HB1xp67_ASAP7_75t_L g1152 ( .A(n_422), .Y(n_1152) );
AND2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g460 ( .A(n_423), .Y(n_460) );
INVx2_ASAP7_75t_L g444 ( .A(n_424), .Y(n_444) );
AND2x2_ASAP7_75t_L g473 ( .A(n_424), .B(n_439), .Y(n_473) );
AND2x4_ASAP7_75t_L g471 ( .A(n_425), .B(n_472), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_425), .A2(n_471), .B1(n_551), .B2(n_570), .C(n_576), .Y(n_569) );
AND2x2_ASAP7_75t_L g781 ( .A(n_425), .B(n_572), .Y(n_781) );
AOI222xp33_ASAP7_75t_L g1266 ( .A1(n_425), .A2(n_565), .B1(n_567), .B2(n_1247), .C1(n_1248), .C2(n_1267), .Y(n_1266) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g499 ( .A(n_426), .B(n_464), .Y(n_499) );
OR2x2_ASAP7_75t_L g501 ( .A(n_426), .B(n_452), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g1312 ( .A1(n_426), .A2(n_1313), .B(n_1314), .C(n_1315), .Y(n_1312) );
INVx1_ASAP7_75t_L g432 ( .A(n_427), .Y(n_432) );
INVx2_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g947 ( .A(n_430), .Y(n_947) );
INVx2_ASAP7_75t_SL g1329 ( .A(n_430), .Y(n_1329) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_435), .Y(n_430) );
AND2x2_ASAP7_75t_L g441 ( .A(n_431), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g495 ( .A(n_431), .Y(n_495) );
AND2x2_ASAP7_75t_L g515 ( .A(n_431), .B(n_487), .Y(n_515) );
AND2x4_ASAP7_75t_L g565 ( .A(n_431), .B(n_435), .Y(n_565) );
AND2x4_ASAP7_75t_L g567 ( .A(n_431), .B(n_442), .Y(n_567) );
BUFx2_ASAP7_75t_L g577 ( .A(n_431), .Y(n_577) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
AND2x4_ASAP7_75t_L g465 ( .A(n_433), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g482 ( .A(n_434), .B(n_466), .Y(n_482) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g634 ( .A(n_436), .Y(n_634) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g487 ( .A(n_438), .B(n_444), .Y(n_487) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g453 ( .A(n_439), .B(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g640 ( .A(n_442), .Y(n_640) );
BUFx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g589 ( .A(n_450), .Y(n_589) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g985 ( .A(n_451), .Y(n_985) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_453), .Y(n_490) );
INVx1_ASAP7_75t_L g629 ( .A(n_453), .Y(n_629) );
INVx1_ASAP7_75t_L g742 ( .A(n_453), .Y(n_742) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_453), .Y(n_780) );
INVx1_ASAP7_75t_L g459 ( .A(n_454), .Y(n_459) );
INVx2_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g699 ( .A(n_458), .Y(n_699) );
INVx1_ASAP7_75t_L g746 ( .A(n_458), .Y(n_746) );
INVx1_ASAP7_75t_L g954 ( .A(n_458), .Y(n_954) );
INVx1_ASAP7_75t_L g981 ( .A(n_458), .Y(n_981) );
BUFx4f_ASAP7_75t_L g1197 ( .A(n_458), .Y(n_1197) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
OR2x2_ASAP7_75t_L g464 ( .A(n_459), .B(n_460), .Y(n_464) );
OAI221xp5_ASAP7_75t_L g977 ( .A1(n_462), .A2(n_978), .B1(n_979), .B2(n_982), .C(n_983), .Y(n_977) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g693 ( .A(n_463), .Y(n_693) );
INVx2_ASAP7_75t_L g955 ( .A(n_463), .Y(n_955) );
INVx2_ASAP7_75t_L g1190 ( .A(n_463), .Y(n_1190) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g574 ( .A(n_464), .Y(n_574) );
BUFx2_ASAP7_75t_L g747 ( .A(n_464), .Y(n_747) );
INVx1_ASAP7_75t_L g1677 ( .A(n_464), .Y(n_1677) );
INVx1_ASAP7_75t_L g596 ( .A(n_465), .Y(n_596) );
AND2x4_ASAP7_75t_L g630 ( .A(n_465), .B(n_514), .Y(n_630) );
AND2x4_ASAP7_75t_L g892 ( .A(n_465), .B(n_514), .Y(n_892) );
INVx2_ASAP7_75t_SL g957 ( .A(n_465), .Y(n_957) );
OAI221xp5_ASAP7_75t_L g1078 ( .A1(n_465), .A2(n_693), .B1(n_746), .B2(n_1044), .C(n_1046), .Y(n_1078) );
OAI221xp5_ASAP7_75t_L g1102 ( .A1(n_465), .A2(n_693), .B1(n_746), .B2(n_1103), .C(n_1104), .Y(n_1102) );
CKINVDCx5p33_ASAP7_75t_R g1276 ( .A(n_465), .Y(n_1276) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g958 ( .A1(n_470), .A2(n_493), .B1(n_942), .B2(n_959), .C(n_963), .Y(n_958) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_471), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g786 ( .A1(n_471), .A2(n_576), .B1(n_787), .B2(n_788), .C(n_789), .Y(n_786) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_471), .Y(n_1080) );
AOI221xp5_ASAP7_75t_L g1105 ( .A1(n_471), .A2(n_576), .B1(n_1106), .B2(n_1107), .C(n_1109), .Y(n_1105) );
INVx2_ASAP7_75t_SL g1143 ( .A(n_471), .Y(n_1143) );
AND2x4_ASAP7_75t_L g576 ( .A(n_472), .B(n_577), .Y(n_576) );
BUFx4f_ASAP7_75t_L g581 ( .A(n_472), .Y(n_581) );
INVx1_ASAP7_75t_L g593 ( .A(n_472), .Y(n_593) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_472), .Y(n_623) );
INVx2_ASAP7_75t_SL g1083 ( .A(n_472), .Y(n_1083) );
AOI22xp5_ASAP7_75t_L g1268 ( .A1(n_472), .A2(n_572), .B1(n_1264), .B2(n_1269), .Y(n_1268) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_473), .Y(n_479) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g756 ( .A(n_478), .Y(n_756) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_479), .Y(n_496) );
INVx1_ASAP7_75t_L g644 ( .A(n_479), .Y(n_644) );
BUFx6f_ASAP7_75t_L g1275 ( .A(n_479), .Y(n_1275) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
BUFx3_ASAP7_75t_L g583 ( .A(n_482), .Y(n_583) );
INVx1_ASAP7_75t_L g617 ( .A(n_482), .Y(n_617) );
INVx2_ASAP7_75t_L g759 ( .A(n_482), .Y(n_759) );
INVx1_ASAP7_75t_L g1327 ( .A(n_482), .Y(n_1327) );
BUFx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g903 ( .A(n_485), .B(n_901), .Y(n_903) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g1321 ( .A(n_486), .Y(n_1321) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx6_ASAP7_75t_L g595 ( .A(n_487), .Y(n_595) );
BUFx2_ASAP7_75t_L g762 ( .A(n_487), .Y(n_762) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI221xp5_ASAP7_75t_SL g578 ( .A1(n_489), .A2(n_530), .B1(n_537), .B2(n_573), .C(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g891 ( .A(n_489), .Y(n_891) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g575 ( .A(n_490), .Y(n_575) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_490), .Y(n_621) );
INVx1_ASAP7_75t_L g881 ( .A(n_490), .Y(n_881) );
HB1xp67_ASAP7_75t_L g1147 ( .A(n_490), .Y(n_1147) );
BUFx6f_ASAP7_75t_L g1278 ( .A(n_490), .Y(n_1278) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g749 ( .A1(n_493), .A2(n_750), .B1(n_751), .B2(n_752), .C(n_760), .Y(n_749) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g877 ( .A(n_496), .Y(n_877) );
BUFx6f_ASAP7_75t_L g961 ( .A(n_496), .Y(n_961) );
INVx1_ASAP7_75t_L g1351 ( .A(n_496), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_498), .A2(n_500), .B1(n_765), .B2(n_766), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_498), .A2(n_500), .B1(n_791), .B2(n_792), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_498), .A2(n_500), .B1(n_1067), .B2(n_1069), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_498), .A2(n_500), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
AOI22xp5_ASAP7_75t_L g1138 ( .A1(n_498), .A2(n_500), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
INVx6_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AOI211xp5_ASAP7_75t_L g945 ( .A1(n_500), .A2(n_939), .B(n_946), .C(n_948), .Y(n_945) );
INVx4_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_SL g1024 ( .A(n_502), .Y(n_1024) );
INVx5_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g1650 ( .A1(n_503), .A2(n_1651), .B(n_1659), .Y(n_1650) );
BUFx8_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
AOI31xp33_ASAP7_75t_L g736 ( .A1(n_504), .A2(n_737), .A3(n_749), .B(n_764), .Y(n_736) );
INVx2_ASAP7_75t_L g1072 ( .A(n_504), .Y(n_1072) );
OAI31xp33_ASAP7_75t_L g1361 ( .A1(n_504), .A2(n_1362), .A3(n_1364), .B(n_1384), .Y(n_1361) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g599 ( .A(n_505), .Y(n_599) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g943 ( .A1(n_509), .A2(n_599), .B1(n_944), .B2(n_966), .Y(n_943) );
INVx5_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g734 ( .A(n_510), .Y(n_734) );
INVx2_ASAP7_75t_SL g794 ( .A(n_510), .Y(n_794) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g1255 ( .A(n_511), .Y(n_1255) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x6_ASAP7_75t_L g870 ( .A(n_513), .B(n_871), .Y(n_870) );
AOI222xp33_ASAP7_75t_L g1386 ( .A1(n_513), .A2(n_903), .B1(n_1374), .B2(n_1377), .C1(n_1381), .C2(n_1387), .Y(n_1386) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g561 ( .A(n_515), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_515), .B(n_1331), .Y(n_1330) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B1(n_701), .B2(n_768), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AO22x2_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_609), .B1(n_610), .B2(n_700), .Y(n_518) );
INVx1_ASAP7_75t_L g700 ( .A(n_519), .Y(n_700) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_557), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_526), .Y(n_521) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g1309 ( .A(n_524), .Y(n_1309) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B1(n_530), .B2(n_531), .Y(n_527) );
OAI221xp5_ASAP7_75t_L g997 ( .A1(n_531), .A2(n_998), .B1(n_999), .B2(n_1000), .C(n_1001), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_531), .A2(n_1097), .B1(n_1112), .B2(n_1130), .Y(n_1129) );
INVx4_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_SL g1303 ( .A(n_532), .Y(n_1303) );
OAI22xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_537), .B2(n_538), .Y(n_533) );
OR2x6_ASAP7_75t_L g667 ( .A(n_535), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g827 ( .A(n_535), .Y(n_827) );
OR2x2_ASAP7_75t_L g866 ( .A(n_535), .B(n_668), .Y(n_866) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx3_ASAP7_75t_L g658 ( .A(n_536), .Y(n_658) );
INVx2_ASAP7_75t_L g863 ( .A(n_536), .Y(n_863) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_536), .Y(n_1056) );
OAI22xp33_ASAP7_75t_L g923 ( .A1(n_538), .A2(n_924), .B1(n_925), .B2(n_926), .Y(n_923) );
OAI22xp33_ASAP7_75t_L g940 ( .A1(n_538), .A2(n_926), .B1(n_941), .B2(n_942), .Y(n_940) );
OAI221xp5_ASAP7_75t_L g1012 ( .A1(n_538), .A2(n_978), .B1(n_982), .B2(n_1013), .C(n_1014), .Y(n_1012) );
OAI221xp5_ASAP7_75t_L g1664 ( .A1(n_538), .A2(n_658), .B1(n_1665), .B2(n_1666), .C(n_1667), .Y(n_1664) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_545), .B2(n_547), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_542), .A2(n_1017), .B1(n_1018), .B2(n_1020), .Y(n_1016) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g1289 ( .A(n_544), .Y(n_1289) );
INVx1_ASAP7_75t_L g1019 ( .A(n_545), .Y(n_1019) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g819 ( .A(n_546), .Y(n_819) );
INVx2_ASAP7_75t_L g824 ( .A(n_546), .Y(n_824) );
INVx2_ASAP7_75t_L g842 ( .A(n_546), .Y(n_842) );
HB1xp67_ASAP7_75t_L g1292 ( .A(n_546), .Y(n_1292) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g1304 ( .A(n_553), .Y(n_1304) );
INVxp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_555), .A2(n_1161), .B1(n_1162), .B2(n_1163), .Y(n_1160) );
INVx1_ASAP7_75t_L g1234 ( .A(n_555), .Y(n_1234) );
AOI21xp5_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_597), .B(n_600), .Y(n_557) );
NAND4xp25_ASAP7_75t_SL g558 ( .A(n_559), .B(n_569), .C(n_578), .D(n_584), .Y(n_558) );
AOI222xp33_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_562), .B1(n_563), .B2(n_566), .C1(n_567), .C2(n_568), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g1273 ( .A1(n_560), .A2(n_1254), .B1(n_1274), .B2(n_1277), .Y(n_1273) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx4_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g784 ( .A(n_565), .Y(n_784) );
INVx1_ASAP7_75t_SL g1155 ( .A(n_565), .Y(n_1155) );
AOI22xp5_ASAP7_75t_L g1202 ( .A1(n_565), .A2(n_567), .B1(n_1203), .B2(n_1204), .Y(n_1202) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_566), .A2(n_605), .B(n_607), .Y(n_604) );
INVx2_ASAP7_75t_SL g785 ( .A(n_567), .Y(n_785) );
INVx2_ASAP7_75t_L g1099 ( .A(n_567), .Y(n_1099) );
OR2x2_ASAP7_75t_L g695 ( .A(n_571), .B(n_694), .Y(n_695) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx4f_ASAP7_75t_L g889 ( .A(n_572), .Y(n_889) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g1355 ( .A(n_575), .Y(n_1355) );
AOI221xp5_ASAP7_75t_L g1079 ( .A1(n_576), .A2(n_1070), .B1(n_1080), .B2(n_1081), .C(n_1085), .Y(n_1079) );
AOI221xp5_ASAP7_75t_L g1141 ( .A1(n_576), .A2(n_1142), .B1(n_1144), .B2(n_1145), .C(n_1146), .Y(n_1141) );
INVx1_ASAP7_75t_L g1199 ( .A(n_576), .Y(n_1199) );
AOI21xp5_ASAP7_75t_L g1270 ( .A1(n_576), .A2(n_1271), .B(n_1272), .Y(n_1270) );
INVx1_ASAP7_75t_L g1315 ( .A(n_576), .Y(n_1315) );
BUFx3_ASAP7_75t_L g586 ( .A(n_580), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_581), .A2(n_900), .B1(n_1298), .B2(n_1300), .Y(n_1314) );
INVx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g962 ( .A(n_583), .Y(n_962) );
INVxp67_ASAP7_75t_L g1084 ( .A(n_583), .Y(n_1084) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_587), .B1(n_588), .B2(n_590), .C(n_591), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_595), .Y(n_626) );
INVx2_ASAP7_75t_L g879 ( .A(n_595), .Y(n_879) );
INVx2_ASAP7_75t_L g1087 ( .A(n_595), .Y(n_1087) );
INVx1_ASAP7_75t_L g1325 ( .A(n_595), .Y(n_1325) );
INVx1_ASAP7_75t_L g748 ( .A(n_596), .Y(n_748) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI21x1_ASAP7_75t_L g646 ( .A1(n_599), .A2(n_647), .B(n_670), .Y(n_646) );
OAI31xp33_ASAP7_75t_L g1311 ( .A1(n_599), .A2(n_1312), .A3(n_1316), .B(n_1328), .Y(n_1311) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_605), .A2(n_607), .B1(n_705), .B2(n_706), .C(n_709), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g1228 ( .A1(n_605), .A2(n_607), .B1(n_706), .B2(n_1203), .C(n_1204), .Y(n_1228) );
AOI221xp5_ASAP7_75t_L g1246 ( .A1(n_605), .A2(n_607), .B1(n_706), .B2(n_1247), .C(n_1248), .Y(n_1246) );
AOI221xp5_ASAP7_75t_L g1332 ( .A1(n_605), .A2(n_607), .B1(n_706), .B2(n_1333), .C(n_1334), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_606), .B(n_873), .Y(n_1008) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_608), .Y(n_729) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR4xp75_ASAP7_75t_L g611 ( .A(n_612), .B(n_646), .C(n_691), .D(n_696), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_631), .Y(n_612) );
AOI33xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_618), .A3(n_622), .B1(n_624), .B2(n_627), .B3(n_630), .Y(n_613) );
INVx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_SL g1672 ( .A1(n_615), .A2(n_986), .B1(n_1673), .B2(n_1675), .Y(n_1672) );
OR2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x4_ASAP7_75t_L g720 ( .A(n_616), .B(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g774 ( .A(n_616), .Y(n_774) );
BUFx2_ASAP7_75t_L g867 ( .A(n_616), .Y(n_867) );
OR2x6_ASAP7_75t_L g883 ( .A(n_616), .B(n_759), .Y(n_883) );
AND2x4_ASAP7_75t_L g1215 ( .A(n_616), .B(n_721), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_616), .B(n_681), .Y(n_1227) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_620), .A2(n_859), .B1(n_861), .B2(n_881), .Y(n_880) );
INVx2_ASAP7_75t_L g900 ( .A(n_620), .Y(n_900) );
INVx1_ASAP7_75t_L g1077 ( .A(n_620), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_621), .A2(n_879), .B1(n_1297), .B2(n_1302), .Y(n_1313) );
INVx1_ASAP7_75t_L g886 ( .A(n_623), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_623), .B(n_645), .Y(n_897) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx4_ASAP7_75t_L g964 ( .A(n_626), .Y(n_964) );
BUFx2_ASAP7_75t_L g1348 ( .A(n_628), .Y(n_1348) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g697 ( .A(n_629), .B(n_694), .Y(n_697) );
OR2x6_ASAP7_75t_L g1027 ( .A(n_629), .B(n_694), .Y(n_1027) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_637), .B1(n_638), .B2(n_641), .C(n_642), .Y(n_631) );
INVx2_ASAP7_75t_L g994 ( .A(n_632), .Y(n_994) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g895 ( .A(n_633), .Y(n_895) );
INVx1_ASAP7_75t_L g1359 ( .A(n_633), .Y(n_1359) );
NAND2x1p5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx2_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
OR2x6_ASAP7_75t_L g639 ( .A(n_636), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g645 ( .A(n_636), .Y(n_645) );
OR2x2_ASAP7_75t_L g896 ( .A(n_636), .B(n_640), .Y(n_896) );
AOI221xp5_ASAP7_75t_L g1357 ( .A1(n_638), .A2(n_642), .B1(n_1358), .B2(n_1359), .C(n_1360), .Y(n_1357) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx2_ASAP7_75t_L g974 ( .A(n_642), .Y(n_974) );
NOR3xp33_ASAP7_75t_L g1670 ( .A(n_642), .B(n_1671), .C(n_1672), .Y(n_1670) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI221x1_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_653), .B1(n_654), .B2(n_655), .C(n_656), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_648), .A2(n_654), .B1(n_851), .B2(n_852), .Y(n_850) );
INVx3_ASAP7_75t_L g1023 ( .A(n_648), .Y(n_1023) );
INVx3_ASAP7_75t_L g1363 ( .A(n_648), .Y(n_1363) );
AOI22xp33_ASAP7_75t_L g1652 ( .A1(n_648), .A2(n_654), .B1(n_1653), .B2(n_1654), .Y(n_1652) );
AND2x4_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
AND2x4_ASAP7_75t_L g682 ( .A(n_649), .B(n_679), .Y(n_682) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g665 ( .A(n_651), .Y(n_665) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g1180 ( .A(n_652), .Y(n_1180) );
INVx3_ASAP7_75t_L g1022 ( .A(n_654), .Y(n_1022) );
INVx3_ASAP7_75t_L g1385 ( .A(n_654), .Y(n_1385) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_662), .B(n_667), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_659), .B(n_660), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g1382 ( .A1(n_658), .A2(n_668), .B(n_1383), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_661), .B(n_873), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_662) );
INVx2_ASAP7_75t_L g930 ( .A(n_663), .Y(n_930) );
INVx1_ASAP7_75t_L g1223 ( .A(n_665), .Y(n_1223) );
INVx1_ASAP7_75t_L g686 ( .A(n_668), .Y(n_686) );
INVx1_ASAP7_75t_L g873 ( .A(n_668), .Y(n_873) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI221xp5_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_675), .B1(n_682), .B2(n_683), .C(n_684), .Y(n_670) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g933 ( .A(n_674), .Y(n_933) );
INVx2_ASAP7_75t_L g1061 ( .A(n_674), .Y(n_1061) );
BUFx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
BUFx6f_ASAP7_75t_L g1003 ( .A(n_677), .Y(n_1003) );
INVx3_ASAP7_75t_L g1226 ( .A(n_677), .Y(n_1226) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g1378 ( .A(n_680), .Y(n_1378) );
INVx2_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g1004 ( .A(n_681), .Y(n_1004) );
INVx8_ASAP7_75t_L g836 ( .A(n_682), .Y(n_836) );
CKINVDCx11_ASAP7_75t_R g1010 ( .A(n_687), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
BUFx3_ASAP7_75t_L g723 ( .A(n_690), .Y(n_723) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
OR2x6_ASAP7_75t_L g698 ( .A(n_694), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g901 ( .A(n_694), .Y(n_901) );
CKINVDCx6p67_ASAP7_75t_R g1389 ( .A(n_698), .Y(n_1389) );
INVx1_ASAP7_75t_L g990 ( .A(n_699), .Y(n_990) );
INVx2_ASAP7_75t_L g768 ( .A(n_701), .Y(n_768) );
XOR2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_767), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_733), .Y(n_702) );
AND4x1_ASAP7_75t_L g703 ( .A(n_704), .B(n_710), .C(n_713), .D(n_717), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_712), .A2(n_714), .B1(n_744), .B2(n_747), .C(n_748), .Y(n_743) );
AOI33xp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_722), .A3(n_726), .B1(n_730), .B2(n_731), .B3(n_732), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g1015 ( .A(n_721), .Y(n_1015) );
BUFx2_ASAP7_75t_SL g1667 ( .A(n_721), .Y(n_1667) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
BUFx3_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B(n_736), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g1071 ( .A1(n_734), .A2(n_1072), .B1(n_1073), .B2(n_1090), .Y(n_1071) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_734), .A2(n_774), .B1(n_1095), .B2(n_1113), .Y(n_1094) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g763 ( .A(n_742), .Y(n_763) );
INVx1_ASAP7_75t_L g952 ( .A(n_742), .Y(n_952) );
OAI211xp5_ASAP7_75t_L g1317 ( .A1(n_744), .A2(n_1318), .B(n_1319), .C(n_1320), .Y(n_1317) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI221xp5_ASAP7_75t_L g987 ( .A1(n_747), .A2(n_988), .B1(n_989), .B2(n_991), .C(n_992), .Y(n_987) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g1030 ( .A(n_769), .Y(n_1030) );
XNOR2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_830), .Y(n_769) );
INVx3_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g828 ( .A(n_772), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_795), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .B1(n_793), .B2(n_794), .Y(n_773) );
NOR2xp67_ASAP7_75t_L g871 ( .A(n_774), .B(n_872), .Y(n_871) );
INVx2_ASAP7_75t_L g1212 ( .A(n_774), .Y(n_1212) );
NAND3xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_786), .C(n_790), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B1(n_781), .B2(n_782), .C(n_783), .Y(n_776) );
BUFx6f_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g1192 ( .A(n_780), .Y(n_1192) );
AOI221xp5_ASAP7_75t_L g1148 ( .A1(n_781), .A2(n_1149), .B1(n_1150), .B2(n_1151), .C(n_1154), .Y(n_1148) );
INVx1_ASAP7_75t_L g1201 ( .A(n_781), .Y(n_1201) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_782), .A2(n_792), .B1(n_815), .B2(n_822), .Y(n_821) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_789), .A2(n_791), .B1(n_809), .B2(n_826), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g1136 ( .A1(n_794), .A2(n_1137), .B1(n_1156), .B2(n_1157), .Y(n_1136) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_804), .C(n_807), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_800), .Y(n_796) );
INVx2_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g1053 ( .A(n_810), .Y(n_1053) );
INVx1_ASAP7_75t_L g1370 ( .A(n_810), .Y(n_1370) );
INVx2_ASAP7_75t_SL g810 ( .A(n_811), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_818), .B1(n_819), .B2(n_820), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_815), .A2(n_1058), .B1(n_1059), .B2(n_1060), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_815), .A2(n_1060), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
BUFx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
BUFx2_ASAP7_75t_L g1301 ( .A(n_816), .Y(n_1301) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
HB1xp67_ASAP7_75t_L g858 ( .A(n_817), .Y(n_858) );
INVx1_ASAP7_75t_L g938 ( .A(n_817), .Y(n_938) );
INVx2_ASAP7_75t_L g998 ( .A(n_817), .Y(n_998) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g1066 ( .A(n_824), .Y(n_1066) );
INVx1_ASAP7_75t_L g1221 ( .A(n_824), .Y(n_1221) );
OAI22xp33_ASAP7_75t_L g1169 ( .A1(n_826), .A2(n_1170), .B1(n_1172), .B2(n_1173), .Y(n_1169) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
XOR2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_967), .Y(n_830) );
XNOR2xp5_ASAP7_75t_L g831 ( .A(n_832), .B(n_906), .Y(n_831) );
NAND4xp25_ASAP7_75t_L g833 ( .A(n_834), .B(n_868), .C(n_874), .D(n_898), .Y(n_833) );
OAI21xp5_ASAP7_75t_SL g834 ( .A1(n_835), .A2(n_853), .B(n_867), .Y(n_834) );
AOI21xp5_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_843), .B(n_849), .Y(n_837) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx2_ASAP7_75t_SL g847 ( .A(n_848), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_851), .A2(n_852), .B1(n_888), .B2(n_890), .Y(n_887) );
CKINVDCx6p67_ASAP7_75t_R g854 ( .A(n_855), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_859), .B1(n_860), .B2(n_861), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_857), .A2(n_1140), .B1(n_1149), .B2(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g1174 ( .A1(n_860), .A2(n_1175), .B1(n_1176), .B2(n_1177), .Y(n_1174) );
OAI21xp5_ASAP7_75t_SL g862 ( .A1(n_863), .A2(n_864), .B(n_865), .Y(n_862) );
OAI22xp33_ASAP7_75t_L g1131 ( .A1(n_863), .A2(n_1106), .B1(n_1111), .B2(n_1132), .Y(n_1131) );
OAI221xp5_ASAP7_75t_L g1368 ( .A1(n_863), .A2(n_1014), .B1(n_1369), .B2(n_1370), .C(n_1371), .Y(n_1368) );
CKINVDCx8_ASAP7_75t_R g1156 ( .A(n_867), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_870), .B(n_972), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g1668 ( .A(n_870), .B(n_1669), .Y(n_1668) );
INVx1_ASAP7_75t_L g1380 ( .A(n_872), .Y(n_1380) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_882), .B1(n_884), .B2(n_892), .C(n_893), .Y(n_874) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g1088 ( .A(n_881), .Y(n_1088) );
INVx1_ASAP7_75t_L g1153 ( .A(n_881), .Y(n_1153) );
INVx1_ASAP7_75t_L g976 ( .A(n_882), .Y(n_976) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g1345 ( .A(n_883), .Y(n_1345) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx4_ASAP7_75t_L g986 ( .A(n_892), .Y(n_986) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_902), .B1(n_903), .B2(n_904), .C(n_905), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g1388 ( .A1(n_899), .A2(n_1373), .B1(n_1376), .B2(n_1389), .Y(n_1388) );
AOI221xp5_ASAP7_75t_L g1681 ( .A1(n_899), .A2(n_903), .B1(n_1682), .B2(n_1683), .C(n_1684), .Y(n_1681) );
AND2x2_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
XNOR2x1_ASAP7_75t_SL g906 ( .A(n_907), .B(n_908), .Y(n_906) );
AND2x2_ASAP7_75t_L g908 ( .A(n_909), .B(n_943), .Y(n_908) );
NOR3xp33_ASAP7_75t_SL g909 ( .A(n_910), .B(n_918), .C(n_920), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_914), .Y(n_910) );
OAI221xp5_ASAP7_75t_L g953 ( .A1(n_913), .A2(n_915), .B1(n_954), .B2(n_955), .C(n_956), .Y(n_953) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
OAI22xp33_ASAP7_75t_L g1181 ( .A1(n_926), .A2(n_1132), .B1(n_1139), .B2(n_1144), .Y(n_1181) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_928), .A2(n_929), .B1(n_931), .B2(n_932), .Y(n_927) );
INVx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g1063 ( .A(n_930), .Y(n_1063) );
INVx2_ASAP7_75t_L g1130 ( .A(n_930), .Y(n_1130) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
NAND3xp33_ASAP7_75t_L g944 ( .A(n_945), .B(n_958), .C(n_965), .Y(n_944) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
BUFx2_ASAP7_75t_L g1347 ( .A(n_951), .Y(n_1347) );
BUFx3_ASAP7_75t_L g1354 ( .A(n_951), .Y(n_1354) );
OAI221xp5_ASAP7_75t_L g1673 ( .A1(n_955), .A2(n_1196), .B1(n_1665), .B2(n_1666), .C(n_1674), .Y(n_1673) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
XNOR2xp5_ASAP7_75t_L g968 ( .A(n_969), .B(n_970), .Y(n_968) );
AND4x1_ASAP7_75t_L g970 ( .A(n_971), .B(n_973), .C(n_995), .D(n_1025), .Y(n_970) );
NOR3xp33_ASAP7_75t_SL g973 ( .A(n_974), .B(n_975), .C(n_993), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_977), .B1(n_986), .B2(n_987), .Y(n_975) );
INVx2_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g1356 ( .A(n_986), .Y(n_1356) );
INVx2_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
OAI31xp33_ASAP7_75t_L g995 ( .A1(n_996), .A2(n_1011), .A3(n_1021), .B(n_1024), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_1006), .A2(n_1007), .B1(n_1009), .B2(n_1010), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx2_ASAP7_75t_SL g1018 ( .A(n_1019), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1028), .Y(n_1025) );
CKINVDCx6p67_ASAP7_75t_R g1387 ( .A(n_1027), .Y(n_1387) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1238), .B1(n_1391), .B2(n_1392), .Y(n_1032) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1033), .Y(n_1392) );
AO22x1_ASAP7_75t_L g1033 ( .A1(n_1034), .A2(n_1035), .B1(n_1133), .B2(n_1237), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
AO22x2_ASAP7_75t_L g1035 ( .A1(n_1036), .A2(n_1037), .B1(n_1091), .B2(n_1092), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
XNOR2xp5_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1039), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1071), .Y(n_1039) );
NOR3xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1048), .C(n_1050), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1045), .Y(n_1041) );
OAI22xp33_ASAP7_75t_L g1051 ( .A1(n_1052), .A2(n_1053), .B1(n_1054), .B2(n_1055), .Y(n_1051) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1064), .B1(n_1065), .B2(n_1067), .Y(n_1062) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
NAND3xp33_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1079), .C(n_1089), .Y(n_1073) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1083), .Y(n_1108) );
BUFx6f_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1114), .Y(n_1093) );
NAND3xp33_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1105), .C(n_1110), .Y(n_1095) );
NOR3xp33_ASAP7_75t_SL g1114 ( .A(n_1115), .B(n_1121), .C(n_1122), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1119), .Y(n_1115) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1133), .Y(n_1237) );
XOR2x2_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1184), .Y(n_1133) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1135), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1158), .Y(n_1135) );
NAND3xp33_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1141), .C(n_1148), .Y(n_1137) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
NOR3xp33_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1167), .C(n_1168), .Y(n_1158) );
NAND2xp5_ASAP7_75t_SL g1159 ( .A(n_1160), .B(n_1164), .Y(n_1159) );
INVx2_ASAP7_75t_L g1233 ( .A(n_1162), .Y(n_1233) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1365 ( .A1(n_1175), .A2(n_1303), .B1(n_1366), .B2(n_1367), .Y(n_1365) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1185), .Y(n_1236) );
NAND4xp75_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1187), .C(n_1213), .D(n_1229), .Y(n_1185) );
OAI31xp33_ASAP7_75t_L g1187 ( .A1(n_1188), .A2(n_1200), .A3(n_1210), .B(n_1211), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_1190), .A2(n_1191), .B1(n_1192), .B2(n_1193), .Y(n_1189) );
OAI21xp33_ASAP7_75t_L g1194 ( .A1(n_1195), .A2(n_1196), .B(n_1198), .Y(n_1194) );
OAI221xp5_ASAP7_75t_L g1675 ( .A1(n_1196), .A2(n_1676), .B1(n_1678), .B2(n_1679), .C(n_1680), .Y(n_1675) );
INVx2_ASAP7_75t_SL g1196 ( .A(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1197), .Y(n_1207) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1197), .Y(n_1323) );
OAI211xp5_ASAP7_75t_L g1205 ( .A1(n_1206), .A2(n_1207), .B(n_1208), .C(n_1209), .Y(n_1205) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
AOI31xp33_ASAP7_75t_SL g1265 ( .A1(n_1212), .A2(n_1266), .A3(n_1270), .B(n_1273), .Y(n_1265) );
AND2x2_ASAP7_75t_SL g1213 ( .A(n_1214), .B(n_1228), .Y(n_1213) );
AOI33xp33_ASAP7_75t_L g1214 ( .A1(n_1215), .A2(n_1216), .A3(n_1218), .B1(n_1222), .B2(n_1224), .B3(n_1227), .Y(n_1214) );
AOI22xp5_ASAP7_75t_L g1249 ( .A1(n_1215), .A2(n_1250), .B1(n_1254), .B2(n_1255), .Y(n_1249) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1238), .Y(n_1391) );
AOI22xp5_ASAP7_75t_L g1238 ( .A1(n_1239), .A2(n_1338), .B1(n_1339), .B2(n_1390), .Y(n_1238) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1239), .Y(n_1390) );
AOI22xp5_ASAP7_75t_L g1239 ( .A1(n_1240), .A2(n_1241), .B1(n_1283), .B2(n_1337), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
HB1xp67_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
NAND2xp5_ASAP7_75t_SL g1243 ( .A(n_1244), .B(n_1279), .Y(n_1243) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1245), .Y(n_1281) );
NAND3xp33_ASAP7_75t_SL g1245 ( .A(n_1246), .B(n_1249), .C(n_1256), .Y(n_1245) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1265), .Y(n_1280) );
NAND3xp33_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1281), .C(n_1282), .Y(n_1279) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1283), .Y(n_1337) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_SL g1336 ( .A(n_1285), .Y(n_1336) );
NAND4xp75_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1307), .C(n_1311), .D(n_1332), .Y(n_1285) );
OAI22xp5_ASAP7_75t_L g1287 ( .A1(n_1288), .A2(n_1289), .B1(n_1290), .B2(n_1291), .Y(n_1287) );
OAI22xp5_ASAP7_75t_L g1660 ( .A1(n_1289), .A2(n_1661), .B1(n_1662), .B2(n_1663), .Y(n_1660) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
OAI211xp5_ASAP7_75t_L g1322 ( .A1(n_1295), .A2(n_1323), .B(n_1324), .C(n_1326), .Y(n_1322) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_1300), .A2(n_1301), .B1(n_1302), .B2(n_1303), .Y(n_1299) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
NOR2x1_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1310), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1322), .Y(n_1316) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
BUFx2_ASAP7_75t_L g1339 ( .A(n_1340), .Y(n_1339) );
BUFx2_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
NAND4xp75_ASAP7_75t_L g1342 ( .A(n_1343), .B(n_1361), .C(n_1386), .D(n_1388), .Y(n_1342) );
AND2x2_ASAP7_75t_SL g1343 ( .A(n_1344), .B(n_1357), .Y(n_1343) );
AOI33xp33_ASAP7_75t_L g1344 ( .A1(n_1345), .A2(n_1346), .A3(n_1349), .B1(n_1352), .B2(n_1353), .B3(n_1356), .Y(n_1344) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
OAI221xp5_ASAP7_75t_L g1364 ( .A1(n_1365), .A2(n_1368), .B1(n_1372), .B2(n_1375), .C(n_1379), .Y(n_1364) );
AOI21xp5_ASAP7_75t_L g1379 ( .A1(n_1380), .A2(n_1381), .B(n_1382), .Y(n_1379) );
OAI221xp5_ASAP7_75t_L g1394 ( .A1(n_1395), .A2(n_1644), .B1(n_1646), .B2(n_1686), .C(n_1690), .Y(n_1394) );
AOI211xp5_ASAP7_75t_L g1395 ( .A1(n_1396), .A2(n_1552), .B(n_1594), .C(n_1626), .Y(n_1395) );
NAND5xp2_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1494), .C(n_1512), .D(n_1541), .E(n_1544), .Y(n_1396) );
AOI321xp33_ASAP7_75t_L g1397 ( .A1(n_1398), .A2(n_1441), .A3(n_1458), .B1(n_1465), .B2(n_1473), .C(n_1484), .Y(n_1397) );
NAND2xp5_ASAP7_75t_L g1398 ( .A(n_1399), .B(n_1437), .Y(n_1398) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1424), .Y(n_1400) );
CKINVDCx6p67_ASAP7_75t_R g1440 ( .A(n_1401), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1401), .B(n_1439), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1486 ( .A(n_1401), .B(n_1487), .Y(n_1486) );
OR2x2_ASAP7_75t_L g1503 ( .A(n_1401), .B(n_1439), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1401), .B(n_1510), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1401), .B(n_1537), .Y(n_1547) );
OR2x2_ASAP7_75t_L g1551 ( .A(n_1401), .B(n_1488), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1401), .B(n_1425), .Y(n_1581) );
A2O1A1Ixp33_ASAP7_75t_SL g1630 ( .A1(n_1401), .A2(n_1631), .B(n_1635), .C(n_1637), .Y(n_1630) );
OR2x6_ASAP7_75t_SL g1401 ( .A(n_1402), .B(n_1414), .Y(n_1401) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1410), .B1(n_1411), .B2(n_1413), .Y(n_1402) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1407), .Y(n_1404) );
AND2x4_ASAP7_75t_L g1412 ( .A(n_1405), .B(n_1408), .Y(n_1412) );
AND2x4_ASAP7_75t_L g1453 ( .A(n_1405), .B(n_1407), .Y(n_1453) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1406), .Y(n_1419) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1409), .B(n_1419), .Y(n_1418) );
OAI22xp5_ASAP7_75t_L g1450 ( .A1(n_1411), .A2(n_1451), .B1(n_1452), .B2(n_1454), .Y(n_1450) );
INVx1_ASAP7_75t_SL g1411 ( .A(n_1412), .Y(n_1411) );
INVx2_ASAP7_75t_L g1464 ( .A(n_1412), .Y(n_1464) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_1415), .A2(n_1420), .B1(n_1421), .B2(n_1423), .Y(n_1414) );
OAI22xp33_ASAP7_75t_L g1445 ( .A1(n_1415), .A2(n_1446), .B1(n_1447), .B2(n_1448), .Y(n_1445) );
OAI22xp33_ASAP7_75t_L g1468 ( .A1(n_1415), .A2(n_1421), .B1(n_1469), .B2(n_1470), .Y(n_1468) );
BUFx3_ASAP7_75t_L g1527 ( .A(n_1415), .Y(n_1527) );
BUFx6f_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
OAI22xp5_ASAP7_75t_L g1434 ( .A1(n_1416), .A2(n_1421), .B1(n_1435), .B2(n_1436), .Y(n_1434) );
OR2x2_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1418), .Y(n_1416) );
OR2x2_ASAP7_75t_L g1421 ( .A(n_1417), .B(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1417), .Y(n_1429) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1418), .Y(n_1428) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1421), .Y(n_1449) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1422), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1424), .B(n_1483), .Y(n_1482) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1424), .Y(n_1489) );
OAI32xp33_ASAP7_75t_L g1556 ( .A1(n_1424), .A2(n_1455), .A3(n_1495), .B1(n_1557), .B2(n_1559), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1424), .B(n_1440), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g1606 ( .A(n_1424), .B(n_1499), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1433), .Y(n_1424) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1425), .Y(n_1439) );
OR2x2_ASAP7_75t_L g1488 ( .A(n_1425), .B(n_1433), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1425), .B(n_1511), .Y(n_1510) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1432), .Y(n_1425) );
AND2x4_ASAP7_75t_L g1427 ( .A(n_1428), .B(n_1429), .Y(n_1427) );
OAI21xp33_ASAP7_75t_SL g1701 ( .A1(n_1428), .A2(n_1694), .B(n_1702), .Y(n_1701) );
AND2x4_ASAP7_75t_L g1430 ( .A(n_1429), .B(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1433), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1433), .B(n_1440), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1537 ( .A(n_1433), .B(n_1439), .Y(n_1537) );
OAI221xp5_ASAP7_75t_L g1513 ( .A1(n_1437), .A2(n_1472), .B1(n_1514), .B2(n_1516), .C(n_1519), .Y(n_1513) );
O2A1O1Ixp33_ASAP7_75t_L g1575 ( .A1(n_1437), .A2(n_1539), .B(n_1576), .C(n_1577), .Y(n_1575) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
A2O1A1Ixp33_ASAP7_75t_L g1590 ( .A1(n_1438), .A2(n_1459), .B(n_1548), .C(n_1591), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1439), .B(n_1440), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1440), .B(n_1460), .Y(n_1499) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_1440), .B(n_1537), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1440), .B(n_1510), .Y(n_1543) );
NOR2xp33_ASAP7_75t_L g1558 ( .A(n_1440), .B(n_1460), .Y(n_1558) );
OR2x2_ASAP7_75t_L g1561 ( .A(n_1440), .B(n_1511), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1440), .B(n_1482), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1440), .B(n_1511), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_1441), .B(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
OAI22xp5_ASAP7_75t_SL g1599 ( .A1(n_1442), .A2(n_1508), .B1(n_1600), .B2(n_1601), .Y(n_1599) );
OR2x2_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1455), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1471 ( .A(n_1443), .B(n_1472), .Y(n_1471) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1443), .Y(n_1478) );
INVx3_ASAP7_75t_L g1540 ( .A(n_1443), .Y(n_1540) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1443), .B(n_1535), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1443), .B(n_1505), .Y(n_1586) );
AOI221xp5_ASAP7_75t_L g1603 ( .A1(n_1443), .A2(n_1604), .B1(n_1605), .B2(n_1607), .C(n_1611), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1443), .B(n_1455), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1637 ( .A(n_1443), .B(n_1493), .Y(n_1637) );
INVx3_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
OR2x2_ASAP7_75t_L g1550 ( .A(n_1444), .B(n_1480), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1444), .B(n_1455), .Y(n_1614) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1450), .Y(n_1444) );
HB1xp67_ASAP7_75t_L g1529 ( .A(n_1448), .Y(n_1529) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1453), .Y(n_1523) );
INVx2_ASAP7_75t_L g1472 ( .A(n_1455), .Y(n_1472) );
OR2x2_ASAP7_75t_L g1480 ( .A(n_1455), .B(n_1467), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1455), .B(n_1467), .Y(n_1493) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1455), .B(n_1502), .Y(n_1501) );
OR2x2_ASAP7_75t_L g1507 ( .A(n_1455), .B(n_1505), .Y(n_1507) );
AND2x2_ASAP7_75t_L g1515 ( .A(n_1455), .B(n_1505), .Y(n_1515) );
AND2x4_ASAP7_75t_L g1455 ( .A(n_1456), .B(n_1457), .Y(n_1455) );
NOR2x1_ASAP7_75t_L g1560 ( .A(n_1458), .B(n_1561), .Y(n_1560) );
NAND2xp5_ASAP7_75t_L g1563 ( .A(n_1458), .B(n_1475), .Y(n_1563) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1458), .B(n_1547), .Y(n_1566) );
OR2x2_ASAP7_75t_L g1577 ( .A(n_1458), .B(n_1507), .Y(n_1577) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1458), .B(n_1565), .Y(n_1600) );
INVx2_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1459), .B(n_1518), .Y(n_1517) );
NAND2xp5_ASAP7_75t_L g1533 ( .A(n_1459), .B(n_1534), .Y(n_1533) );
NAND2xp5_ASAP7_75t_L g1546 ( .A(n_1459), .B(n_1547), .Y(n_1546) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1459), .B(n_1640), .Y(n_1639) );
INVx2_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx4_ASAP7_75t_L g1483 ( .A(n_1460), .Y(n_1483) );
NAND2xp5_ASAP7_75t_L g1504 ( .A(n_1460), .B(n_1505), .Y(n_1504) );
OR2x2_ASAP7_75t_L g1555 ( .A(n_1460), .B(n_1488), .Y(n_1555) );
NAND2xp5_ASAP7_75t_L g1576 ( .A(n_1460), .B(n_1535), .Y(n_1576) );
OR2x2_ASAP7_75t_L g1622 ( .A(n_1460), .B(n_1534), .Y(n_1622) );
NAND2xp5_ASAP7_75t_L g1629 ( .A(n_1460), .B(n_1509), .Y(n_1629) );
OR2x2_ASAP7_75t_L g1636 ( .A(n_1460), .B(n_1551), .Y(n_1636) );
AND2x6_ASAP7_75t_L g1460 ( .A(n_1461), .B(n_1462), .Y(n_1460) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
OAI22xp5_ASAP7_75t_L g1521 ( .A1(n_1464), .A2(n_1522), .B1(n_1523), .B2(n_1524), .Y(n_1521) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1465), .Y(n_1604) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1466), .B(n_1471), .Y(n_1465) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1466), .Y(n_1598) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1466), .B(n_1602), .Y(n_1601) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1466), .Y(n_1608) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1466), .Y(n_1625) );
HB1xp67_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
INVx2_ASAP7_75t_SL g1505 ( .A(n_1467), .Y(n_1505) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1472), .Y(n_1496) );
OAI22xp5_ASAP7_75t_L g1473 ( .A1(n_1474), .A2(n_1476), .B1(n_1478), .B2(n_1481), .Y(n_1473) );
INVxp67_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1475), .B(n_1483), .Y(n_1573) );
INVxp67_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1478), .B(n_1479), .Y(n_1477) );
AOI21xp5_ASAP7_75t_L g1589 ( .A1(n_1478), .A2(n_1497), .B(n_1519), .Y(n_1589) );
AOI22xp5_ASAP7_75t_L g1615 ( .A1(n_1478), .A2(n_1616), .B1(n_1619), .B2(n_1623), .Y(n_1615) );
OAI211xp5_ASAP7_75t_L g1552 ( .A1(n_1479), .A2(n_1553), .B(n_1564), .C(n_1578), .Y(n_1552) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVxp67_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1483), .Y(n_1492) );
NAND2xp5_ASAP7_75t_L g1514 ( .A(n_1483), .B(n_1515), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1483), .B(n_1543), .Y(n_1542) );
AOI21xp5_ASAP7_75t_L g1484 ( .A1(n_1485), .A2(n_1489), .B(n_1490), .Y(n_1484) );
AND2x2_ASAP7_75t_L g1617 ( .A(n_1485), .B(n_1618), .Y(n_1617) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
OAI31xp33_ASAP7_75t_L g1638 ( .A1(n_1486), .A2(n_1517), .A3(n_1639), .B(n_1641), .Y(n_1638) );
NAND2xp5_ASAP7_75t_L g1498 ( .A(n_1487), .B(n_1499), .Y(n_1498) );
NAND2xp5_ASAP7_75t_L g1610 ( .A(n_1487), .B(n_1558), .Y(n_1610) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1493), .Y(n_1491) );
NAND2xp5_ASAP7_75t_L g1580 ( .A(n_1492), .B(n_1581), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1492), .B(n_1510), .Y(n_1591) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1493), .Y(n_1593) );
AOI211xp5_ASAP7_75t_SL g1494 ( .A1(n_1495), .A2(n_1497), .B(n_1500), .C(n_1506), .Y(n_1494) );
OAI22xp5_ASAP7_75t_L g1579 ( .A1(n_1495), .A2(n_1580), .B1(n_1582), .B2(n_1583), .Y(n_1579) );
AOI21xp5_ASAP7_75t_L g1595 ( .A1(n_1495), .A2(n_1596), .B(n_1599), .Y(n_1595) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g1597 ( .A(n_1497), .B(n_1598), .Y(n_1597) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
OR2x2_ASAP7_75t_L g1624 ( .A(n_1498), .B(n_1625), .Y(n_1624) );
INVxp67_ASAP7_75t_SL g1500 ( .A(n_1501), .Y(n_1500) );
INVxp33_ASAP7_75t_L g1612 ( .A(n_1502), .Y(n_1612) );
NOR2xp33_ASAP7_75t_L g1502 ( .A(n_1503), .B(n_1504), .Y(n_1502) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1503), .Y(n_1640) );
INVx2_ASAP7_75t_SL g1535 ( .A(n_1505), .Y(n_1535) );
NOR2xp33_ASAP7_75t_L g1506 ( .A(n_1507), .B(n_1508), .Y(n_1506) );
INVx2_ASAP7_75t_L g1565 ( .A(n_1507), .Y(n_1565) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
OAI21xp33_ASAP7_75t_SL g1572 ( .A1(n_1509), .A2(n_1573), .B(n_1574), .Y(n_1572) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1510), .Y(n_1633) );
OAI21xp5_ASAP7_75t_L g1512 ( .A1(n_1513), .A2(n_1530), .B(n_1538), .Y(n_1512) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1515), .Y(n_1582) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
INVxp67_ASAP7_75t_L g1583 ( .A(n_1518), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1538 ( .A(n_1519), .B(n_1539), .Y(n_1538) );
CKINVDCx5p33_ASAP7_75t_R g1519 ( .A(n_1520), .Y(n_1519) );
OR2x6_ASAP7_75t_SL g1520 ( .A(n_1521), .B(n_1525), .Y(n_1520) );
OAI22xp5_ASAP7_75t_L g1525 ( .A1(n_1526), .A2(n_1527), .B1(n_1528), .B2(n_1529), .Y(n_1525) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1527), .Y(n_1645) );
INVxp67_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
NAND2xp5_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1536), .Y(n_1531) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
AOI221xp5_ASAP7_75t_L g1553 ( .A1(n_1535), .A2(n_1540), .B1(n_1554), .B2(n_1556), .C(n_1562), .Y(n_1553) );
NOR2xp33_ASAP7_75t_L g1562 ( .A(n_1535), .B(n_1563), .Y(n_1562) );
NAND2xp5_ASAP7_75t_L g1571 ( .A(n_1535), .B(n_1555), .Y(n_1571) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1535), .Y(n_1643) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1537), .Y(n_1634) );
AOI211xp5_ASAP7_75t_L g1578 ( .A1(n_1539), .A2(n_1579), .B(n_1584), .C(n_1592), .Y(n_1578) );
NOR2xp33_ASAP7_75t_L g1621 ( .A(n_1539), .B(n_1622), .Y(n_1621) );
INVx1_ASAP7_75t_SL g1539 ( .A(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1543), .Y(n_1618) );
AOI21xp5_ASAP7_75t_L g1544 ( .A1(n_1545), .A2(n_1548), .B(n_1549), .Y(n_1544) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
NOR2xp33_ASAP7_75t_L g1549 ( .A(n_1550), .B(n_1551), .Y(n_1549) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1550), .Y(n_1574) );
NOR2xp33_ASAP7_75t_L g1592 ( .A(n_1551), .B(n_1593), .Y(n_1592) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
AOI211xp5_ASAP7_75t_L g1564 ( .A1(n_1565), .A2(n_1566), .B(n_1567), .C(n_1575), .Y(n_1564) );
OAI21xp33_ASAP7_75t_L g1567 ( .A1(n_1568), .A2(n_1570), .B(n_1572), .Y(n_1567) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
INVxp67_ASAP7_75t_SL g1570 ( .A(n_1571), .Y(n_1570) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_1577), .B(n_1620), .Y(n_1619) );
OAI211xp5_ASAP7_75t_L g1584 ( .A1(n_1585), .A2(n_1587), .B(n_1589), .C(n_1590), .Y(n_1584) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
AOI21xp33_ASAP7_75t_SL g1611 ( .A1(n_1587), .A2(n_1612), .B(n_1613), .Y(n_1611) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
NAND3xp33_ASAP7_75t_L g1594 ( .A(n_1595), .B(n_1603), .C(n_1615), .Y(n_1594) );
INVxp67_ASAP7_75t_SL g1596 ( .A(n_1597), .Y(n_1596) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1608), .B(n_1609), .Y(n_1607) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
INVxp67_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
INVxp67_ASAP7_75t_SL g1620 ( .A(n_1621), .Y(n_1620) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
OAI211xp5_ASAP7_75t_L g1626 ( .A1(n_1627), .A2(n_1629), .B(n_1630), .C(n_1638), .Y(n_1626) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1628), .Y(n_1627) );
NAND2xp5_ASAP7_75t_L g1642 ( .A(n_1628), .B(n_1643), .Y(n_1642) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1633), .B(n_1634), .Y(n_1632) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
CKINVDCx16_ASAP7_75t_R g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
HB1xp67_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1649), .Y(n_1685) );
NAND4xp25_ASAP7_75t_L g1649 ( .A(n_1650), .B(n_1668), .C(n_1670), .D(n_1681), .Y(n_1649) );
AOI21xp5_ASAP7_75t_L g1655 ( .A1(n_1656), .A2(n_1657), .B(n_1658), .Y(n_1655) );
INVx2_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
HB1xp67_ASAP7_75t_L g1698 ( .A(n_1685), .Y(n_1698) );
INVx2_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
CKINVDCx5p33_ASAP7_75t_R g1692 ( .A(n_1693), .Y(n_1692) );
INVxp33_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1698), .Y(n_1699) );
HB1xp67_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
endmodule