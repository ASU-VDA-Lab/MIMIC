module fake_jpeg_29730_n_112 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_51),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_48),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_15),
.B1(n_35),
.B2(n_34),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_46),
.B1(n_39),
.B2(n_41),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_1),
.B(n_3),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_3),
.Y(n_61)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_48),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_69),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_4),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_40),
.B1(n_43),
.B2(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_4),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_68),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_47),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_73),
.B1(n_76),
.B2(n_80),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_40),
.B1(n_45),
.B2(n_16),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_14),
.C(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_77),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_36),
.B1(n_31),
.B2(n_30),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_82),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_29),
.B1(n_28),
.B2(n_23),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_19),
.A3(n_17),
.B1(n_6),
.B2(n_7),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_76),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_69),
.B1(n_58),
.B2(n_65),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_58),
.B(n_6),
.C(n_7),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_72),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_92),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_94),
.B1(n_96),
.B2(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_5),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_8),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_73),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_71),
.C(n_10),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_101),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_10),
.C(n_11),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_102),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_97),
.B(n_85),
.C(n_87),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_85),
.B(n_100),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_99),
.C(n_102),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_106),
.A2(n_107),
.B(n_103),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_98),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_87),
.B1(n_95),
.B2(n_91),
.Y(n_110)
);

AOI322xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_87),
.C1(n_95),
.C2(n_104),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_111),
.Y(n_112)
);


endmodule