module fake_netlist_1_2108_n_1472 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1472);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1472;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_386;
wire n_659;
wire n_432;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1439;
wire n_374;
wire n_718;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_250), .Y(n_344) );
INVxp33_ASAP7_75t_SL g345 ( .A(n_68), .Y(n_345) );
INVxp33_ASAP7_75t_SL g346 ( .A(n_64), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_92), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_71), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_127), .Y(n_349) );
CKINVDCx14_ASAP7_75t_R g350 ( .A(n_113), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_223), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_331), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_30), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_332), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_309), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_107), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_172), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_185), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_80), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_174), .Y(n_360) );
INVxp33_ASAP7_75t_SL g361 ( .A(n_192), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_87), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_53), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_212), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_195), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_75), .Y(n_366) );
INVxp33_ASAP7_75t_L g367 ( .A(n_334), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_81), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_208), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_253), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_307), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_56), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_1), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_89), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_148), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_19), .Y(n_376) );
INVxp33_ASAP7_75t_SL g377 ( .A(n_342), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_244), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_292), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_278), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_63), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_264), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_215), .Y(n_383) );
INVxp33_ASAP7_75t_L g384 ( .A(n_255), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_32), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_82), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_38), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_56), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_160), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_16), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_218), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_330), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_62), .Y(n_393) );
INVxp67_ASAP7_75t_SL g394 ( .A(n_14), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_64), .Y(n_395) );
CKINVDCx14_ASAP7_75t_R g396 ( .A(n_299), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_273), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_90), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_282), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_135), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_211), .Y(n_401) );
CKINVDCx14_ASAP7_75t_R g402 ( .A(n_260), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_128), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_240), .B(n_177), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_193), .Y(n_405) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_33), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_52), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_28), .Y(n_408) );
CKINVDCx14_ASAP7_75t_R g409 ( .A(n_270), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g410 ( .A(n_229), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_322), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_335), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_10), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_29), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_38), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_109), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_47), .Y(n_417) );
INVxp33_ASAP7_75t_L g418 ( .A(n_176), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_235), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_252), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_184), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_65), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_52), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_257), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_243), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_78), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_221), .Y(n_427) );
BUFx3_ASAP7_75t_L g428 ( .A(n_317), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_18), .Y(n_429) );
INVx2_ASAP7_75t_SL g430 ( .A(n_258), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_327), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_222), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_324), .Y(n_433) );
INVx1_ASAP7_75t_SL g434 ( .A(n_29), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_261), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_202), .Y(n_436) );
INVxp67_ASAP7_75t_L g437 ( .A(n_207), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_256), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_101), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_161), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_74), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_275), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_333), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_201), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_225), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_84), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_216), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_186), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_228), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_166), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_205), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_279), .Y(n_452) );
INVx4_ASAP7_75t_R g453 ( .A(n_269), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_114), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_180), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_117), .Y(n_456) );
INVxp33_ASAP7_75t_L g457 ( .A(n_20), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_62), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_102), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_110), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_266), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_140), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_129), .B(n_144), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_0), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_112), .Y(n_465) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_162), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_48), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_111), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_343), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_74), .Y(n_470) );
CKINVDCx14_ASAP7_75t_R g471 ( .A(n_167), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_226), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_182), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_73), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_67), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_262), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_147), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_100), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_12), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_220), .Y(n_480) );
INVxp33_ASAP7_75t_SL g481 ( .A(n_42), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_171), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_173), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_106), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_75), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_123), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_311), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_115), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_198), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_122), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_233), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_283), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_339), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_158), .Y(n_494) );
INVxp33_ASAP7_75t_L g495 ( .A(n_150), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_95), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_83), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_178), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_2), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_267), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_217), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_248), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_100), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_131), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_12), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_70), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_164), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g508 ( .A(n_98), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_316), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_305), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_136), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_312), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_230), .Y(n_513) );
INVx3_ASAP7_75t_L g514 ( .A(n_423), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_513), .B(n_0), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_382), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_513), .B(n_1), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_391), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_382), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_383), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_356), .Y(n_521) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_356), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_383), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_356), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_389), .Y(n_525) );
AND3x2_ASAP7_75t_L g526 ( .A(n_353), .B(n_2), .C(n_3), .Y(n_526) );
XNOR2xp5_ASAP7_75t_L g527 ( .A(n_347), .B(n_3), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_389), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_356), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_502), .Y(n_530) );
CKINVDCx11_ASAP7_75t_R g531 ( .A(n_347), .Y(n_531) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_356), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_502), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_423), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_358), .Y(n_535) );
NOR2xp33_ASAP7_75t_SL g536 ( .A(n_344), .B(n_105), .Y(n_536) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_391), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_430), .B(n_4), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_386), .Y(n_539) );
INVx4_ASAP7_75t_L g540 ( .A(n_423), .Y(n_540) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_428), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_353), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_358), .Y(n_543) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_428), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_457), .B(n_4), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_386), .Y(n_546) );
BUFx2_ASAP7_75t_L g547 ( .A(n_439), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_369), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_390), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_390), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_413), .Y(n_551) );
NOR2xp33_ASAP7_75t_SL g552 ( .A(n_410), .B(n_108), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_547), .B(n_430), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_542), .B(n_457), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_547), .B(n_357), .Y(n_555) );
BUFx3_ASAP7_75t_L g556 ( .A(n_538), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_531), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_538), .B(n_369), .Y(n_558) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_522), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_517), .B(n_512), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_517), .B(n_474), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_532), .Y(n_562) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_522), .Y(n_563) );
INVx2_ASAP7_75t_SL g564 ( .A(n_518), .Y(n_564) );
OAI221xp5_ASAP7_75t_L g565 ( .A1(n_542), .A2(n_406), .B1(n_394), .B2(n_376), .C(n_387), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_532), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_535), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_545), .Y(n_568) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_522), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_547), .B(n_367), .Y(n_570) );
BUFx3_ASAP7_75t_L g571 ( .A(n_538), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_545), .B(n_367), .Y(n_572) );
INVx5_ASAP7_75t_L g573 ( .A(n_522), .Y(n_573) );
NAND2x1p5_ASAP7_75t_L g574 ( .A(n_517), .B(n_349), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_540), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_517), .B(n_474), .Y(n_576) );
INVx4_ASAP7_75t_SL g577 ( .A(n_538), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_535), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_538), .B(n_400), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_516), .B(n_384), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_532), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_516), .B(n_400), .Y(n_582) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_522), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_535), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_532), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_519), .B(n_370), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_543), .Y(n_587) );
INVx3_ASAP7_75t_L g588 ( .A(n_540), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_532), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_532), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_543), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_519), .B(n_416), .Y(n_592) );
AOI21x1_ASAP7_75t_L g593 ( .A1(n_521), .A2(n_431), .B(n_416), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_532), .Y(n_594) );
NOR2x1p5_ASAP7_75t_L g595 ( .A(n_515), .B(n_362), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_522), .Y(n_596) );
INVx2_ASAP7_75t_SL g597 ( .A(n_518), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_517), .B(n_439), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_557), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_572), .A2(n_545), .B1(n_552), .B2(n_536), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_577), .B(n_536), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g602 ( .A(n_572), .B(n_381), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_572), .A2(n_552), .B1(n_515), .B2(n_346), .Y(n_603) );
NOR2xp67_ASAP7_75t_L g604 ( .A(n_565), .B(n_520), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_580), .B(n_520), .Y(n_605) );
O2A1O1Ixp5_ASAP7_75t_L g606 ( .A1(n_558), .A2(n_418), .B(n_495), .C(n_384), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_580), .B(n_523), .Y(n_607) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_556), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_568), .Y(n_609) );
OR2x2_ASAP7_75t_SL g610 ( .A(n_555), .B(n_531), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_570), .Y(n_611) );
BUFx2_ASAP7_75t_L g612 ( .A(n_554), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_568), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_593), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_554), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_593), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_561), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_570), .B(n_586), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_570), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_577), .B(n_523), .Y(n_620) );
OR2x6_ASAP7_75t_L g621 ( .A(n_560), .B(n_527), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_555), .Y(n_622) );
BUFx3_ASAP7_75t_L g623 ( .A(n_556), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_586), .B(n_525), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_593), .Y(n_625) );
INVxp67_ASAP7_75t_L g626 ( .A(n_553), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_556), .A2(n_528), .B1(n_530), .B2(n_525), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_561), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_556), .Y(n_629) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_571), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_553), .B(n_528), .Y(n_631) );
INVx4_ASAP7_75t_L g632 ( .A(n_577), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_560), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_560), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_598), .B(n_530), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_571), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_595), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_598), .B(n_533), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_561), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_595), .Y(n_640) );
OR2x6_ASAP7_75t_L g641 ( .A(n_560), .B(n_527), .Y(n_641) );
BUFx3_ASAP7_75t_L g642 ( .A(n_571), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_561), .Y(n_643) );
INVx2_ASAP7_75t_SL g644 ( .A(n_574), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_577), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_577), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_561), .B(n_533), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_577), .B(n_504), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_576), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_576), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_576), .Y(n_651) );
INVx2_ASAP7_75t_SL g652 ( .A(n_574), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_565), .B(n_508), .Y(n_653) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_574), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_576), .A2(n_346), .B1(n_481), .B2(n_345), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_576), .B(n_418), .Y(n_656) );
NOR2xp67_ASAP7_75t_L g657 ( .A(n_567), .B(n_449), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_567), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_574), .B(n_351), .Y(n_659) );
INVx3_ASAP7_75t_SL g660 ( .A(n_598), .Y(n_660) );
BUFx3_ASAP7_75t_L g661 ( .A(n_564), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_578), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_598), .B(n_352), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_598), .A2(n_481), .B1(n_345), .B2(n_397), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_558), .B(n_518), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_578), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_579), .A2(n_397), .B1(n_424), .B2(n_360), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_579), .B(n_518), .Y(n_668) );
NOR2xp67_ASAP7_75t_L g669 ( .A(n_584), .B(n_480), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_584), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_587), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_587), .B(n_495), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_591), .B(n_489), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_591), .Y(n_674) );
BUFx4f_ASAP7_75t_SL g675 ( .A(n_582), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_582), .B(n_526), .Y(n_676) );
BUFx3_ASAP7_75t_L g677 ( .A(n_564), .Y(n_677) );
INVx5_ASAP7_75t_L g678 ( .A(n_575), .Y(n_678) );
OR2x6_ASAP7_75t_L g679 ( .A(n_592), .B(n_527), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_564), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_592), .Y(n_681) );
BUFx12f_ASAP7_75t_L g682 ( .A(n_597), .Y(n_682) );
INVx2_ASAP7_75t_SL g683 ( .A(n_644), .Y(n_683) );
BUFx12f_ASAP7_75t_L g684 ( .A(n_599), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_611), .A2(n_377), .B1(n_361), .B2(n_499), .Y(n_685) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_652), .Y(n_686) );
BUFx3_ASAP7_75t_L g687 ( .A(n_646), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_658), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_658), .Y(n_689) );
BUFx6f_ASAP7_75t_SL g690 ( .A(n_621), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_618), .A2(n_377), .B1(n_361), .B2(n_499), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_662), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_662), .Y(n_693) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_632), .Y(n_694) );
INVx4_ASAP7_75t_L g695 ( .A(n_633), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_660), .Y(n_696) );
BUFx4_ASAP7_75t_SL g697 ( .A(n_599), .Y(n_697) );
BUFx8_ASAP7_75t_L g698 ( .A(n_612), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_666), .Y(n_699) );
INVx3_ASAP7_75t_L g700 ( .A(n_632), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_631), .A2(n_543), .B(n_548), .C(n_546), .Y(n_701) );
AO22x1_ASAP7_75t_L g702 ( .A1(n_619), .A2(n_426), .B1(n_478), .B2(n_362), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_666), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_617), .Y(n_704) );
BUFx2_ASAP7_75t_SL g705 ( .A(n_646), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_670), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g707 ( .A(n_621), .Y(n_707) );
BUFx3_ASAP7_75t_L g708 ( .A(n_608), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_615), .A2(n_350), .B1(n_402), .B2(n_396), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_626), .A2(n_409), .B1(n_471), .B2(n_422), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_628), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_622), .B(n_426), .Y(n_712) );
INVx5_ASAP7_75t_L g713 ( .A(n_608), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_621), .Y(n_714) );
BUFx3_ASAP7_75t_L g715 ( .A(n_608), .Y(n_715) );
INVx4_ASAP7_75t_L g716 ( .A(n_634), .Y(n_716) );
OAI22xp33_ASAP7_75t_L g717 ( .A1(n_641), .A2(n_414), .B1(n_422), .B2(n_360), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_670), .Y(n_718) );
BUFx2_ASAP7_75t_L g719 ( .A(n_641), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_629), .Y(n_720) );
INVx3_ASAP7_75t_L g721 ( .A(n_608), .Y(n_721) );
OR2x6_ASAP7_75t_L g722 ( .A(n_641), .B(n_381), .Y(n_722) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_630), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_602), .B(n_478), .Y(n_724) );
BUFx6f_ASAP7_75t_L g725 ( .A(n_630), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_639), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_602), .B(n_485), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_631), .B(n_485), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_629), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_643), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_654), .A2(n_424), .B1(n_450), .B2(n_436), .Y(n_731) );
AND2x4_ASAP7_75t_L g732 ( .A(n_609), .B(n_526), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_649), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_624), .B(n_479), .Y(n_734) );
BUFx3_ASAP7_75t_L g735 ( .A(n_630), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_613), .A2(n_414), .B1(n_488), .B2(n_465), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_650), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_604), .A2(n_488), .B1(n_359), .B2(n_363), .Y(n_738) );
BUFx2_ASAP7_75t_L g739 ( .A(n_660), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_605), .B(n_539), .Y(n_740) );
INVx4_ASAP7_75t_L g741 ( .A(n_630), .Y(n_741) );
AND2x4_ASAP7_75t_L g742 ( .A(n_640), .B(n_539), .Y(n_742) );
INVx3_ASAP7_75t_L g743 ( .A(n_636), .Y(n_743) );
AND2x2_ASAP7_75t_SL g744 ( .A(n_600), .B(n_387), .Y(n_744) );
BUFx10_ASAP7_75t_L g745 ( .A(n_676), .Y(n_745) );
INVx2_ASAP7_75t_SL g746 ( .A(n_623), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_636), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_659), .A2(n_597), .B(n_588), .Y(n_748) );
BUFx6f_ASAP7_75t_L g749 ( .A(n_636), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_607), .B(n_546), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_627), .A2(n_355), .B1(n_412), .B2(n_375), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_651), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_671), .Y(n_753) );
BUFx3_ASAP7_75t_L g754 ( .A(n_636), .Y(n_754) );
AND2x4_ASAP7_75t_L g755 ( .A(n_676), .B(n_549), .Y(n_755) );
INVx3_ASAP7_75t_L g756 ( .A(n_623), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_635), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_659), .A2(n_597), .B(n_588), .Y(n_758) );
CKINVDCx5p33_ASAP7_75t_R g759 ( .A(n_667), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_674), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_645), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_627), .A2(n_355), .B1(n_412), .B2(n_375), .Y(n_762) );
OR2x2_ASAP7_75t_L g763 ( .A(n_679), .B(n_385), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_638), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_672), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_645), .Y(n_766) );
CKINVDCx6p67_ASAP7_75t_R g767 ( .A(n_679), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_680), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_679), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_647), .Y(n_770) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_642), .Y(n_771) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_657), .Y(n_772) );
INVx1_ASAP7_75t_SL g773 ( .A(n_673), .Y(n_773) );
INVx2_ASAP7_75t_SL g774 ( .A(n_642), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_680), .Y(n_775) );
INVxp67_ASAP7_75t_L g776 ( .A(n_669), .Y(n_776) );
INVx2_ASAP7_75t_SL g777 ( .A(n_620), .Y(n_777) );
AND2x4_ASAP7_75t_L g778 ( .A(n_676), .B(n_549), .Y(n_778) );
AO22x1_ASAP7_75t_L g779 ( .A1(n_637), .A2(n_420), .B1(n_460), .B2(n_421), .Y(n_779) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_661), .Y(n_780) );
BUFx2_ASAP7_75t_L g781 ( .A(n_664), .Y(n_781) );
NOR2x1_ASAP7_75t_L g782 ( .A(n_653), .B(n_348), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g783 ( .A(n_601), .B(n_575), .Y(n_783) );
NAND2xp5_ASAP7_75t_SL g784 ( .A(n_601), .B(n_575), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_647), .B(n_550), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_603), .B(n_575), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_663), .Y(n_787) );
INVx2_ASAP7_75t_SL g788 ( .A(n_620), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_655), .A2(n_420), .B1(n_460), .B2(n_421), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_656), .B(n_550), .Y(n_790) );
BUFx6f_ASAP7_75t_L g791 ( .A(n_661), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_656), .B(n_486), .Y(n_792) );
AND2x4_ASAP7_75t_L g793 ( .A(n_663), .B(n_551), .Y(n_793) );
AND2x4_ASAP7_75t_L g794 ( .A(n_648), .B(n_551), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_681), .B(n_575), .Y(n_795) );
INVx3_ASAP7_75t_L g796 ( .A(n_682), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_665), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_614), .Y(n_798) );
INVx3_ASAP7_75t_L g799 ( .A(n_682), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_668), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_606), .Y(n_801) );
INVx3_ASAP7_75t_L g802 ( .A(n_678), .Y(n_802) );
INVxp67_ASAP7_75t_L g803 ( .A(n_648), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g804 ( .A1(n_614), .A2(n_588), .B(n_596), .Y(n_804) );
BUFx3_ASAP7_75t_L g805 ( .A(n_678), .Y(n_805) );
BUFx6f_ASAP7_75t_L g806 ( .A(n_677), .Y(n_806) );
BUFx12f_ASAP7_75t_L g807 ( .A(n_610), .Y(n_807) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_722), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_755), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_724), .B(n_434), .Y(n_810) );
BUFx3_ASAP7_75t_L g811 ( .A(n_684), .Y(n_811) );
INVx6_ASAP7_75t_L g812 ( .A(n_684), .Y(n_812) );
INVx2_ASAP7_75t_SL g813 ( .A(n_697), .Y(n_813) );
OA21x2_ASAP7_75t_L g814 ( .A1(n_783), .A2(n_625), .B(n_616), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_770), .B(n_678), .Y(n_815) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_773), .A2(n_372), .B1(n_373), .B2(n_368), .C(n_366), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_755), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_744), .A2(n_616), .B1(n_625), .B2(n_548), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_744), .A2(n_548), .B1(n_388), .B2(n_505), .Y(n_819) );
NOR2xp67_ASAP7_75t_L g820 ( .A(n_731), .B(n_5), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_755), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_781), .A2(n_675), .B1(n_677), .B2(n_393), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_688), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_778), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_722), .A2(n_675), .B1(n_395), .B2(n_398), .Y(n_825) );
BUFx2_ASAP7_75t_L g826 ( .A(n_698), .Y(n_826) );
AOI21xp5_ASAP7_75t_L g827 ( .A1(n_783), .A2(n_588), .B(n_466), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_724), .B(n_388), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_759), .B(n_588), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_727), .B(n_505), .Y(n_830) );
NAND2x1p5_ASAP7_75t_L g831 ( .A(n_716), .B(n_423), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_727), .B(n_374), .Y(n_832) );
INVx2_ASAP7_75t_SL g833 ( .A(n_698), .Y(n_833) );
INVx1_ASAP7_75t_SL g834 ( .A(n_696), .Y(n_834) );
AO31x2_ASAP7_75t_L g835 ( .A1(n_701), .A2(n_524), .A3(n_529), .B(n_521), .Y(n_835) );
AO22x1_ASAP7_75t_SL g836 ( .A1(n_717), .A2(n_408), .B1(n_415), .B2(n_407), .Y(n_836) );
AND2x4_ASAP7_75t_L g837 ( .A(n_716), .B(n_417), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_688), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_757), .B(n_441), .Y(n_839) );
CKINVDCx14_ASAP7_75t_R g840 ( .A(n_714), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g841 ( .A1(n_722), .A2(n_759), .B1(n_714), .B2(n_707), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_722), .A2(n_429), .B1(n_503), .B2(n_413), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_778), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_769), .A2(n_446), .B1(n_459), .B2(n_458), .Y(n_844) );
INVx6_ASAP7_75t_L g845 ( .A(n_698), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_778), .Y(n_846) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_784), .A2(n_596), .B(n_566), .Y(n_847) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_686), .Y(n_848) );
AOI22xp33_ASAP7_75t_SL g849 ( .A1(n_690), .A2(n_498), .B1(n_486), .B2(n_467), .Y(n_849) );
AOI21xp5_ASAP7_75t_R g850 ( .A1(n_732), .A2(n_453), .B(n_5), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_689), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_690), .A2(n_464), .B1(n_475), .B2(n_470), .Y(n_852) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_707), .A2(n_498), .B1(n_503), .B2(n_429), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_689), .Y(n_854) );
NAND2x1p5_ASAP7_75t_L g855 ( .A(n_716), .B(n_423), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_690), .A2(n_497), .B1(n_506), .B2(n_496), .Y(n_856) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_695), .Y(n_857) );
OR2x2_ASAP7_75t_L g858 ( .A(n_736), .B(n_6), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_753), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_760), .A2(n_364), .B1(n_365), .B2(n_354), .Y(n_860) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_695), .Y(n_861) );
AND2x4_ASAP7_75t_L g862 ( .A(n_695), .B(n_371), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_760), .A2(n_379), .B1(n_380), .B2(n_378), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_712), .A2(n_719), .B1(n_732), .B2(n_767), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_793), .Y(n_865) );
INVx4_ASAP7_75t_L g866 ( .A(n_686), .Y(n_866) );
CKINVDCx11_ASAP7_75t_R g867 ( .A(n_807), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_793), .Y(n_868) );
AOI21xp5_ASAP7_75t_L g869 ( .A1(n_784), .A2(n_596), .B(n_566), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_793), .Y(n_870) );
NAND2xp5_ASAP7_75t_SL g871 ( .A(n_686), .B(n_443), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_764), .B(n_392), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_794), .Y(n_873) );
NAND2x1p5_ASAP7_75t_L g874 ( .A(n_796), .B(n_445), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_794), .Y(n_875) );
NAND3x1_ASAP7_75t_L g876 ( .A(n_782), .B(n_403), .C(n_401), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_712), .A2(n_405), .B1(n_419), .B2(n_411), .Y(n_877) );
INVx3_ASAP7_75t_L g878 ( .A(n_686), .Y(n_878) );
AOI21xp33_ASAP7_75t_L g879 ( .A1(n_801), .A2(n_427), .B(n_425), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_732), .A2(n_433), .B1(n_435), .B2(n_432), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_767), .A2(n_447), .B1(n_448), .B2(n_440), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_765), .B(n_451), .Y(n_882) );
INVx1_ASAP7_75t_SL g883 ( .A(n_739), .Y(n_883) );
INVx1_ASAP7_75t_SL g884 ( .A(n_713), .Y(n_884) );
BUFx2_ASAP7_75t_L g885 ( .A(n_687), .Y(n_885) );
O2A1O1Ixp33_ASAP7_75t_SL g886 ( .A1(n_701), .A2(n_455), .B(n_456), .C(n_454), .Y(n_886) );
OAI21x1_ASAP7_75t_L g887 ( .A1(n_804), .A2(n_438), .B(n_431), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_763), .A2(n_462), .B1(n_468), .B2(n_461), .Y(n_888) );
BUFx2_ASAP7_75t_L g889 ( .A(n_687), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_794), .Y(n_890) );
OAI211xp5_ASAP7_75t_L g891 ( .A1(n_710), .A2(n_437), .B(n_442), .C(n_399), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_742), .Y(n_892) );
AND2x4_ASAP7_75t_L g893 ( .A(n_796), .B(n_469), .Y(n_893) );
AO31x2_ASAP7_75t_L g894 ( .A1(n_798), .A2(n_524), .A3(n_529), .B(n_521), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_702), .Y(n_895) );
INVx1_ASAP7_75t_SL g896 ( .A(n_713), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_786), .A2(n_472), .B1(n_476), .B2(n_473), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_786), .A2(n_477), .B1(n_484), .B2(n_483), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_742), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_742), .Y(n_900) );
BUFx2_ASAP7_75t_L g901 ( .A(n_796), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_692), .A2(n_490), .B1(n_491), .B2(n_487), .Y(n_902) );
BUFx6f_ASAP7_75t_L g903 ( .A(n_780), .Y(n_903) );
BUFx3_ASAP7_75t_L g904 ( .A(n_799), .Y(n_904) );
CKINVDCx11_ASAP7_75t_R g905 ( .A(n_807), .Y(n_905) );
AND2x6_ASAP7_75t_L g906 ( .A(n_780), .B(n_438), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_728), .A2(n_492), .B1(n_494), .B2(n_493), .Y(n_907) );
OR2x6_ASAP7_75t_L g908 ( .A(n_705), .B(n_482), .Y(n_908) );
INVx2_ASAP7_75t_L g909 ( .A(n_692), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_740), .Y(n_910) );
AND2x4_ASAP7_75t_L g911 ( .A(n_799), .B(n_500), .Y(n_911) );
OR2x2_ASAP7_75t_L g912 ( .A(n_728), .B(n_6), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_779), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_693), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_799), .Y(n_915) );
HB1xp67_ASAP7_75t_L g916 ( .A(n_683), .Y(n_916) );
NAND2x1p5_ASAP7_75t_L g917 ( .A(n_683), .B(n_445), .Y(n_917) );
OAI211xp5_ASAP7_75t_L g918 ( .A1(n_709), .A2(n_444), .B(n_452), .C(n_501), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_704), .B(n_507), .Y(n_919) );
AND2x4_ASAP7_75t_L g920 ( .A(n_713), .B(n_509), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_738), .A2(n_789), .B1(n_787), .B2(n_745), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_750), .Y(n_922) );
OR2x6_ASAP7_75t_L g923 ( .A(n_694), .B(n_482), .Y(n_923) );
AO31x2_ASAP7_75t_L g924 ( .A1(n_798), .A2(n_529), .A3(n_524), .B(n_540), .Y(n_924) );
CKINVDCx20_ASAP7_75t_R g925 ( .A(n_751), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_776), .B(n_510), .Y(n_926) );
CKINVDCx20_ASAP7_75t_R g927 ( .A(n_762), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_693), .Y(n_928) );
AO31x2_ASAP7_75t_L g929 ( .A1(n_699), .A2(n_540), .A3(n_511), .B(n_463), .Y(n_929) );
BUFx3_ASAP7_75t_L g930 ( .A(n_805), .Y(n_930) );
NOR2xp67_ASAP7_75t_SL g931 ( .A(n_713), .B(n_541), .Y(n_931) );
OAI21x1_ASAP7_75t_L g932 ( .A1(n_748), .A2(n_566), .B(n_562), .Y(n_932) );
A2O1A1Ixp33_ASAP7_75t_L g933 ( .A1(n_750), .A2(n_404), .B(n_534), .C(n_514), .Y(n_933) );
AOI21xp5_ASAP7_75t_L g934 ( .A1(n_758), .A2(n_581), .B(n_562), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_699), .A2(n_541), .B1(n_544), .B2(n_537), .Y(n_935) );
AND2x4_ASAP7_75t_L g936 ( .A(n_713), .B(n_7), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_785), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_703), .A2(n_541), .B1(n_544), .B2(n_537), .Y(n_938) );
BUFx2_ASAP7_75t_R g939 ( .A(n_805), .Y(n_939) );
OAI22xp33_ASAP7_75t_L g940 ( .A1(n_734), .A2(n_537), .B1(n_544), .B2(n_541), .Y(n_940) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_703), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_790), .A2(n_537), .B1(n_544), .B2(n_541), .Y(n_942) );
AND2x4_ASAP7_75t_L g943 ( .A(n_785), .B(n_7), .Y(n_943) );
CKINVDCx20_ASAP7_75t_R g944 ( .A(n_772), .Y(n_944) );
AOI221xp5_ASAP7_75t_L g945 ( .A1(n_691), .A2(n_537), .B1(n_541), .B2(n_544), .C(n_514), .Y(n_945) );
AOI221xp5_ASAP7_75t_L g946 ( .A1(n_819), .A2(n_790), .B1(n_685), .B2(n_792), .C(n_711), .Y(n_946) );
OA21x2_ASAP7_75t_L g947 ( .A1(n_887), .A2(n_718), .B(n_706), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_943), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g949 ( .A1(n_879), .A2(n_800), .B(n_797), .Y(n_949) );
AOI22xp33_ASAP7_75t_SL g950 ( .A1(n_819), .A2(n_803), .B1(n_706), .B2(n_718), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_943), .A2(n_795), .B1(n_726), .B2(n_733), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_859), .Y(n_952) );
INVx4_ASAP7_75t_L g953 ( .A(n_845), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_912), .Y(n_954) );
BUFx3_ASAP7_75t_L g955 ( .A(n_845), .Y(n_955) );
AOI22xp33_ASAP7_75t_SL g956 ( .A1(n_925), .A2(n_795), .B1(n_791), .B2(n_780), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_910), .Y(n_957) );
OAI22xp33_ASAP7_75t_L g958 ( .A1(n_820), .A2(n_927), .B1(n_841), .B2(n_858), .Y(n_958) );
OAI21x1_ASAP7_75t_L g959 ( .A1(n_932), .A2(n_775), .B(n_768), .Y(n_959) );
AOI221xp5_ASAP7_75t_L g960 ( .A1(n_816), .A2(n_730), .B1(n_752), .B2(n_737), .C(n_802), .Y(n_960) );
OAI211xp5_ASAP7_75t_SL g961 ( .A1(n_852), .A2(n_534), .B(n_514), .C(n_802), .Y(n_961) );
BUFx6f_ASAP7_75t_L g962 ( .A(n_848), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_922), .A2(n_756), .B1(n_802), .B2(n_774), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_941), .Y(n_964) );
AOI221xp5_ASAP7_75t_L g965 ( .A1(n_832), .A2(n_729), .B1(n_720), .B2(n_788), .C(n_777), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_842), .A2(n_756), .B1(n_774), .B2(n_746), .Y(n_966) );
AND2x2_ASAP7_75t_L g967 ( .A(n_810), .B(n_720), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_839), .Y(n_968) );
BUFx6f_ASAP7_75t_L g969 ( .A(n_848), .Y(n_969) );
AOI21xp33_ASAP7_75t_L g970 ( .A1(n_818), .A2(n_747), .B(n_746), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_839), .Y(n_971) );
OAI221xp5_ASAP7_75t_L g972 ( .A1(n_856), .A2(n_788), .B1(n_777), .B2(n_756), .C(n_700), .Y(n_972) );
BUFx12f_ASAP7_75t_L g973 ( .A(n_813), .Y(n_973) );
BUFx8_ASAP7_75t_SL g974 ( .A(n_826), .Y(n_974) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_913), .A2(n_806), .B1(n_780), .B2(n_791), .Y(n_975) );
AND2x6_ASAP7_75t_SL g976 ( .A(n_867), .B(n_8), .Y(n_976) );
BUFx3_ASAP7_75t_L g977 ( .A(n_811), .Y(n_977) );
AO21x2_ASAP7_75t_L g978 ( .A1(n_879), .A2(n_747), .B(n_761), .Y(n_978) );
AO31x2_ASAP7_75t_L g979 ( .A1(n_933), .A2(n_775), .A3(n_768), .B(n_761), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_842), .A2(n_771), .B1(n_741), .B2(n_700), .Y(n_980) );
AOI221xp5_ASAP7_75t_L g981 ( .A1(n_828), .A2(n_729), .B1(n_771), .B2(n_741), .C(n_766), .Y(n_981) );
AO21x1_ASAP7_75t_SL g982 ( .A1(n_808), .A2(n_741), .B(n_715), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_895), .A2(n_771), .B1(n_700), .B2(n_754), .Y(n_983) );
AND2x4_ASAP7_75t_L g984 ( .A(n_937), .B(n_694), .Y(n_984) );
OAI21xp5_ASAP7_75t_L g985 ( .A1(n_818), .A2(n_766), .B(n_721), .Y(n_985) );
INVx6_ASAP7_75t_L g986 ( .A(n_866), .Y(n_986) );
A2O1A1Ixp33_ASAP7_75t_L g987 ( .A1(n_829), .A2(n_708), .B(n_715), .C(n_735), .Y(n_987) );
INVx3_ASAP7_75t_L g988 ( .A(n_866), .Y(n_988) );
AND2x4_ASAP7_75t_L g989 ( .A(n_809), .B(n_694), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g990 ( .A1(n_830), .A2(n_771), .B1(n_544), .B2(n_743), .C(n_721), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_850), .A2(n_806), .B1(n_791), .B2(n_723), .Y(n_991) );
OAI22xp33_ASAP7_75t_L g992 ( .A1(n_908), .A2(n_806), .B1(n_791), .B2(n_694), .Y(n_992) );
CKINVDCx5p33_ASAP7_75t_R g993 ( .A(n_905), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_837), .A2(n_754), .B1(n_735), .B2(n_708), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_837), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_823), .Y(n_996) );
AOI22xp33_ASAP7_75t_SL g997 ( .A1(n_840), .A2(n_806), .B1(n_725), .B2(n_749), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g998 ( .A1(n_923), .A2(n_725), .B1(n_749), .B2(n_723), .Y(n_998) );
OR2x2_ASAP7_75t_L g999 ( .A(n_836), .B(n_721), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_923), .A2(n_723), .B1(n_749), .B2(n_725), .Y(n_1000) );
CKINVDCx5p33_ASAP7_75t_R g1001 ( .A(n_812), .Y(n_1001) );
AOI222xp33_ASAP7_75t_L g1002 ( .A1(n_864), .A2(n_743), .B1(n_749), .B2(n_725), .C1(n_723), .C2(n_534), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_883), .B(n_8), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_883), .B(n_9), .Y(n_1004) );
OR2x2_ASAP7_75t_L g1005 ( .A(n_834), .B(n_743), .Y(n_1005) );
AOI21xp5_ASAP7_75t_L g1006 ( .A1(n_934), .A2(n_581), .B(n_562), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_923), .A2(n_544), .B1(n_534), .B2(n_514), .Y(n_1007) );
OA21x2_ASAP7_75t_L g1008 ( .A1(n_847), .A2(n_585), .B(n_581), .Y(n_1008) );
INVx3_ASAP7_75t_L g1009 ( .A(n_936), .Y(n_1009) );
OAI21xp5_ASAP7_75t_L g1010 ( .A1(n_815), .A2(n_534), .B(n_514), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1011 ( .A1(n_872), .A2(n_522), .B1(n_11), .B2(n_9), .Y(n_1011) );
AOI221xp5_ASAP7_75t_L g1012 ( .A1(n_844), .A2(n_522), .B1(n_590), .B2(n_589), .C(n_585), .Y(n_1012) );
INVx2_ASAP7_75t_L g1013 ( .A(n_838), .Y(n_1013) );
OAI211xp5_ASAP7_75t_L g1014 ( .A1(n_918), .A2(n_585), .B(n_590), .C(n_589), .Y(n_1014) );
BUFx4f_ASAP7_75t_SL g1015 ( .A(n_833), .Y(n_1015) );
OAI221xp5_ASAP7_75t_L g1016 ( .A1(n_877), .A2(n_594), .B1(n_590), .B2(n_589), .C(n_583), .Y(n_1016) );
INVx2_ASAP7_75t_L g1017 ( .A(n_851), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g1018 ( .A1(n_888), .A2(n_594), .B1(n_583), .B2(n_569), .C(n_563), .Y(n_1018) );
CKINVDCx5p33_ASAP7_75t_R g1019 ( .A(n_812), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_908), .A2(n_594), .B1(n_563), .B2(n_569), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_908), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_865), .B(n_10), .Y(n_1022) );
INVxp67_ASAP7_75t_L g1023 ( .A(n_834), .Y(n_1023) );
AOI211xp5_ASAP7_75t_L g1024 ( .A1(n_853), .A2(n_563), .B(n_569), .C(n_559), .Y(n_1024) );
AOI221xp5_ASAP7_75t_L g1025 ( .A1(n_907), .A2(n_583), .B1(n_569), .B2(n_563), .C(n_559), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_868), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_825), .B(n_13), .Y(n_1027) );
INVx2_ASAP7_75t_L g1028 ( .A(n_854), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_870), .B(n_13), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_873), .Y(n_1030) );
OAI211xp5_ASAP7_75t_L g1031 ( .A1(n_881), .A2(n_573), .B(n_563), .C(n_569), .Y(n_1031) );
OAI21x1_ASAP7_75t_L g1032 ( .A1(n_869), .A2(n_563), .B(n_559), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_872), .A2(n_16), .B1(n_14), .B2(n_15), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_893), .A2(n_563), .B1(n_569), .B2(n_559), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_875), .Y(n_1035) );
AOI222xp33_ASAP7_75t_SL g1036 ( .A1(n_860), .A2(n_15), .B1(n_17), .B2(n_18), .C1(n_19), .C2(n_20), .Y(n_1036) );
BUFx6f_ASAP7_75t_SL g1037 ( .A(n_893), .Y(n_1037) );
NAND3xp33_ASAP7_75t_L g1038 ( .A(n_945), .B(n_563), .C(n_559), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_831), .A2(n_22), .B1(n_17), .B2(n_21), .Y(n_1039) );
OR2x2_ASAP7_75t_L g1040 ( .A(n_882), .B(n_21), .Y(n_1040) );
HB1xp67_ASAP7_75t_L g1041 ( .A(n_857), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_890), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_892), .B(n_22), .Y(n_1043) );
AOI22xp33_ASAP7_75t_SL g1044 ( .A1(n_885), .A2(n_25), .B1(n_23), .B2(n_24), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_911), .A2(n_569), .B1(n_583), .B2(n_559), .Y(n_1045) );
HB1xp67_ASAP7_75t_L g1046 ( .A(n_861), .Y(n_1046) );
AOI21xp5_ASAP7_75t_L g1047 ( .A1(n_886), .A2(n_569), .B(n_559), .Y(n_1047) );
AOI21xp33_ASAP7_75t_L g1048 ( .A1(n_920), .A2(n_26), .B(n_27), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_882), .Y(n_1049) );
CKINVDCx8_ASAP7_75t_R g1050 ( .A(n_915), .Y(n_1050) );
AO22x2_ASAP7_75t_L g1051 ( .A1(n_936), .A2(n_28), .B1(n_26), .B2(n_27), .Y(n_1051) );
OAI21xp33_ASAP7_75t_SL g1052 ( .A1(n_815), .A2(n_30), .B(n_31), .Y(n_1052) );
BUFx3_ASAP7_75t_L g1053 ( .A(n_904), .Y(n_1053) );
OAI33xp33_ASAP7_75t_L g1054 ( .A1(n_860), .A2(n_31), .A3(n_32), .B1(n_33), .B2(n_34), .B3(n_35), .Y(n_1054) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_926), .A2(n_583), .B1(n_559), .B2(n_36), .C(n_37), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_919), .Y(n_1056) );
OAI221xp5_ASAP7_75t_L g1057 ( .A1(n_921), .A2(n_34), .B1(n_35), .B2(n_36), .C(n_37), .Y(n_1057) );
AOI221xp5_ASAP7_75t_L g1058 ( .A1(n_863), .A2(n_583), .B1(n_40), .B2(n_41), .C(n_42), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_911), .A2(n_583), .B1(n_573), .B2(n_41), .Y(n_1059) );
INVxp67_ASAP7_75t_L g1060 ( .A(n_862), .Y(n_1060) );
INVx2_ASAP7_75t_L g1061 ( .A(n_909), .Y(n_1061) );
OAI211xp5_ASAP7_75t_L g1062 ( .A1(n_891), .A2(n_573), .B(n_583), .C(n_43), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_849), .B(n_39), .Y(n_1063) );
AO31x2_ASAP7_75t_L g1064 ( .A1(n_935), .A2(n_39), .A3(n_40), .B(n_43), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_862), .A2(n_573), .B1(n_45), .B2(n_46), .Y(n_1065) );
OAI21x1_ASAP7_75t_L g1066 ( .A1(n_814), .A2(n_118), .B(n_116), .Y(n_1066) );
INVx11_ASAP7_75t_L g1067 ( .A(n_906), .Y(n_1067) );
AO21x2_ASAP7_75t_L g1068 ( .A1(n_940), .A2(n_120), .B(n_119), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_919), .Y(n_1069) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_831), .A2(n_44), .B1(n_45), .B2(n_46), .Y(n_1070) );
OAI211xp5_ASAP7_75t_L g1071 ( .A1(n_897), .A2(n_573), .B(n_47), .C(n_48), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_899), .A2(n_573), .B1(n_49), .B2(n_50), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_900), .A2(n_573), .B1(n_49), .B2(n_50), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_889), .B(n_44), .Y(n_1074) );
AOI21xp5_ASAP7_75t_L g1075 ( .A1(n_814), .A2(n_573), .B(n_124), .Y(n_1075) );
AOI221xp5_ASAP7_75t_L g1076 ( .A1(n_863), .A2(n_898), .B1(n_902), .B2(n_880), .C(n_822), .Y(n_1076) );
AND2x2_ASAP7_75t_SL g1077 ( .A(n_920), .B(n_51), .Y(n_1077) );
OAI22xp33_ASAP7_75t_L g1078 ( .A1(n_916), .A2(n_51), .B1(n_53), .B2(n_54), .Y(n_1078) );
AOI222xp33_ASAP7_75t_L g1079 ( .A1(n_817), .A2(n_54), .B1(n_55), .B2(n_57), .C1(n_58), .C2(n_59), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_901), .Y(n_1080) );
OAI22xp33_ASAP7_75t_L g1081 ( .A1(n_855), .A2(n_55), .B1(n_57), .B2(n_58), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_952), .Y(n_1082) );
AO21x2_ASAP7_75t_L g1083 ( .A1(n_970), .A2(n_938), .B(n_935), .Y(n_1083) );
OAI211xp5_ASAP7_75t_L g1084 ( .A1(n_1079), .A2(n_871), .B(n_944), .C(n_902), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_958), .A2(n_821), .B1(n_824), .B2(n_843), .Y(n_1085) );
AOI221xp5_ASAP7_75t_L g1086 ( .A1(n_954), .A2(n_846), .B1(n_942), .B2(n_827), .C(n_938), .Y(n_1086) );
OAI21x1_ASAP7_75t_L g1087 ( .A1(n_1032), .A2(n_855), .B(n_878), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_968), .B(n_876), .Y(n_1088) );
OR2x2_ASAP7_75t_L g1089 ( .A(n_964), .B(n_917), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1077), .B(n_874), .Y(n_1090) );
INVx2_ASAP7_75t_L g1091 ( .A(n_996), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_971), .B(n_930), .Y(n_1092) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_1023), .B(n_917), .Y(n_1093) );
NOR2xp33_ASAP7_75t_L g1094 ( .A(n_1049), .B(n_939), .Y(n_1094) );
INVx3_ASAP7_75t_L g1095 ( .A(n_1067), .Y(n_1095) );
AOI22xp5_ASAP7_75t_L g1096 ( .A1(n_1076), .A2(n_884), .B1(n_896), .B2(n_906), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1097 ( .A1(n_951), .A2(n_939), .B1(n_884), .B2(n_896), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1013), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_967), .B(n_914), .Y(n_1099) );
OAI22xp5_ASAP7_75t_SL g1100 ( .A1(n_1015), .A2(n_848), .B1(n_878), .B2(n_928), .Y(n_1100) );
INVxp33_ASAP7_75t_L g1101 ( .A(n_1041), .Y(n_1101) );
OAI221xp5_ASAP7_75t_L g1102 ( .A1(n_1060), .A2(n_903), .B1(n_931), .B2(n_929), .C(n_835), .Y(n_1102) );
OAI211xp5_ASAP7_75t_SL g1103 ( .A1(n_1079), .A2(n_929), .B(n_60), .C(n_61), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_957), .Y(n_1104) );
INVx2_ASAP7_75t_L g1105 ( .A(n_1017), .Y(n_1105) );
OAI22xp5_ASAP7_75t_L g1106 ( .A1(n_948), .A2(n_903), .B1(n_906), .B2(n_929), .Y(n_1106) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1028), .Y(n_1107) );
OAI21xp5_ASAP7_75t_L g1108 ( .A1(n_949), .A2(n_906), .B(n_835), .Y(n_1108) );
NOR2xp33_ASAP7_75t_L g1109 ( .A(n_1056), .B(n_903), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1051), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1003), .B(n_59), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_1057), .A2(n_835), .B1(n_924), .B2(n_894), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_1057), .A2(n_924), .B1(n_894), .B2(n_63), .Y(n_1113) );
OA21x2_ASAP7_75t_L g1114 ( .A1(n_985), .A2(n_894), .B(n_924), .Y(n_1114) );
OA21x2_ASAP7_75t_L g1115 ( .A1(n_985), .A2(n_125), .B(n_121), .Y(n_1115) );
NOR2xp33_ASAP7_75t_R g1116 ( .A(n_1001), .B(n_61), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_1069), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_1117) );
OAI21xp5_ASAP7_75t_L g1118 ( .A1(n_949), .A2(n_66), .B(n_68), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1051), .Y(n_1119) );
INVx3_ASAP7_75t_L g1120 ( .A(n_986), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1061), .Y(n_1121) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_984), .B(n_69), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1051), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1026), .Y(n_1124) );
BUFx2_ASAP7_75t_L g1125 ( .A(n_974), .Y(n_1125) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1030), .Y(n_1126) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1035), .Y(n_1127) );
OR2x2_ASAP7_75t_L g1128 ( .A(n_1046), .B(n_69), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1027), .B(n_70), .Y(n_1129) );
OAI221xp5_ASAP7_75t_SL g1130 ( .A1(n_1052), .A2(n_71), .B1(n_72), .B2(n_73), .C(n_76), .Y(n_1130) );
AOI33xp33_ASAP7_75t_L g1131 ( .A1(n_1044), .A2(n_72), .A3(n_76), .B1(n_77), .B2(n_78), .B3(n_79), .Y(n_1131) );
INVx2_ASAP7_75t_SL g1132 ( .A(n_977), .Y(n_1132) );
NOR2xp33_ASAP7_75t_L g1133 ( .A(n_995), .B(n_77), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1042), .Y(n_1134) );
AND2x4_ASAP7_75t_SL g1135 ( .A(n_953), .B(n_79), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_946), .B(n_80), .Y(n_1136) );
OR2x2_ASAP7_75t_L g1137 ( .A(n_1040), .B(n_82), .Y(n_1137) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_984), .B(n_83), .Y(n_1138) );
AOI222xp33_ASAP7_75t_L g1139 ( .A1(n_1037), .A2(n_84), .B1(n_85), .B2(n_86), .C1(n_87), .C2(n_88), .Y(n_1139) );
NAND2xp5_ASAP7_75t_SL g1140 ( .A(n_991), .B(n_85), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g1141 ( .A1(n_1033), .A2(n_86), .B1(n_88), .B2(n_89), .C(n_90), .Y(n_1141) );
AOI221xp5_ASAP7_75t_L g1142 ( .A1(n_1033), .A2(n_91), .B1(n_92), .B2(n_93), .C(n_94), .Y(n_1142) );
AOI22xp5_ASAP7_75t_L g1143 ( .A1(n_1036), .A2(n_91), .B1(n_93), .B2(n_94), .Y(n_1143) );
NAND4xp25_ASAP7_75t_L g1144 ( .A(n_1063), .B(n_95), .C(n_96), .D(n_97), .Y(n_1144) );
HB1xp67_ASAP7_75t_L g1145 ( .A(n_998), .Y(n_1145) );
INVx2_ASAP7_75t_L g1146 ( .A(n_1043), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1021), .B(n_96), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1022), .Y(n_1148) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1043), .Y(n_1149) );
INVx1_ASAP7_75t_SL g1150 ( .A(n_1019), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_1054), .A2(n_99), .B1(n_102), .B2(n_103), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_1011), .A2(n_103), .B1(n_104), .B2(n_126), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_999), .B(n_104), .Y(n_1153) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_1004), .B(n_130), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_960), .B(n_341), .Y(n_1155) );
OAI221xp5_ASAP7_75t_SL g1156 ( .A1(n_1065), .A2(n_132), .B1(n_133), .B2(n_134), .C(n_137), .Y(n_1156) );
AOI21xp33_ASAP7_75t_L g1157 ( .A1(n_991), .A2(n_138), .B(n_139), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1080), .B(n_141), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_1011), .A2(n_142), .B1(n_143), .B2(n_145), .Y(n_1159) );
OAI221xp5_ASAP7_75t_L g1160 ( .A1(n_950), .A2(n_146), .B1(n_149), .B2(n_151), .C(n_152), .Y(n_1160) );
AOI21xp33_ASAP7_75t_L g1161 ( .A1(n_1062), .A2(n_153), .B(n_154), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1074), .B(n_155), .Y(n_1162) );
OAI21xp5_ASAP7_75t_L g1163 ( .A1(n_1071), .A2(n_156), .B(n_157), .Y(n_1163) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_1009), .A2(n_159), .B1(n_163), .B2(n_165), .Y(n_1164) );
OA21x2_ASAP7_75t_L g1165 ( .A1(n_970), .A2(n_168), .B(n_169), .Y(n_1165) );
BUFx3_ASAP7_75t_L g1166 ( .A(n_986), .Y(n_1166) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1005), .Y(n_1167) );
AOI22xp33_ASAP7_75t_SL g1168 ( .A1(n_1037), .A2(n_170), .B1(n_175), .B2(n_179), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1169 ( .A(n_998), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1053), .B(n_181), .Y(n_1170) );
INVx1_ASAP7_75t_SL g1171 ( .A(n_955), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1050), .B(n_183), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_1058), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_1173) );
OAI211xp5_ASAP7_75t_L g1174 ( .A1(n_1048), .A2(n_190), .B(n_191), .C(n_194), .Y(n_1174) );
INVxp33_ASAP7_75t_SL g1175 ( .A(n_993), .Y(n_1175) );
INVxp67_ASAP7_75t_L g1176 ( .A(n_982), .Y(n_1176) );
OR2x6_ASAP7_75t_L g1177 ( .A(n_1009), .B(n_196), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1022), .B(n_197), .Y(n_1178) );
OAI22xp5_ASAP7_75t_L g1179 ( .A1(n_956), .A2(n_199), .B1(n_200), .B2(n_203), .Y(n_1179) );
AOI22xp5_ASAP7_75t_L g1180 ( .A1(n_1036), .A2(n_204), .B1(n_206), .B2(n_209), .Y(n_1180) );
OAI221xp5_ASAP7_75t_L g1181 ( .A1(n_1055), .A2(n_210), .B1(n_213), .B2(n_214), .C(n_219), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_1078), .A2(n_224), .B1(n_227), .B2(n_231), .Y(n_1182) );
OAI332xp33_ASAP7_75t_L g1183 ( .A1(n_1039), .A2(n_232), .A3(n_234), .B1(n_236), .B2(n_237), .B3(n_238), .C1(n_239), .C2(n_241), .Y(n_1183) );
NAND3xp33_ASAP7_75t_L g1184 ( .A(n_1048), .B(n_242), .C(n_245), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_965), .A2(n_246), .B1(n_247), .B2(n_249), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_1039), .A2(n_251), .B1(n_254), .B2(n_259), .Y(n_1186) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1029), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_972), .B(n_263), .Y(n_1188) );
OAI221xp5_ASAP7_75t_L g1189 ( .A1(n_966), .A2(n_265), .B1(n_268), .B2(n_271), .C(n_272), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_1070), .A2(n_274), .B1(n_276), .B2(n_277), .Y(n_1190) );
AOI221xp5_ASAP7_75t_L g1191 ( .A1(n_1081), .A2(n_280), .B1(n_281), .B2(n_284), .C(n_285), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_1070), .A2(n_286), .B1(n_287), .B2(n_288), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_1029), .A2(n_289), .B1(n_290), .B2(n_291), .Y(n_1193) );
NOR2xp33_ASAP7_75t_L g1194 ( .A(n_961), .B(n_293), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1082), .Y(n_1195) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1114), .Y(n_1196) );
HB1xp67_ASAP7_75t_L g1197 ( .A(n_1145), .Y(n_1197) );
INVx2_ASAP7_75t_L g1198 ( .A(n_1114), .Y(n_1198) );
OR2x2_ASAP7_75t_L g1199 ( .A(n_1167), .B(n_1064), .Y(n_1199) );
AND2x4_ASAP7_75t_L g1200 ( .A(n_1176), .B(n_988), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1099), .B(n_988), .Y(n_1201) );
INVx2_ASAP7_75t_L g1202 ( .A(n_1114), .Y(n_1202) );
OR2x2_ASAP7_75t_SL g1203 ( .A(n_1128), .B(n_976), .Y(n_1203) );
AND2x4_ASAP7_75t_L g1204 ( .A(n_1110), .B(n_962), .Y(n_1204) );
OA211x2_ASAP7_75t_L g1205 ( .A1(n_1140), .A2(n_980), .B(n_981), .C(n_1020), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1206 ( .A(n_1101), .B(n_1064), .Y(n_1206) );
INVx2_ASAP7_75t_SL g1207 ( .A(n_1132), .Y(n_1207) );
AND2x4_ASAP7_75t_L g1208 ( .A(n_1119), .B(n_1064), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1111), .B(n_1101), .Y(n_1209) );
OAI21xp5_ASAP7_75t_L g1210 ( .A1(n_1118), .A2(n_1073), .B(n_1072), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1104), .B(n_989), .Y(n_1211) );
BUFx5_ASAP7_75t_L g1212 ( .A(n_1166), .Y(n_1212) );
NAND2xp5_ASAP7_75t_SL g1213 ( .A(n_1140), .B(n_1106), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1124), .Y(n_1214) );
OAI31xp33_ASAP7_75t_L g1215 ( .A1(n_1084), .A2(n_992), .A3(n_1007), .B(n_1031), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1134), .Y(n_1216) );
OAI33xp33_ASAP7_75t_L g1217 ( .A1(n_1144), .A2(n_1007), .A3(n_975), .B1(n_1000), .B2(n_1038), .B3(n_1059), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1126), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1127), .Y(n_1219) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1091), .Y(n_1220) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_1085), .A2(n_1024), .B1(n_997), .B2(n_994), .Y(n_1221) );
INVx2_ASAP7_75t_L g1222 ( .A(n_1098), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1090), .B(n_989), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1224 ( .A(n_1089), .B(n_1000), .Y(n_1224) );
OAI21xp5_ASAP7_75t_SL g1225 ( .A1(n_1139), .A2(n_1002), .B(n_990), .Y(n_1225) );
NOR2xp33_ASAP7_75t_L g1226 ( .A(n_1088), .B(n_973), .Y(n_1226) );
OAI22xp5_ASAP7_75t_L g1227 ( .A1(n_1085), .A2(n_963), .B1(n_986), .B2(n_983), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1105), .Y(n_1228) );
AOI33xp33_ASAP7_75t_L g1229 ( .A1(n_1143), .A2(n_1045), .A3(n_1034), .B1(n_1012), .B2(n_1025), .B3(n_1002), .Y(n_1229) );
AOI22xp5_ASAP7_75t_L g1230 ( .A1(n_1094), .A2(n_1014), .B1(n_978), .B2(n_1068), .Y(n_1230) );
AOI211xp5_ASAP7_75t_L g1231 ( .A1(n_1116), .A2(n_1010), .B(n_987), .C(n_1075), .Y(n_1231) );
NOR3xp33_ASAP7_75t_L g1232 ( .A(n_1103), .B(n_1130), .C(n_1183), .Y(n_1232) );
BUFx2_ASAP7_75t_L g1233 ( .A(n_1166), .Y(n_1233) );
INVx2_ASAP7_75t_SL g1234 ( .A(n_1125), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1122), .B(n_979), .Y(n_1235) );
NAND4xp25_ASAP7_75t_L g1236 ( .A(n_1153), .B(n_1006), .C(n_1047), .D(n_1018), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1107), .Y(n_1237) );
OAI321xp33_ASAP7_75t_L g1238 ( .A1(n_1180), .A2(n_1016), .A3(n_969), .B1(n_962), .B2(n_1068), .C(n_298), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_1123), .B(n_978), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1121), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1092), .Y(n_1241) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1146), .Y(n_1242) );
INVxp67_ASAP7_75t_L g1243 ( .A(n_1102), .Y(n_1243) );
NAND2x1p5_ASAP7_75t_L g1244 ( .A(n_1095), .B(n_969), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1138), .Y(n_1245) );
AOI221xp5_ASAP7_75t_L g1246 ( .A1(n_1133), .A2(n_969), .B1(n_962), .B2(n_979), .C(n_1008), .Y(n_1246) );
INVx2_ASAP7_75t_L g1247 ( .A(n_1149), .Y(n_1247) );
NOR3xp33_ASAP7_75t_L g1248 ( .A(n_1136), .B(n_1066), .C(n_959), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1109), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1109), .Y(n_1250) );
OAI21x1_ASAP7_75t_L g1251 ( .A1(n_1087), .A2(n_1008), .B(n_947), .Y(n_1251) );
AOI22xp5_ASAP7_75t_L g1252 ( .A1(n_1094), .A2(n_947), .B1(n_979), .B2(n_296), .Y(n_1252) );
AOI21xp33_ASAP7_75t_L g1253 ( .A1(n_1097), .A2(n_294), .B(n_295), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1148), .B(n_340), .Y(n_1254) );
INVx2_ASAP7_75t_L g1255 ( .A(n_1187), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1116), .B(n_297), .Y(n_1256) );
AND2x4_ASAP7_75t_L g1257 ( .A(n_1145), .B(n_300), .Y(n_1257) );
INVx5_ASAP7_75t_SL g1258 ( .A(n_1177), .Y(n_1258) );
OAI222xp33_ASAP7_75t_L g1259 ( .A1(n_1177), .A2(n_301), .B1(n_302), .B2(n_303), .C1(n_304), .C2(n_306), .Y(n_1259) );
HB1xp67_ASAP7_75t_L g1260 ( .A(n_1169), .Y(n_1260) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1093), .Y(n_1261) );
INVxp67_ASAP7_75t_SL g1262 ( .A(n_1169), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1137), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1147), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1133), .B(n_308), .Y(n_1265) );
AOI33xp33_ASAP7_75t_L g1266 ( .A1(n_1117), .A2(n_310), .A3(n_313), .B1(n_314), .B2(n_315), .B3(n_318), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1131), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1162), .B(n_319), .Y(n_1268) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1083), .Y(n_1269) );
AO22x1_ASAP7_75t_L g1270 ( .A1(n_1175), .A2(n_320), .B1(n_321), .B2(n_323), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1135), .B(n_325), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1170), .B(n_326), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1172), .B(n_328), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1131), .Y(n_1274) );
INVx2_ASAP7_75t_L g1275 ( .A(n_1083), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1120), .B(n_329), .Y(n_1276) );
OAI33xp33_ASAP7_75t_L g1277 ( .A1(n_1129), .A2(n_336), .A3(n_337), .B1(n_338), .B2(n_1154), .B3(n_1158), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1278 ( .A(n_1171), .B(n_1150), .Y(n_1278) );
INVx2_ASAP7_75t_L g1279 ( .A(n_1115), .Y(n_1279) );
INVx2_ASAP7_75t_L g1280 ( .A(n_1115), .Y(n_1280) );
BUFx3_ASAP7_75t_L g1281 ( .A(n_1120), .Y(n_1281) );
AOI21xp5_ASAP7_75t_SL g1282 ( .A1(n_1177), .A2(n_1115), .B(n_1179), .Y(n_1282) );
OAI31xp33_ASAP7_75t_L g1283 ( .A1(n_1188), .A2(n_1156), .A3(n_1174), .B(n_1152), .Y(n_1283) );
INVxp67_ASAP7_75t_L g1284 ( .A(n_1108), .Y(n_1284) );
INVx2_ASAP7_75t_L g1285 ( .A(n_1165), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1195), .Y(n_1286) );
NOR3xp33_ASAP7_75t_SL g1287 ( .A(n_1225), .B(n_1141), .C(n_1142), .Y(n_1287) );
BUFx3_ASAP7_75t_L g1288 ( .A(n_1200), .Y(n_1288) );
OAI31xp33_ASAP7_75t_L g1289 ( .A1(n_1267), .A2(n_1100), .A3(n_1117), .B(n_1160), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1209), .B(n_1096), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_1261), .B(n_1152), .Y(n_1291) );
NAND3xp33_ASAP7_75t_L g1292 ( .A(n_1243), .B(n_1151), .C(n_1186), .Y(n_1292) );
HB1xp67_ASAP7_75t_L g1293 ( .A(n_1197), .Y(n_1293) );
NOR2x1_ASAP7_75t_L g1294 ( .A(n_1200), .B(n_1184), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1201), .B(n_1112), .Y(n_1295) );
BUFx3_ASAP7_75t_L g1296 ( .A(n_1200), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_1218), .B(n_1113), .Y(n_1297) );
OR2x2_ASAP7_75t_L g1298 ( .A(n_1219), .B(n_1113), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1214), .Y(n_1299) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_1263), .B(n_1112), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1208), .B(n_1151), .Y(n_1301) );
INVx1_ASAP7_75t_SL g1302 ( .A(n_1207), .Y(n_1302) );
AND2x4_ASAP7_75t_L g1303 ( .A(n_1208), .B(n_1163), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1223), .B(n_1190), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1241), .B(n_1086), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1216), .B(n_1155), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1249), .B(n_1178), .Y(n_1307) );
INVx1_ASAP7_75t_SL g1308 ( .A(n_1278), .Y(n_1308) );
INVx2_ASAP7_75t_L g1309 ( .A(n_1196), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1242), .Y(n_1310) );
OAI22xp5_ASAP7_75t_L g1311 ( .A1(n_1258), .A2(n_1186), .B1(n_1190), .B2(n_1192), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1247), .Y(n_1312) );
NAND2x1_ASAP7_75t_L g1313 ( .A(n_1282), .B(n_1165), .Y(n_1313) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1196), .Y(n_1314) );
OAI31xp33_ASAP7_75t_L g1315 ( .A1(n_1274), .A2(n_1181), .A3(n_1189), .B(n_1164), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1255), .Y(n_1316) );
NOR2xp33_ASAP7_75t_L g1317 ( .A(n_1264), .B(n_1194), .Y(n_1317) );
NAND2xp33_ASAP7_75t_L g1318 ( .A(n_1232), .B(n_1159), .Y(n_1318) );
INVx2_ASAP7_75t_L g1319 ( .A(n_1198), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1255), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1250), .B(n_1182), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1228), .Y(n_1322) );
AND2x2_ASAP7_75t_SL g1323 ( .A(n_1257), .B(n_1193), .Y(n_1323) );
AOI31xp67_ASAP7_75t_SL g1324 ( .A1(n_1258), .A2(n_1168), .A3(n_1157), .B(n_1185), .Y(n_1324) );
OAI322xp33_ASAP7_75t_L g1325 ( .A1(n_1206), .A2(n_1194), .A3(n_1173), .B1(n_1191), .B2(n_1185), .C1(n_1193), .C2(n_1161), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1237), .B(n_1173), .Y(n_1326) );
NAND4xp25_ASAP7_75t_SL g1327 ( .A(n_1256), .B(n_1232), .C(n_1271), .D(n_1266), .Y(n_1327) );
NOR2x1_ASAP7_75t_L g1328 ( .A(n_1259), .B(n_1233), .Y(n_1328) );
AND2x2_ASAP7_75t_SL g1329 ( .A(n_1257), .B(n_1235), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1240), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1245), .B(n_1220), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1211), .B(n_1220), .Y(n_1332) );
NOR2xp33_ASAP7_75t_L g1333 ( .A(n_1217), .B(n_1203), .Y(n_1333) );
AND2x4_ASAP7_75t_L g1334 ( .A(n_1208), .B(n_1204), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1222), .Y(n_1335) );
AOI21xp33_ASAP7_75t_L g1336 ( .A1(n_1243), .A2(n_1284), .B(n_1283), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1284), .B(n_1198), .Y(n_1337) );
OAI22xp33_ASAP7_75t_L g1338 ( .A1(n_1221), .A2(n_1224), .B1(n_1227), .B2(n_1210), .Y(n_1338) );
AND3x1_ASAP7_75t_L g1339 ( .A(n_1234), .B(n_1226), .C(n_1273), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1222), .B(n_1281), .Y(n_1340) );
OAI22xp5_ASAP7_75t_L g1341 ( .A1(n_1257), .A2(n_1231), .B1(n_1205), .B2(n_1268), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1281), .B(n_1226), .Y(n_1342) );
NAND2xp5_ASAP7_75t_SL g1343 ( .A(n_1246), .B(n_1212), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1344 ( .A(n_1199), .B(n_1197), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1260), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1260), .B(n_1262), .Y(n_1346) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1202), .Y(n_1347) );
INVx2_ASAP7_75t_SL g1348 ( .A(n_1212), .Y(n_1348) );
OAI221xp5_ASAP7_75t_L g1349 ( .A1(n_1215), .A2(n_1230), .B1(n_1252), .B2(n_1213), .C(n_1253), .Y(n_1349) );
INVx1_ASAP7_75t_SL g1350 ( .A(n_1244), .Y(n_1350) );
INVxp67_ASAP7_75t_SL g1351 ( .A(n_1202), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1337), .B(n_1262), .Y(n_1352) );
AND2x4_ASAP7_75t_SL g1353 ( .A(n_1342), .B(n_1204), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1286), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1290), .B(n_1239), .Y(n_1355) );
OAI211xp5_ASAP7_75t_L g1356 ( .A1(n_1333), .A2(n_1213), .B(n_1272), .C(n_1265), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1337), .B(n_1275), .Y(n_1357) );
NOR2xp33_ASAP7_75t_L g1358 ( .A(n_1302), .B(n_1308), .Y(n_1358) );
INVx1_ASAP7_75t_SL g1359 ( .A(n_1339), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1331), .B(n_1212), .Y(n_1360) );
OR2x2_ASAP7_75t_L g1361 ( .A(n_1344), .B(n_1275), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1335), .Y(n_1362) );
NAND2xp5_ASAP7_75t_SL g1363 ( .A(n_1328), .B(n_1212), .Y(n_1363) );
XNOR2x1_ASAP7_75t_L g1364 ( .A(n_1338), .B(n_1270), .Y(n_1364) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1300), .B(n_1212), .Y(n_1365) );
OAI21xp5_ASAP7_75t_L g1366 ( .A1(n_1333), .A2(n_1266), .B(n_1238), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1334), .B(n_1269), .Y(n_1367) );
NOR2xp33_ASAP7_75t_L g1368 ( .A(n_1336), .B(n_1244), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1334), .B(n_1269), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1299), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1334), .B(n_1280), .Y(n_1371) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1346), .B(n_1280), .Y(n_1372) );
INVx1_ASAP7_75t_SL g1373 ( .A(n_1340), .Y(n_1373) );
INVx1_ASAP7_75t_SL g1374 ( .A(n_1350), .Y(n_1374) );
NOR2x1_ASAP7_75t_L g1375 ( .A(n_1294), .B(n_1236), .Y(n_1375) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1309), .Y(n_1376) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1322), .Y(n_1377) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1330), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1301), .B(n_1279), .Y(n_1379) );
INVxp67_ASAP7_75t_SL g1380 ( .A(n_1351), .Y(n_1380) );
AOI21xp5_ASAP7_75t_L g1381 ( .A1(n_1323), .A2(n_1277), .B(n_1217), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1301), .B(n_1279), .Y(n_1382) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1345), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1332), .Y(n_1384) );
INVxp67_ASAP7_75t_L g1385 ( .A(n_1317), .Y(n_1385) );
OAI21xp33_ASAP7_75t_L g1386 ( .A1(n_1338), .A2(n_1254), .B(n_1229), .Y(n_1386) );
INVx1_ASAP7_75t_SL g1387 ( .A(n_1288), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1295), .B(n_1285), .Y(n_1388) );
INVx2_ASAP7_75t_L g1389 ( .A(n_1309), .Y(n_1389) );
CKINVDCx16_ASAP7_75t_R g1390 ( .A(n_1288), .Y(n_1390) );
OR2x2_ASAP7_75t_L g1391 ( .A(n_1293), .B(n_1285), .Y(n_1391) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1310), .Y(n_1392) );
OR2x2_ASAP7_75t_L g1393 ( .A(n_1293), .B(n_1251), .Y(n_1393) );
AOI21xp33_ASAP7_75t_L g1394 ( .A1(n_1341), .A2(n_1276), .B(n_1277), .Y(n_1394) );
INVx2_ASAP7_75t_SL g1395 ( .A(n_1296), .Y(n_1395) );
NOR3xp33_ASAP7_75t_L g1396 ( .A(n_1327), .B(n_1248), .C(n_1229), .Y(n_1396) );
HB1xp67_ASAP7_75t_L g1397 ( .A(n_1312), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1388), .B(n_1351), .Y(n_1398) );
NAND2x1_ASAP7_75t_SL g1399 ( .A(n_1375), .B(n_1303), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1361), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1384), .B(n_1320), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1388), .B(n_1303), .Y(n_1402) );
INVx1_ASAP7_75t_SL g1403 ( .A(n_1387), .Y(n_1403) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1361), .Y(n_1404) );
INVx2_ASAP7_75t_L g1405 ( .A(n_1376), .Y(n_1405) );
NOR2xp33_ASAP7_75t_L g1406 ( .A(n_1359), .B(n_1305), .Y(n_1406) );
XNOR2xp5_ASAP7_75t_L g1407 ( .A(n_1364), .B(n_1329), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g1408 ( .A(n_1385), .B(n_1321), .Y(n_1408) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1397), .Y(n_1409) );
BUFx2_ASAP7_75t_L g1410 ( .A(n_1380), .Y(n_1410) );
HB1xp67_ASAP7_75t_L g1411 ( .A(n_1373), .Y(n_1411) );
INVx2_ASAP7_75t_L g1412 ( .A(n_1389), .Y(n_1412) );
OAI322xp33_ASAP7_75t_L g1413 ( .A1(n_1364), .A2(n_1291), .A3(n_1298), .B1(n_1297), .B2(n_1349), .C1(n_1307), .C2(n_1313), .Y(n_1413) );
INVx2_ASAP7_75t_SL g1414 ( .A(n_1353), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1372), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1379), .B(n_1303), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1372), .Y(n_1417) );
OR2x2_ASAP7_75t_L g1418 ( .A(n_1355), .B(n_1347), .Y(n_1418) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1354), .Y(n_1419) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1383), .B(n_1316), .Y(n_1420) );
XOR2x2_ASAP7_75t_L g1421 ( .A(n_1363), .B(n_1329), .Y(n_1421) );
INVx2_ASAP7_75t_L g1422 ( .A(n_1391), .Y(n_1422) );
INVxp67_ASAP7_75t_L g1423 ( .A(n_1358), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1379), .B(n_1347), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1377), .B(n_1319), .Y(n_1425) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1382), .B(n_1319), .Y(n_1426) );
NOR2xp33_ASAP7_75t_L g1427 ( .A(n_1374), .B(n_1318), .Y(n_1427) );
NOR2xp33_ASAP7_75t_L g1428 ( .A(n_1386), .B(n_1292), .Y(n_1428) );
AOI22xp5_ASAP7_75t_L g1429 ( .A1(n_1396), .A2(n_1323), .B1(n_1311), .B2(n_1287), .Y(n_1429) );
XNOR2x1_ASAP7_75t_L g1430 ( .A(n_1366), .B(n_1304), .Y(n_1430) );
AOI22xp33_ASAP7_75t_L g1431 ( .A1(n_1381), .A2(n_1289), .B1(n_1306), .B2(n_1343), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1370), .Y(n_1432) );
OAI21xp5_ASAP7_75t_L g1433 ( .A1(n_1363), .A2(n_1343), .B(n_1315), .Y(n_1433) );
INVxp67_ASAP7_75t_L g1434 ( .A(n_1393), .Y(n_1434) );
XOR2xp5_ASAP7_75t_L g1435 ( .A(n_1390), .B(n_1296), .Y(n_1435) );
NOR2xp33_ASAP7_75t_L g1436 ( .A(n_1368), .B(n_1325), .Y(n_1436) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1378), .Y(n_1437) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1362), .Y(n_1438) );
INVx2_ASAP7_75t_L g1439 ( .A(n_1357), .Y(n_1439) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1362), .Y(n_1440) );
NOR2xp33_ASAP7_75t_L g1441 ( .A(n_1356), .B(n_1326), .Y(n_1441) );
AOI22xp5_ASAP7_75t_L g1442 ( .A1(n_1365), .A2(n_1348), .B1(n_1324), .B2(n_1314), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1392), .Y(n_1443) );
OAI321xp33_ASAP7_75t_L g1444 ( .A1(n_1433), .A2(n_1429), .A3(n_1442), .B1(n_1428), .B2(n_1436), .C(n_1431), .Y(n_1444) );
INVx1_ASAP7_75t_SL g1445 ( .A(n_1403), .Y(n_1445) );
AOI211xp5_ASAP7_75t_SL g1446 ( .A1(n_1413), .A2(n_1436), .B(n_1441), .C(n_1394), .Y(n_1446) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1409), .Y(n_1447) );
INVx2_ASAP7_75t_L g1448 ( .A(n_1410), .Y(n_1448) );
OAI211xp5_ASAP7_75t_L g1449 ( .A1(n_1431), .A2(n_1399), .B(n_1427), .C(n_1441), .Y(n_1449) );
OAI321xp33_ASAP7_75t_L g1450 ( .A1(n_1414), .A2(n_1434), .A3(n_1406), .B1(n_1423), .B2(n_1410), .C(n_1395), .Y(n_1450) );
OAI21xp5_ASAP7_75t_SL g1451 ( .A1(n_1407), .A2(n_1430), .B(n_1435), .Y(n_1451) );
O2A1O1Ixp33_ASAP7_75t_L g1452 ( .A1(n_1434), .A2(n_1403), .B(n_1411), .C(n_1408), .Y(n_1452) );
AOI221x1_ASAP7_75t_SL g1453 ( .A1(n_1415), .A2(n_1417), .B1(n_1400), .B2(n_1404), .C(n_1409), .Y(n_1453) );
AOI22xp33_ASAP7_75t_SL g1454 ( .A1(n_1414), .A2(n_1353), .B1(n_1421), .B2(n_1398), .Y(n_1454) );
OA22x2_ASAP7_75t_L g1455 ( .A1(n_1421), .A2(n_1400), .B1(n_1437), .B2(n_1432), .Y(n_1455) );
OAI22xp5_ASAP7_75t_L g1456 ( .A1(n_1454), .A2(n_1418), .B1(n_1402), .B2(n_1439), .Y(n_1456) );
A2O1A1Ixp33_ASAP7_75t_L g1457 ( .A1(n_1451), .A2(n_1419), .B(n_1401), .C(n_1416), .Y(n_1457) );
AOI222xp33_ASAP7_75t_L g1458 ( .A1(n_1444), .A2(n_1419), .B1(n_1401), .B2(n_1422), .C1(n_1440), .C2(n_1443), .Y(n_1458) );
AOI21xp5_ASAP7_75t_L g1459 ( .A1(n_1450), .A2(n_1420), .B(n_1425), .Y(n_1459) );
OAI21xp5_ASAP7_75t_SL g1460 ( .A1(n_1446), .A2(n_1367), .B(n_1369), .Y(n_1460) );
NAND5xp2_ASAP7_75t_L g1461 ( .A(n_1449), .B(n_1352), .C(n_1371), .D(n_1382), .E(n_1367), .Y(n_1461) );
AOI211xp5_ASAP7_75t_SL g1462 ( .A1(n_1455), .A2(n_1393), .B(n_1360), .C(n_1369), .Y(n_1462) );
NAND4xp25_ASAP7_75t_L g1463 ( .A(n_1458), .B(n_1453), .C(n_1445), .D(n_1452), .Y(n_1463) );
NAND4xp25_ASAP7_75t_L g1464 ( .A(n_1457), .B(n_1448), .C(n_1447), .D(n_1352), .Y(n_1464) );
NAND4xp25_ASAP7_75t_L g1465 ( .A(n_1457), .B(n_1371), .C(n_1420), .D(n_1425), .Y(n_1465) );
OR2x2_ASAP7_75t_L g1466 ( .A(n_1465), .B(n_1461), .Y(n_1466) );
NOR4xp25_ASAP7_75t_L g1467 ( .A(n_1463), .B(n_1460), .C(n_1456), .D(n_1462), .Y(n_1467) );
AOI21xp33_ASAP7_75t_SL g1468 ( .A1(n_1467), .A2(n_1464), .B(n_1459), .Y(n_1468) );
OAI221xp5_ASAP7_75t_L g1469 ( .A1(n_1468), .A2(n_1466), .B1(n_1348), .B2(n_1422), .C(n_1438), .Y(n_1469) );
INVxp67_ASAP7_75t_L g1470 ( .A(n_1469), .Y(n_1470) );
INVxp67_ASAP7_75t_L g1471 ( .A(n_1470), .Y(n_1471) );
AOI221xp5_ASAP7_75t_L g1472 ( .A1(n_1471), .A2(n_1405), .B1(n_1412), .B2(n_1424), .C(n_1426), .Y(n_1472) );
endmodule