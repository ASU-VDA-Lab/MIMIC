module fake_jpeg_11663_n_136 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_7),
.Y(n_32)
);

NOR2xp67_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_41),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_0),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_39),
.B1(n_42),
.B2(n_38),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_55),
.B1(n_61),
.B2(n_30),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_23),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_19),
.C(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_1),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_15),
.B1(n_22),
.B2(n_27),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_60),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_26),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_28),
.C(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_29),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_27),
.B1(n_22),
.B2(n_26),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_34),
.B1(n_36),
.B2(n_22),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_68),
.B1(n_46),
.B2(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_30),
.B1(n_21),
.B2(n_28),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_40),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_72),
.B(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_25),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_20),
.B1(n_17),
.B2(n_40),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_48),
.C(n_53),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_51),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_87),
.B1(n_90),
.B2(n_63),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_43),
.B1(n_58),
.B2(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_71),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_68),
.C(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_49),
.B1(n_48),
.B2(n_51),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_74),
.Y(n_97)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_56),
.A3(n_53),
.B1(n_6),
.B2(n_3),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_70),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_87),
.B1(n_83),
.B2(n_66),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_103),
.B1(n_81),
.B2(n_85),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_95),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_98),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_104),
.C(n_53),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_77),
.B1(n_64),
.B2(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_13),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_13),
.Y(n_109)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_70),
.B1(n_64),
.B2(n_67),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_113),
.B1(n_103),
.B2(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_94),
.C(n_93),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_116),
.C(n_117),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_96),
.C(n_98),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_100),
.C(n_102),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_86),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_108),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_125),
.C(n_53),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_105),
.B(n_112),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_86),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_12),
.C1(n_76),
.C2(n_5),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_129),
.C(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_121),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_9),
.C(n_10),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_131),
.C(n_12),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);


endmodule