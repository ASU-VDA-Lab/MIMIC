module fake_netlist_5_2378_n_1666 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1666);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1666;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx5_ASAP7_75t_L g151 ( 
.A(n_39),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_27),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_72),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_74),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_60),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_36),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_130),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_67),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_90),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_19),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_107),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_53),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_99),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_7),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_6),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_50),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_68),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_55),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_129),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_89),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_50),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_31),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_113),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_136),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_48),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_111),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_43),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_0),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_86),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_114),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_36),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_106),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_125),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_85),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_128),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_95),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_54),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_135),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_137),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_1),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_134),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_51),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_94),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_126),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_23),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_4),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_22),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_109),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_31),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_96),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_123),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_10),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_147),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_122),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_92),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_145),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_140),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_18),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_62),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_13),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_46),
.Y(n_218)
);

BUFx8_ASAP7_75t_SL g219 ( 
.A(n_93),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_39),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_14),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_102),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_53),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_119),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_118),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_101),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_28),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_48),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_115),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_112),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_3),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_117),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_63),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_24),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_131),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_120),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_139),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_56),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_73),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_10),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_103),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_38),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_17),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_19),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_76),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_49),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_88),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_57),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_23),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_91),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_0),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_22),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_132),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_33),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_110),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_17),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_51),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_14),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_13),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_24),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_49),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_43),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_100),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_64),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_8),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_25),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_16),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_142),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_116),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_35),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_59),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_84),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_28),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_121),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_7),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_69),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_83),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_2),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_105),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_5),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_20),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_47),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_6),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_38),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_124),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_5),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_81),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_9),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_150),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_46),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_8),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_66),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_133),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_54),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_77),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_58),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_45),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_75),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_25),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_11),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_1),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_82),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_40),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_151),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_151),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_151),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_219),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_159),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_151),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_192),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_178),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_151),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_180),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_151),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_186),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_241),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_151),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_194),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_187),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_151),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_189),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_196),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_198),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_262),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_226),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_262),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_253),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_262),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_262),
.B(n_2),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_262),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_220),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_200),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_220),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_220),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_184),
.B(n_3),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_201),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_209),
.B(n_4),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_268),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_220),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_220),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_205),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_234),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_223),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_207),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_238),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_269),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_167),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_273),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_167),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_208),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_211),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_184),
.B(n_9),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_259),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_259),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_193),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_233),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_212),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_281),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_241),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_213),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_179),
.B(n_11),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_281),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_288),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_214),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_222),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_288),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_225),
.B(n_12),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_225),
.B(n_12),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_179),
.Y(n_375)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_152),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_224),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_230),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_152),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_209),
.B(n_15),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_232),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_239),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_228),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_157),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_245),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_228),
.Y(n_386)
);

INVxp33_ASAP7_75t_SL g387 ( 
.A(n_157),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_162),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_247),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_338),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_336),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_320),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_330),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_312),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_352),
.B(n_191),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_339),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_314),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_229),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_316),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_344),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_345),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_R g406 ( 
.A(n_309),
.B(n_248),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_338),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_229),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_305),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_321),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_306),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_374),
.B(n_340),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_332),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_318),
.B(n_154),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_358),
.B(n_154),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_306),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_307),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_304),
.A2(n_275),
.B1(n_243),
.B2(n_258),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_160),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_307),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_365),
.B(n_153),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_310),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_310),
.B(n_160),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_313),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_352),
.B(n_191),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_343),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_313),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_323),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_315),
.B(n_163),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_315),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_319),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_319),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_325),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_326),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_362),
.B(n_191),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_322),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_322),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_361),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_347),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_324),
.Y(n_440)
);

AND2x6_ASAP7_75t_L g441 ( 
.A(n_324),
.B(n_255),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_328),
.B(n_163),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_328),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_365),
.B(n_153),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_337),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_341),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_R g447 ( 
.A(n_308),
.B(n_250),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_329),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_329),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_351),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_331),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_342),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_346),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_331),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_376),
.B(n_155),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_349),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_366),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_L g458 ( 
.A(n_356),
.B(n_168),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_377),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_333),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_375),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_357),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_379),
.B(n_216),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_412),
.B(n_363),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_461),
.B(n_388),
.Y(n_465)
);

AND2x2_ASAP7_75t_SL g466 ( 
.A(n_412),
.B(n_158),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_455),
.B(n_158),
.Y(n_468)
);

AND2x2_ASAP7_75t_SL g469 ( 
.A(n_402),
.B(n_408),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_396),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_455),
.B(n_171),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_452),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_L g473 ( 
.A(n_415),
.B(n_255),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_423),
.B(n_171),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_421),
.B(n_375),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_402),
.B(n_210),
.Y(n_476)
);

NAND3xp33_ASAP7_75t_L g477 ( 
.A(n_415),
.B(n_419),
.C(n_423),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_397),
.B(n_291),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_396),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_402),
.B(n_370),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_421),
.B(n_383),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_457),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_401),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_461),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_421),
.B(n_383),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_414),
.B(n_317),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_429),
.B(n_210),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_401),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_408),
.A2(n_334),
.B1(n_342),
.B2(n_300),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_408),
.A2(n_291),
.B1(n_300),
.B2(n_380),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_419),
.B(n_371),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_429),
.B(n_381),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_442),
.A2(n_311),
.B1(n_348),
.B2(n_387),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_401),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_442),
.B(n_414),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_452),
.B(n_235),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_416),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_390),
.B(n_427),
.Y(n_498)
);

INVx5_ASAP7_75t_L g499 ( 
.A(n_441),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_447),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_439),
.B(n_354),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_394),
.B(n_235),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_399),
.B(n_237),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_427),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_459),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_444),
.B(n_353),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_430),
.A2(n_384),
.B1(n_286),
.B2(n_242),
.Y(n_507)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_439),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_450),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_450),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_392),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_393),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_430),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_425),
.B(n_386),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_438),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_463),
.B(n_385),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_407),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_431),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_407),
.Y(n_519)
);

AND2x2_ASAP7_75t_SL g520 ( 
.A(n_458),
.B(n_237),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_438),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_409),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_403),
.B(n_271),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_443),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_437),
.A2(n_454),
.B1(n_451),
.B2(n_449),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_407),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_410),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_444),
.B(n_386),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_437),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_449),
.B(n_271),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_451),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_454),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_422),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_411),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_422),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_428),
.B(n_255),
.Y(n_537)
);

NAND2x1p5_ASAP7_75t_L g538 ( 
.A(n_444),
.B(n_161),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_422),
.Y(n_539)
);

BUFx8_ASAP7_75t_SL g540 ( 
.A(n_413),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_426),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_433),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_434),
.A2(n_389),
.B1(n_382),
.B2(n_378),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_406),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_438),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_411),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_443),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_462),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_443),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_448),
.B(n_335),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_418),
.B(n_270),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_391),
.B(n_353),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_411),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_391),
.B(n_372),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_448),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_417),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_417),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_417),
.B(n_255),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_420),
.Y(n_559)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_441),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_441),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_418),
.B(n_372),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_445),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_446),
.B(n_350),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_395),
.B(n_369),
.Y(n_565)
);

INVx6_ASAP7_75t_L g566 ( 
.A(n_441),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_441),
.Y(n_567)
);

AND2x6_ASAP7_75t_L g568 ( 
.A(n_424),
.B(n_255),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_424),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_441),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_424),
.B(n_156),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_435),
.B(n_369),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_453),
.A2(n_173),
.B1(n_287),
.B2(n_289),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_432),
.B(n_165),
.Y(n_574)
);

AO21x2_ASAP7_75t_L g575 ( 
.A1(n_432),
.A2(n_190),
.B(n_188),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_456),
.B(n_183),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_432),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_440),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_440),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_440),
.B(n_176),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_395),
.B(n_236),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_460),
.B(n_335),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_460),
.Y(n_583)
);

AND2x2_ASAP7_75t_SL g584 ( 
.A(n_460),
.B(n_195),
.Y(n_584)
);

INVx6_ASAP7_75t_L g585 ( 
.A(n_441),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_398),
.A2(n_256),
.B1(n_266),
.B2(n_252),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_400),
.B(n_182),
.C(n_181),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_404),
.B(n_355),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_404),
.B(n_292),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_466),
.B(n_405),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_464),
.B(n_166),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_501),
.B(n_168),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_472),
.B(n_493),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_552),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_466),
.A2(n_254),
.B1(n_215),
.B2(n_203),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_491),
.B(n_405),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_477),
.A2(n_280),
.B1(n_246),
.B2(n_231),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_557),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_469),
.B(n_166),
.Y(n_599)
);

BUFx5_ASAP7_75t_L g600 ( 
.A(n_476),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_552),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_484),
.B(n_355),
.Y(n_602)
);

O2A1O1Ixp33_ASAP7_75t_L g603 ( 
.A1(n_468),
.A2(n_368),
.B(n_364),
.C(n_360),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_557),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_520),
.B(n_193),
.Y(n_605)
);

O2A1O1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_468),
.A2(n_368),
.B(n_364),
.C(n_360),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_472),
.B(n_273),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_486),
.B(n_170),
.Y(n_608)
);

O2A1O1Ixp5_ASAP7_75t_L g609 ( 
.A1(n_474),
.A2(n_361),
.B(n_263),
.C(n_295),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_554),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_L g611 ( 
.A(n_471),
.B(n_202),
.C(n_261),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_521),
.B(n_545),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_554),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_559),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_509),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_565),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_486),
.B(n_173),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_559),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_565),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_475),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_534),
.A2(n_274),
.B(n_279),
.Y(n_621)
);

AOI221xp5_ASAP7_75t_L g622 ( 
.A1(n_551),
.A2(n_294),
.B1(n_303),
.B2(n_301),
.C(n_299),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_545),
.B(n_492),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_475),
.Y(n_624)
);

AOI221xp5_ASAP7_75t_L g625 ( 
.A1(n_551),
.A2(n_294),
.B1(n_303),
.B2(n_301),
.C(n_299),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_484),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_588),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_569),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_510),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g630 ( 
.A(n_498),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_513),
.B(n_264),
.Y(n_631)
);

AO221x1_ASAP7_75t_L g632 ( 
.A1(n_586),
.A2(n_218),
.B1(n_199),
.B2(n_282),
.C(n_260),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_480),
.B(n_174),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_576),
.B(n_174),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_572),
.B(n_177),
.Y(n_635)
);

BUFx5_ASAP7_75t_L g636 ( 
.A(n_476),
.Y(n_636)
);

AND2x6_ASAP7_75t_L g637 ( 
.A(n_536),
.B(n_267),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_520),
.A2(n_272),
.B1(n_277),
.B2(n_276),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_501),
.B(n_169),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_506),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_506),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_506),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_481),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_465),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_507),
.B(n_257),
.C(n_197),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_467),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_516),
.B(n_538),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_L g648 ( 
.A(n_502),
.B(n_177),
.C(n_302),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_467),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_481),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_476),
.A2(n_293),
.B1(n_298),
.B2(n_289),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_470),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_476),
.A2(n_293),
.B1(n_298),
.B2(n_285),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_572),
.B(n_285),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_497),
.B(n_287),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_504),
.B(n_296),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_538),
.B(n_296),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_500),
.B(n_216),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_518),
.B(n_193),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_SL g660 ( 
.A(n_500),
.B(n_164),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_524),
.B(n_193),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_530),
.B(n_193),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_465),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_532),
.B(n_193),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_502),
.B(n_216),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_533),
.B(n_193),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_470),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_503),
.B(n_244),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_474),
.A2(n_185),
.B1(n_297),
.B2(n_290),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_503),
.B(n_249),
.C(n_204),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_508),
.B(n_273),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_514),
.A2(n_251),
.B1(n_206),
.B2(n_217),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_479),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_485),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_485),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_479),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_555),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_523),
.B(n_227),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_541),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_523),
.B(n_278),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_529),
.Y(n_681)
);

OAI221xp5_ASAP7_75t_L g682 ( 
.A1(n_489),
.A2(n_221),
.B1(n_283),
.B2(n_290),
.C(n_297),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_529),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_562),
.B(n_169),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_548),
.B(n_359),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_540),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_514),
.A2(n_175),
.B1(n_172),
.B2(n_359),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_573),
.B(n_175),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_562),
.B(n_172),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_580),
.B(n_146),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_487),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_581),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_514),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_584),
.B(n_61),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_584),
.B(n_144),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_539),
.B(n_141),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_548),
.B(n_21),
.Y(n_697)
);

AO221x1_ASAP7_75t_L g698 ( 
.A1(n_543),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.C(n_29),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_508),
.B(n_542),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_511),
.B(n_26),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_537),
.B(n_29),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_526),
.B(n_65),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_580),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_537),
.B(n_544),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_487),
.B(n_138),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_514),
.Y(n_706)
);

AND2x6_ASAP7_75t_SL g707 ( 
.A(n_564),
.B(n_30),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_575),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_708)
);

BUFx8_ASAP7_75t_L g709 ( 
.A(n_540),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_580),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_522),
.B(n_108),
.Y(n_711)
);

BUFx5_ASAP7_75t_L g712 ( 
.A(n_531),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_483),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_525),
.B(n_104),
.Y(n_714)
);

AND2x6_ASAP7_75t_L g715 ( 
.A(n_535),
.B(n_98),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_496),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_483),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_488),
.Y(n_718)
);

NOR3xp33_ASAP7_75t_L g719 ( 
.A(n_587),
.B(n_32),
.C(n_34),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_580),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_630),
.B(n_589),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_692),
.B(n_699),
.Y(n_722)
);

NOR2x1_ASAP7_75t_L g723 ( 
.A(n_647),
.B(n_563),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_612),
.A2(n_550),
.B(n_582),
.Y(n_724)
);

CKINVDCx10_ASAP7_75t_R g725 ( 
.A(n_709),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_677),
.Y(n_726)
);

AOI21x1_ASAP7_75t_L g727 ( 
.A1(n_605),
.A2(n_578),
.B(n_577),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_598),
.Y(n_728)
);

OR2x6_ASAP7_75t_L g729 ( 
.A(n_629),
.B(n_478),
.Y(n_729)
);

OAI21xp33_ASAP7_75t_L g730 ( 
.A1(n_591),
.A2(n_490),
.B(n_478),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_692),
.A2(n_716),
.B1(n_591),
.B2(n_596),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_SL g732 ( 
.A(n_615),
.B(n_528),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_634),
.B(n_496),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_L g734 ( 
.A(n_634),
.B(n_512),
.C(n_482),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_716),
.B(n_549),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_633),
.B(n_505),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_700),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_640),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_604),
.Y(n_739)
);

NOR3xp33_ASAP7_75t_L g740 ( 
.A(n_658),
.B(n_541),
.C(n_473),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_633),
.B(n_547),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_677),
.Y(n_742)
);

NOR3xp33_ASAP7_75t_SL g743 ( 
.A(n_682),
.B(n_478),
.C(n_528),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_642),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_668),
.A2(n_473),
.B(n_583),
.C(n_547),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_642),
.B(n_528),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_635),
.B(n_478),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_650),
.B(n_549),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_650),
.A2(n_546),
.B(n_556),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_685),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_626),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_675),
.A2(n_535),
.B(n_553),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_685),
.Y(n_753)
);

BUFx2_ASAP7_75t_SL g754 ( 
.A(n_686),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_654),
.B(n_579),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_595),
.A2(n_585),
.B1(n_566),
.B2(n_561),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_685),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_626),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_595),
.A2(n_585),
.B1(n_566),
.B2(n_561),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_641),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_654),
.B(n_579),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_681),
.A2(n_683),
.B(n_705),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_680),
.A2(n_553),
.B(n_494),
.C(n_488),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_620),
.B(n_494),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_660),
.B(n_570),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_624),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_607),
.B(n_575),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_643),
.B(n_531),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_644),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_674),
.B(n_531),
.Y(n_770)
);

OAI21xp33_ASAP7_75t_L g771 ( 
.A1(n_684),
.A2(n_527),
.B(n_519),
.Y(n_771)
);

BUFx12f_ASAP7_75t_L g772 ( 
.A(n_709),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_680),
.A2(n_517),
.B(n_519),
.C(n_527),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_599),
.A2(n_517),
.B(n_531),
.C(n_571),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_669),
.B(n_499),
.C(n_560),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_593),
.B(n_585),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_594),
.B(n_574),
.Y(n_777)
);

O2A1O1Ixp5_ASAP7_75t_L g778 ( 
.A1(n_694),
.A2(n_574),
.B(n_571),
.C(n_568),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_601),
.B(n_567),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_610),
.B(n_574),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_684),
.B(n_566),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_R g782 ( 
.A(n_679),
.B(n_566),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_613),
.B(n_574),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_711),
.A2(n_567),
.B(n_560),
.Y(n_784)
);

CKINVDCx8_ASAP7_75t_R g785 ( 
.A(n_707),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_714),
.A2(n_567),
.B(n_560),
.Y(n_786)
);

NOR2xp67_ASAP7_75t_L g787 ( 
.A(n_638),
.B(n_79),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_694),
.A2(n_567),
.B(n_560),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_616),
.B(n_574),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_663),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_619),
.B(n_499),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_695),
.A2(n_499),
.B(n_571),
.Y(n_792)
);

AOI21xp33_ASAP7_75t_L g793 ( 
.A1(n_689),
.A2(n_37),
.B(n_40),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_695),
.A2(n_571),
.B(n_568),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_627),
.B(n_568),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_704),
.B(n_688),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_690),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_602),
.B(n_558),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_608),
.B(n_37),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_602),
.B(n_558),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_646),
.Y(n_801)
);

NOR2x1_ASAP7_75t_L g802 ( 
.A(n_611),
.B(n_87),
.Y(n_802)
);

O2A1O1Ixp33_ASAP7_75t_SL g803 ( 
.A1(n_702),
.A2(n_558),
.B(n_42),
.C(n_44),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_659),
.A2(n_558),
.B(n_80),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_661),
.A2(n_70),
.B(n_42),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_649),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_662),
.A2(n_41),
.B(n_44),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_652),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_664),
.A2(n_45),
.B(n_47),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_666),
.A2(n_52),
.B(n_631),
.Y(n_810)
);

BUFx8_ASAP7_75t_SL g811 ( 
.A(n_671),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_701),
.A2(n_52),
.B(n_697),
.C(n_708),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_667),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_673),
.A2(n_676),
.B(n_718),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_648),
.B(n_670),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_669),
.B(n_622),
.C(n_625),
.Y(n_816)
);

NOR3xp33_ASAP7_75t_L g817 ( 
.A(n_617),
.B(n_657),
.C(n_665),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_713),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_592),
.B(n_639),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_SL g820 ( 
.A(n_690),
.B(n_693),
.Y(n_820)
);

AO22x1_ASAP7_75t_L g821 ( 
.A1(n_719),
.A2(n_648),
.B1(n_670),
.B2(n_706),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_708),
.A2(n_651),
.B1(n_653),
.B2(n_691),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_597),
.B(n_672),
.C(n_645),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_720),
.A2(n_710),
.B(n_703),
.C(n_621),
.Y(n_824)
);

OAI321xp33_ASAP7_75t_L g825 ( 
.A1(n_691),
.A2(n_597),
.A3(n_687),
.B1(n_678),
.B2(n_656),
.C(n_655),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_637),
.A2(n_628),
.B1(n_618),
.B2(n_614),
.Y(n_826)
);

BUFx12f_ASAP7_75t_L g827 ( 
.A(n_715),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_637),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_637),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_717),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_609),
.A2(n_696),
.B(n_603),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_637),
.B(n_600),
.Y(n_832)
);

NAND3xp33_ASAP7_75t_L g833 ( 
.A(n_606),
.B(n_632),
.C(n_698),
.Y(n_833)
);

NAND2x1p5_ASAP7_75t_L g834 ( 
.A(n_600),
.B(n_636),
.Y(n_834)
);

NAND2x1p5_ASAP7_75t_L g835 ( 
.A(n_600),
.B(n_636),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_715),
.A2(n_471),
.B(n_468),
.C(n_650),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_715),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_715),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_636),
.A2(n_466),
.B1(n_591),
.B2(n_692),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_712),
.A2(n_612),
.B(n_515),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_715),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_712),
.B(n_692),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_712),
.A2(n_612),
.B(n_515),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_712),
.A2(n_477),
.B(n_495),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_650),
.A2(n_471),
.B(n_468),
.C(n_590),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_598),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_709),
.Y(n_847)
);

NAND2x1p5_ASAP7_75t_L g848 ( 
.A(n_642),
.B(n_690),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_692),
.B(n_548),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_692),
.B(n_548),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_598),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_630),
.B(n_596),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_642),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_612),
.A2(n_623),
.B(n_630),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_650),
.A2(n_471),
.B(n_468),
.C(n_590),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_612),
.A2(n_623),
.B(n_630),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_612),
.A2(n_623),
.B(n_630),
.Y(n_857)
);

BUFx8_ASAP7_75t_L g858 ( 
.A(n_629),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_642),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_630),
.B(n_596),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_591),
.A2(n_634),
.B(n_464),
.C(n_477),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_612),
.A2(n_623),
.B(n_630),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_640),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_591),
.A2(n_466),
.B1(n_692),
.B2(n_623),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_612),
.A2(n_623),
.B(n_630),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_861),
.A2(n_793),
.B(n_731),
.C(n_815),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_852),
.B(n_860),
.Y(n_867)
);

OAI21x1_ASAP7_75t_L g868 ( 
.A1(n_840),
.A2(n_843),
.B(n_727),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_822),
.A2(n_856),
.B(n_854),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_738),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_816),
.A2(n_733),
.B1(n_864),
.B2(n_839),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_858),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_858),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_721),
.B(n_722),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_760),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_736),
.B(n_747),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_820),
.B(n_751),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_753),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_781),
.B(n_776),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_751),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_730),
.A2(n_812),
.B(n_823),
.C(n_825),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_857),
.A2(n_865),
.B(n_862),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_799),
.A2(n_845),
.B(n_855),
.C(n_796),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_863),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_SL g885 ( 
.A1(n_834),
.A2(n_835),
.B(n_832),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_767),
.B(n_755),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_766),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_737),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_764),
.Y(n_889)
);

AO31x2_ASAP7_75t_L g890 ( 
.A1(n_745),
.A2(n_763),
.A3(n_773),
.B(n_824),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_761),
.B(n_819),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_734),
.B(n_757),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_787),
.A2(n_833),
.B1(n_817),
.B2(n_790),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_797),
.B(n_750),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_811),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_748),
.B(n_762),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_859),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_797),
.A2(n_848),
.B1(n_743),
.B2(n_775),
.Y(n_898)
);

AND2x6_ASAP7_75t_SL g899 ( 
.A(n_729),
.B(n_725),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_751),
.B(n_758),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_821),
.B(n_848),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_772),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_849),
.B(n_850),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_754),
.B(n_729),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_728),
.B(n_739),
.Y(n_905)
);

AO21x1_ASAP7_75t_L g906 ( 
.A1(n_844),
.A2(n_836),
.B(n_810),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_729),
.B(n_723),
.Y(n_907)
);

NOR2x1_ASAP7_75t_R g908 ( 
.A(n_847),
.B(n_758),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_782),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_846),
.B(n_851),
.Y(n_910)
);

OAI222xp33_ASAP7_75t_L g911 ( 
.A1(n_807),
.A2(n_809),
.B1(n_785),
.B2(n_810),
.C1(n_805),
.C2(n_802),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_732),
.B(n_740),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_744),
.Y(n_913)
);

AND2x6_ASAP7_75t_SL g914 ( 
.A(n_765),
.B(n_735),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_741),
.B(n_742),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_758),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_756),
.A2(n_759),
.B1(n_837),
.B2(n_841),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_742),
.B(n_769),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_853),
.B(n_859),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_726),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_803),
.A2(n_746),
.B(n_777),
.C(n_780),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_853),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_744),
.B(n_818),
.Y(n_923)
);

AO21x1_ASAP7_75t_L g924 ( 
.A1(n_831),
.A2(n_805),
.B(n_842),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_801),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_837),
.A2(n_841),
.B1(n_838),
.B2(n_828),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_771),
.B(n_744),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_806),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_726),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_778),
.A2(n_774),
.B(n_783),
.C(n_789),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_813),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_749),
.B(n_726),
.Y(n_932)
);

AO31x2_ASAP7_75t_L g933 ( 
.A1(n_794),
.A2(n_724),
.A3(n_792),
.B(n_807),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_830),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_808),
.B(n_752),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_SL g936 ( 
.A(n_827),
.B(n_829),
.Y(n_936)
);

AOI21xp33_ASAP7_75t_L g937 ( 
.A1(n_768),
.A2(n_770),
.B(n_795),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_794),
.A2(n_792),
.B(n_724),
.C(n_826),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_837),
.B(n_809),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_814),
.Y(n_940)
);

AND2x2_ASAP7_75t_SL g941 ( 
.A(n_798),
.B(n_800),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_779),
.B(n_791),
.Y(n_942)
);

AO31x2_ASAP7_75t_L g943 ( 
.A1(n_804),
.A2(n_788),
.A3(n_784),
.B(n_786),
.Y(n_943)
);

NOR2x1_ASAP7_75t_L g944 ( 
.A(n_849),
.B(n_850),
.Y(n_944)
);

AOI221xp5_ASAP7_75t_SL g945 ( 
.A1(n_861),
.A2(n_822),
.B1(n_595),
.B2(n_812),
.C(n_864),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_822),
.A2(n_865),
.B(n_856),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_852),
.B(n_860),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_852),
.B(n_860),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_725),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_852),
.B(n_860),
.Y(n_950)
);

OAI21x1_ASAP7_75t_SL g951 ( 
.A1(n_844),
.A2(n_836),
.B(n_812),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_861),
.A2(n_747),
.B(n_591),
.C(n_730),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_751),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_822),
.A2(n_865),
.B(n_856),
.Y(n_954)
);

AOI221xp5_ASAP7_75t_SL g955 ( 
.A1(n_861),
.A2(n_822),
.B1(n_595),
.B2(n_812),
.C(n_864),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_852),
.B(n_860),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_861),
.A2(n_747),
.B(n_591),
.C(n_730),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_840),
.A2(n_843),
.B(n_727),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_840),
.A2(n_843),
.B(n_727),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_738),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_852),
.B(n_860),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_852),
.B(n_860),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_738),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_751),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_722),
.B(n_511),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_858),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_861),
.A2(n_747),
.B(n_591),
.C(n_730),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_852),
.B(n_860),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_722),
.Y(n_969)
);

NOR2x1_ASAP7_75t_L g970 ( 
.A(n_849),
.B(n_850),
.Y(n_970)
);

AO31x2_ASAP7_75t_L g971 ( 
.A1(n_745),
.A2(n_864),
.A3(n_839),
.B(n_822),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_858),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_852),
.B(n_860),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_738),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_751),
.Y(n_975)
);

OAI22x1_ASAP7_75t_L g976 ( 
.A1(n_816),
.A2(n_747),
.B1(n_736),
.B2(n_799),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_722),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_861),
.A2(n_747),
.B(n_591),
.C(n_730),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_731),
.B(n_548),
.Y(n_979)
);

OAI21x1_ASAP7_75t_SL g980 ( 
.A1(n_844),
.A2(n_836),
.B(n_812),
.Y(n_980)
);

CKINVDCx8_ASAP7_75t_R g981 ( 
.A(n_725),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_822),
.A2(n_865),
.B(n_856),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_722),
.Y(n_983)
);

OAI21x1_ASAP7_75t_SL g984 ( 
.A1(n_844),
.A2(n_836),
.B(n_812),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_722),
.B(n_819),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_822),
.A2(n_865),
.B(n_856),
.Y(n_986)
);

AO31x2_ASAP7_75t_L g987 ( 
.A1(n_745),
.A2(n_864),
.A3(n_839),
.B(n_822),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_797),
.B(n_853),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_852),
.B(n_860),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_736),
.B(n_692),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_858),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_897),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_976),
.A2(n_876),
.B1(n_871),
.B2(n_891),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_894),
.B(n_900),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_894),
.B(n_900),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_870),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_990),
.B(n_965),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_880),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_875),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_884),
.Y(n_1000)
);

INVxp67_ASAP7_75t_SL g1001 ( 
.A(n_867),
.Y(n_1001)
);

CKINVDCx6p67_ASAP7_75t_R g1002 ( 
.A(n_902),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_985),
.B(n_969),
.Y(n_1003)
);

AND2x6_ASAP7_75t_L g1004 ( 
.A(n_897),
.B(n_922),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_878),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_977),
.B(n_983),
.Y(n_1006)
);

OAI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_867),
.A2(n_973),
.B1(n_968),
.B2(n_962),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_874),
.B(n_962),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_968),
.B(n_973),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_989),
.B(n_947),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_960),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_907),
.B(n_904),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_887),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_880),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_963),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_904),
.B(n_913),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_974),
.Y(n_1017)
);

AOI21xp33_ASAP7_75t_SL g1018 ( 
.A1(n_903),
.A2(n_949),
.B(n_912),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_928),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_981),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_979),
.A2(n_948),
.B1(n_961),
.B2(n_956),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_904),
.B(n_964),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_879),
.B(n_888),
.Y(n_1023)
);

OR2x6_ASAP7_75t_SL g1024 ( 
.A(n_909),
.B(n_901),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_892),
.B(n_889),
.Y(n_1025)
);

BUFx4f_ASAP7_75t_L g1026 ( 
.A(n_880),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_950),
.A2(n_952),
.B1(n_978),
.B2(n_957),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_916),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_905),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_872),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_910),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_964),
.B(n_975),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_916),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_967),
.A2(n_883),
.B(n_881),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_922),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_916),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_886),
.B(n_879),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_945),
.B(n_955),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_953),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_923),
.B(n_925),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_951),
.A2(n_984),
.B1(n_980),
.B2(n_954),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_890),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_890),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_908),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_953),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_869),
.A2(n_982),
.B1(n_954),
.B2(n_986),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_931),
.B(n_944),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_890),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_945),
.B(n_955),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_893),
.B(n_896),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_896),
.B(n_970),
.Y(n_1051)
);

BUFx10_ASAP7_75t_L g1052 ( 
.A(n_899),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_934),
.B(n_939),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_918),
.Y(n_1054)
);

HAxp5_ASAP7_75t_L g1055 ( 
.A(n_914),
.B(n_972),
.CON(n_1055),
.SN(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_933),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_929),
.B(n_877),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_895),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_927),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_869),
.A2(n_982),
.B1(n_946),
.B2(n_906),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_941),
.B(n_917),
.Y(n_1061)
);

AOI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_921),
.A2(n_942),
.B(n_932),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_924),
.A2(n_940),
.B1(n_935),
.B2(n_882),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_975),
.B(n_929),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_920),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_933),
.Y(n_1066)
);

AND2x6_ASAP7_75t_L g1067 ( 
.A(n_953),
.B(n_920),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_927),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_920),
.B(n_918),
.Y(n_1069)
);

AND2x6_ASAP7_75t_L g1070 ( 
.A(n_915),
.B(n_935),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_898),
.B(n_926),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_971),
.B(n_987),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_919),
.Y(n_1073)
);

BUFx12f_ASAP7_75t_L g1074 ( 
.A(n_991),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_966),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_919),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_971),
.B(n_987),
.Y(n_1077)
);

INVx3_ASAP7_75t_SL g1078 ( 
.A(n_873),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_911),
.A2(n_938),
.B(n_930),
.C(n_937),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_971),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_936),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_987),
.B(n_988),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_885),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_868),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_958),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_943),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_959),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_943),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_943),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_894),
.B(n_900),
.Y(n_1090)
);

CKINVDCx8_ASAP7_75t_R g1091 ( 
.A(n_899),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_887),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_870),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_981),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_880),
.Y(n_1095)
);

BUFx4f_ASAP7_75t_L g1096 ( 
.A(n_880),
.Y(n_1096)
);

BUFx4f_ASAP7_75t_L g1097 ( 
.A(n_880),
.Y(n_1097)
);

BUFx10_ASAP7_75t_L g1098 ( 
.A(n_949),
.Y(n_1098)
);

INVxp67_ASAP7_75t_SL g1099 ( 
.A(n_867),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_891),
.B(n_876),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_965),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_878),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_SL g1103 ( 
.A1(n_876),
.A2(n_816),
.B1(n_822),
.B2(n_660),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_870),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_876),
.B(n_990),
.Y(n_1105)
);

NAND2x1p5_ASAP7_75t_L g1106 ( 
.A(n_900),
.B(n_964),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_876),
.B(n_990),
.Y(n_1107)
);

INVx8_ASAP7_75t_L g1108 ( 
.A(n_900),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_878),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_880),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_952),
.A2(n_861),
.B(n_957),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_952),
.A2(n_861),
.B(n_967),
.C(n_957),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_969),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_985),
.B(n_722),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_SL g1115 ( 
.A1(n_883),
.A2(n_822),
.B(n_861),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_952),
.A2(n_861),
.B(n_967),
.C(n_957),
.Y(n_1116)
);

BUFx12f_ASAP7_75t_L g1117 ( 
.A(n_949),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_870),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_969),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_866),
.A2(n_816),
.B(n_861),
.C(n_876),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_876),
.A2(n_861),
.B1(n_962),
.B2(n_867),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_870),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_894),
.B(n_900),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_969),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_870),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_880),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_965),
.Y(n_1127)
);

BUFx12f_ASAP7_75t_L g1128 ( 
.A(n_949),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_985),
.B(n_722),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_894),
.B(n_900),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_894),
.B(n_900),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1069),
.B(n_1012),
.Y(n_1132)
);

INVx6_ASAP7_75t_L g1133 ( 
.A(n_1039),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_1108),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_1069),
.B(n_1012),
.Y(n_1135)
);

BUFx12f_ASAP7_75t_L g1136 ( 
.A(n_1020),
.Y(n_1136)
);

NAND2x1p5_ASAP7_75t_L g1137 ( 
.A(n_1039),
.B(n_1076),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1004),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_1108),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_993),
.B(n_1103),
.Y(n_1140)
);

BUFx12f_ASAP7_75t_L g1141 ( 
.A(n_1094),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1105),
.B(n_1107),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1026),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1125),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_993),
.B(n_1103),
.Y(n_1145)
);

OAI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1100),
.A2(n_1107),
.B1(n_1105),
.B2(n_1010),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_996),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_999),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1034),
.A2(n_1111),
.B1(n_1046),
.B2(n_1027),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1026),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_SL g1151 ( 
.A1(n_1091),
.A2(n_997),
.B1(n_1081),
.B2(n_1030),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1120),
.A2(n_1115),
.B(n_1121),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1011),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1015),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1017),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_1096),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1046),
.A2(n_1050),
.B1(n_1041),
.B2(n_1114),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_997),
.B(n_1101),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1129),
.B(n_1008),
.Y(n_1159)
);

BUFx2_ASAP7_75t_SL g1160 ( 
.A(n_1013),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1127),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1053),
.B(n_1022),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1041),
.A2(n_1061),
.B1(n_1071),
.B2(n_1037),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1120),
.A2(n_1021),
.B(n_1007),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1023),
.A2(n_1025),
.B1(n_1003),
.B2(n_1099),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1061),
.A2(n_1071),
.B1(n_1060),
.B2(n_1023),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1009),
.B(n_1001),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1059),
.B(n_1068),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1096),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1068),
.B(n_1054),
.Y(n_1170)
);

OAI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1001),
.A2(n_1099),
.B1(n_1024),
.B2(n_1018),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1093),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1104),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1118),
.Y(n_1174)
);

INVx1_ASAP7_75t_SL g1175 ( 
.A(n_1005),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1122),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1119),
.Y(n_1177)
);

BUFx2_ASAP7_75t_R g1178 ( 
.A(n_1058),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1060),
.A2(n_1021),
.B1(n_1051),
.B2(n_1007),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_SL g1180 ( 
.A1(n_1038),
.A2(n_1049),
.B1(n_1083),
.B2(n_1044),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1070),
.A2(n_1082),
.B1(n_1006),
.B2(n_1102),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1019),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_SL g1183 ( 
.A1(n_1047),
.A2(n_1124),
.B1(n_1119),
.B2(n_1057),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1004),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_1112),
.B(n_1116),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_1109),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1029),
.B(n_1031),
.Y(n_1187)
);

INVx6_ASAP7_75t_L g1188 ( 
.A(n_994),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1097),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1124),
.Y(n_1190)
);

INVx8_ASAP7_75t_L g1191 ( 
.A(n_1067),
.Y(n_1191)
);

BUFx4f_ASAP7_75t_SL g1192 ( 
.A(n_1117),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1084),
.A2(n_1086),
.B(n_1079),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1070),
.A2(n_1080),
.B1(n_1062),
.B2(n_1077),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1040),
.B(n_1113),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1113),
.B(n_1092),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1070),
.A2(n_1072),
.B1(n_1088),
.B2(n_1016),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1004),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1042),
.B(n_1043),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1028),
.Y(n_1200)
);

BUFx2_ASAP7_75t_SL g1201 ( 
.A(n_998),
.Y(n_1201)
);

CKINVDCx11_ASAP7_75t_R g1202 ( 
.A(n_1098),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1028),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1022),
.A2(n_1075),
.B1(n_994),
.B2(n_995),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_995),
.B(n_1131),
.Y(n_1205)
);

OA21x2_ASAP7_75t_L g1206 ( 
.A1(n_1063),
.A2(n_1066),
.B(n_1056),
.Y(n_1206)
);

NAND2x1p5_ASAP7_75t_L g1207 ( 
.A(n_1076),
.B(n_992),
.Y(n_1207)
);

CKINVDCx6p67_ASAP7_75t_R g1208 ( 
.A(n_1128),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1043),
.B(n_1048),
.Y(n_1209)
);

BUFx4f_ASAP7_75t_SL g1210 ( 
.A(n_1074),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1090),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1090),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1063),
.B(n_1035),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1089),
.Y(n_1214)
);

AO21x1_ASAP7_75t_SL g1215 ( 
.A1(n_1073),
.A2(n_1070),
.B(n_1087),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1016),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1097),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1123),
.B(n_1131),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1085),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1085),
.A2(n_1073),
.B(n_1130),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1123),
.B(n_1130),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1085),
.A2(n_1106),
.B(n_1045),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_998),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1070),
.A2(n_1078),
.B1(n_1052),
.B2(n_1064),
.Y(n_1224)
);

AOI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1064),
.A2(n_1032),
.B(n_1065),
.Y(n_1225)
);

INVxp67_ASAP7_75t_SL g1226 ( 
.A(n_1106),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1014),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1014),
.Y(n_1228)
);

INVx4_ASAP7_75t_L g1229 ( 
.A(n_1067),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1045),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1098),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1110),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1032),
.A2(n_1126),
.B(n_1033),
.Y(n_1233)
);

CKINVDCx6p67_ASAP7_75t_R g1234 ( 
.A(n_1002),
.Y(n_1234)
);

INVx4_ASAP7_75t_SL g1235 ( 
.A(n_1067),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1055),
.A2(n_1036),
.B(n_1095),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1095),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1095),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1126),
.A2(n_876),
.B1(n_1100),
.B2(n_1105),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1126),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1052),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1000),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1177),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1199),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1199),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1202),
.Y(n_1246)
);

AO21x1_ASAP7_75t_SL g1247 ( 
.A1(n_1152),
.A2(n_1164),
.B(n_1149),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1199),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_1175),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1185),
.B(n_1165),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1199),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1190),
.Y(n_1252)
);

OAI21xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1163),
.A2(n_1166),
.B(n_1145),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1209),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1209),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1170),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1185),
.B(n_1167),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1186),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1215),
.Y(n_1259)
);

OA21x2_ASAP7_75t_L g1260 ( 
.A1(n_1193),
.A2(n_1194),
.B(n_1179),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1140),
.B(n_1145),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1206),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1214),
.A2(n_1213),
.B(n_1171),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1140),
.B(n_1213),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1146),
.B(n_1142),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1185),
.B(n_1170),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1202),
.Y(n_1267)
);

AO21x2_ASAP7_75t_L g1268 ( 
.A1(n_1219),
.A2(n_1220),
.B(n_1236),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1185),
.B(n_1168),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1168),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1147),
.A2(n_1182),
.B(n_1176),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1222),
.B(n_1138),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1157),
.B(n_1242),
.Y(n_1273)
);

AO21x2_ASAP7_75t_L g1274 ( 
.A1(n_1148),
.A2(n_1153),
.B(n_1174),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1142),
.B(n_1159),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1239),
.B(n_1180),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_1192),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1161),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1158),
.Y(n_1279)
);

AOI21xp33_ASAP7_75t_L g1280 ( 
.A1(n_1158),
.A2(n_1187),
.B(n_1195),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1197),
.B(n_1181),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1144),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1200),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1138),
.A2(n_1198),
.B(n_1184),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1162),
.B(n_1132),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1154),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1155),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1162),
.B(n_1132),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1235),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1172),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1203),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1162),
.B(n_1132),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1228),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1173),
.Y(n_1294)
);

INVx8_ASAP7_75t_L g1295 ( 
.A(n_1191),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1225),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1133),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1225),
.Y(n_1298)
);

NOR2xp67_ASAP7_75t_R g1299 ( 
.A(n_1156),
.B(n_1229),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1135),
.B(n_1211),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1215),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1135),
.B(n_1183),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1184),
.A2(n_1198),
.B(n_1224),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1216),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1232),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1204),
.A2(n_1151),
.B1(n_1160),
.B2(n_1212),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1135),
.B(n_1237),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1207),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1207),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1230),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1241),
.A2(n_1231),
.B1(n_1196),
.B2(n_1188),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1272),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1272),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1262),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1272),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1257),
.B(n_1196),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1269),
.B(n_1238),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1269),
.B(n_1238),
.Y(n_1318)
);

NOR2x1_ASAP7_75t_L g1319 ( 
.A(n_1296),
.B(n_1298),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1264),
.B(n_1238),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1257),
.B(n_1226),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1263),
.B(n_1250),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1264),
.B(n_1240),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1272),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1255),
.B(n_1218),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1255),
.B(n_1218),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1293),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1255),
.B(n_1218),
.Y(n_1328)
);

OAI221xp5_ASAP7_75t_L g1329 ( 
.A1(n_1276),
.A2(n_1241),
.B1(n_1221),
.B2(n_1205),
.C(n_1188),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1303),
.Y(n_1330)
);

AOI221xp5_ASAP7_75t_L g1331 ( 
.A1(n_1253),
.A2(n_1231),
.B1(n_1156),
.B2(n_1217),
.C(n_1150),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1262),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1271),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1263),
.B(n_1223),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1265),
.B(n_1223),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1271),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1266),
.B(n_1188),
.Y(n_1337)
);

NOR2x1_ASAP7_75t_L g1338 ( 
.A(n_1296),
.B(n_1233),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1266),
.B(n_1188),
.Y(n_1339)
);

AND2x2_ASAP7_75t_SL g1340 ( 
.A(n_1260),
.B(n_1229),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1254),
.B(n_1227),
.Y(n_1341)
);

INVxp67_ASAP7_75t_SL g1342 ( 
.A(n_1298),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1284),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1244),
.B(n_1245),
.Y(n_1344)
);

NAND2xp33_ASAP7_75t_R g1345 ( 
.A(n_1246),
.B(n_1178),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1271),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1274),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1268),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1254),
.B(n_1227),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1303),
.Y(n_1350)
);

NAND2x1_ASAP7_75t_L g1351 ( 
.A(n_1289),
.B(n_1229),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1261),
.B(n_1137),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1305),
.Y(n_1353)
);

INVx4_ASAP7_75t_L g1354 ( 
.A(n_1289),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1263),
.B(n_1235),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1263),
.B(n_1235),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1261),
.B(n_1137),
.Y(n_1357)
);

OR2x6_ASAP7_75t_L g1358 ( 
.A(n_1259),
.B(n_1191),
.Y(n_1358)
);

OAI221xp5_ASAP7_75t_L g1359 ( 
.A1(n_1253),
.A2(n_1156),
.B1(n_1169),
.B2(n_1217),
.C(n_1150),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1312),
.B(n_1324),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1316),
.B(n_1243),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1329),
.A2(n_1311),
.B(n_1280),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1331),
.A2(n_1311),
.B(n_1306),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1331),
.A2(n_1247),
.B1(n_1329),
.B2(n_1359),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1359),
.A2(n_1247),
.B1(n_1250),
.B2(n_1281),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_SL g1366 ( 
.A(n_1354),
.B(n_1267),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1316),
.B(n_1278),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1353),
.B(n_1252),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_L g1369 ( 
.A(n_1335),
.B(n_1279),
.C(n_1275),
.Y(n_1369)
);

AND2x2_ASAP7_75t_SL g1370 ( 
.A(n_1340),
.B(n_1260),
.Y(n_1370)
);

NAND3xp33_ASAP7_75t_L g1371 ( 
.A(n_1335),
.B(n_1283),
.C(n_1291),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1321),
.B(n_1249),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1327),
.B(n_1252),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1324),
.B(n_1313),
.Y(n_1374)
);

NAND4xp25_ASAP7_75t_L g1375 ( 
.A(n_1321),
.B(n_1258),
.C(n_1287),
.D(n_1286),
.Y(n_1375)
);

NAND3xp33_ASAP7_75t_L g1376 ( 
.A(n_1322),
.B(n_1281),
.C(n_1304),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1323),
.B(n_1256),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1340),
.A2(n_1299),
.B(n_1260),
.Y(n_1378)
);

OAI21xp33_ASAP7_75t_L g1379 ( 
.A1(n_1322),
.A2(n_1273),
.B(n_1302),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1352),
.B(n_1285),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1352),
.B(n_1292),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1357),
.B(n_1288),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1323),
.B(n_1270),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1357),
.A2(n_1289),
.B1(n_1301),
.B2(n_1259),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1320),
.B(n_1270),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1358),
.A2(n_1289),
.B1(n_1259),
.B2(n_1301),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1337),
.A2(n_1302),
.B1(n_1273),
.B2(n_1260),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1313),
.B(n_1245),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1320),
.B(n_1287),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1325),
.B(n_1290),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1325),
.B(n_1290),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1313),
.B(n_1248),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1337),
.B(n_1288),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1334),
.B(n_1294),
.C(n_1310),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1326),
.B(n_1282),
.Y(n_1395)
);

NOR3xp33_ASAP7_75t_L g1396 ( 
.A(n_1338),
.B(n_1308),
.C(n_1309),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1355),
.A2(n_1301),
.B(n_1259),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_SL g1398 ( 
.A1(n_1355),
.A2(n_1301),
.B(n_1259),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1315),
.B(n_1251),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1339),
.B(n_1300),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1315),
.B(n_1344),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_L g1402 ( 
.A(n_1334),
.B(n_1310),
.C(n_1308),
.Y(n_1402)
);

OAI221xp5_ASAP7_75t_SL g1403 ( 
.A1(n_1356),
.A2(n_1234),
.B1(n_1208),
.B2(n_1251),
.C(n_1169),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1328),
.B(n_1341),
.Y(n_1404)
);

OAI221xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1356),
.A2(n_1234),
.B1(n_1208),
.B2(n_1309),
.C(n_1307),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1339),
.B(n_1307),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1340),
.A2(n_1259),
.B1(n_1301),
.B2(n_1295),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1401),
.Y(n_1408)
);

NOR2x1_ASAP7_75t_L g1409 ( 
.A(n_1402),
.B(n_1338),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1390),
.B(n_1314),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1370),
.B(n_1401),
.Y(n_1411)
);

NAND3xp33_ASAP7_75t_L g1412 ( 
.A(n_1362),
.B(n_1319),
.C(n_1341),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1388),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1388),
.Y(n_1414)
);

OAI221xp5_ASAP7_75t_L g1415 ( 
.A1(n_1363),
.A2(n_1345),
.B1(n_1349),
.B2(n_1351),
.C(n_1330),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1394),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1367),
.B(n_1342),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1370),
.B(n_1330),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1394),
.Y(n_1419)
);

INVxp67_ASAP7_75t_L g1420 ( 
.A(n_1369),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1391),
.B(n_1314),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1370),
.B(n_1330),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1374),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1374),
.B(n_1330),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1360),
.Y(n_1425)
);

INVxp67_ASAP7_75t_R g1426 ( 
.A(n_1386),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1392),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1376),
.B(n_1333),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1360),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1399),
.B(n_1343),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1399),
.Y(n_1431)
);

INVxp67_ASAP7_75t_SL g1432 ( 
.A(n_1402),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1378),
.B(n_1350),
.Y(n_1433)
);

NOR2x1_ASAP7_75t_L g1434 ( 
.A(n_1371),
.B(n_1319),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1389),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1361),
.B(n_1342),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1373),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1404),
.B(n_1350),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1395),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1368),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1379),
.B(n_1350),
.Y(n_1441)
);

INVxp67_ASAP7_75t_SL g1442 ( 
.A(n_1371),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1383),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1376),
.B(n_1332),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1379),
.B(n_1350),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1387),
.B(n_1348),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1411),
.B(n_1396),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1420),
.A2(n_1364),
.B1(n_1365),
.B2(n_1369),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1416),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1411),
.B(n_1407),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1416),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1419),
.B(n_1377),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1419),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1420),
.B(n_1380),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1440),
.B(n_1381),
.Y(n_1455)
);

OAI211xp5_ASAP7_75t_L g1456 ( 
.A1(n_1442),
.A2(n_1375),
.B(n_1372),
.C(n_1403),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1425),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1444),
.B(n_1385),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1411),
.B(n_1397),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1437),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1415),
.A2(n_1301),
.B1(n_1366),
.B2(n_1384),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1425),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1410),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1418),
.B(n_1398),
.Y(n_1464)
);

NAND2x1p5_ASAP7_75t_L g1465 ( 
.A(n_1409),
.B(n_1348),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1418),
.B(n_1343),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1444),
.B(n_1333),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1410),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1440),
.B(n_1382),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1437),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1413),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1418),
.B(n_1317),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1443),
.B(n_1136),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1442),
.B(n_1336),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1432),
.B(n_1336),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1413),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1440),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1413),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1421),
.Y(n_1479)
);

AOI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1412),
.A2(n_1400),
.B1(n_1405),
.B2(n_1406),
.C(n_1393),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1422),
.B(n_1317),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1414),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1422),
.B(n_1343),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1414),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1422),
.B(n_1318),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1463),
.B(n_1432),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1463),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1459),
.B(n_1426),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1459),
.B(n_1426),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1449),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1465),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1468),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1454),
.B(n_1412),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1449),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1457),
.B(n_1409),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1468),
.Y(n_1496)
);

OAI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1448),
.A2(n_1415),
.B1(n_1434),
.B2(n_1358),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1457),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1479),
.B(n_1428),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1479),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1460),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1451),
.B(n_1428),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1451),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1450),
.B(n_1434),
.Y(n_1504)
);

INVxp67_ASAP7_75t_L g1505 ( 
.A(n_1452),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1453),
.B(n_1428),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1448),
.B(n_1443),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1478),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1464),
.B(n_1433),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1455),
.B(n_1435),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1452),
.B(n_1435),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1453),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1478),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1456),
.B(n_1439),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1464),
.B(n_1433),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1478),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1450),
.B(n_1447),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1462),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1482),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1447),
.B(n_1433),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1458),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1482),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1447),
.B(n_1430),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1482),
.Y(n_1524)
);

AOI311xp33_ASAP7_75t_L g1525 ( 
.A1(n_1470),
.A2(n_1439),
.A3(n_1417),
.B(n_1436),
.C(n_1431),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1484),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1458),
.B(n_1417),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1484),
.A2(n_1347),
.B(n_1346),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1503),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1501),
.B(n_1480),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1486),
.B(n_1474),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1488),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1503),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1495),
.B(n_1447),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1498),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1493),
.B(n_1472),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1528),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1486),
.B(n_1474),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1514),
.B(n_1472),
.Y(n_1539)
);

AOI22x1_ASAP7_75t_L g1540 ( 
.A1(n_1504),
.A2(n_1465),
.B1(n_1141),
.B2(n_1136),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1488),
.B(n_1481),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1497),
.A2(n_1461),
.B1(n_1473),
.B2(n_1446),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1507),
.B(n_1481),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1489),
.B(n_1485),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1528),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1512),
.Y(n_1546)
);

NAND3x1_ASAP7_75t_L g1547 ( 
.A(n_1489),
.B(n_1469),
.C(n_1445),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1517),
.B(n_1485),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1512),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1517),
.B(n_1466),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1490),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1509),
.B(n_1466),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1504),
.A2(n_1446),
.B1(n_1441),
.B2(n_1445),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1527),
.B(n_1475),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1494),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1509),
.B(n_1466),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1498),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1515),
.B(n_1466),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1495),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1504),
.B(n_1477),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1527),
.B(n_1475),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1521),
.A2(n_1520),
.B1(n_1515),
.B2(n_1505),
.Y(n_1562)
);

INVxp67_ASAP7_75t_SL g1563 ( 
.A(n_1495),
.Y(n_1563)
);

AOI222xp33_ASAP7_75t_L g1564 ( 
.A1(n_1518),
.A2(n_1446),
.B1(n_1441),
.B2(n_1445),
.C1(n_1436),
.C2(n_1438),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1529),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1559),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1541),
.B(n_1520),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1532),
.B(n_1518),
.Y(n_1568)
);

O2A1O1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1530),
.A2(n_1465),
.B(n_1491),
.C(n_1506),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1535),
.Y(n_1570)
);

O2A1O1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1532),
.A2(n_1491),
.B(n_1506),
.C(n_1502),
.Y(n_1571)
);

AOI322xp5_ASAP7_75t_L g1572 ( 
.A1(n_1542),
.A2(n_1441),
.A3(n_1525),
.B1(n_1523),
.B2(n_1511),
.C1(n_1491),
.C2(n_1487),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1529),
.Y(n_1573)
);

NAND2x1_ASAP7_75t_L g1574 ( 
.A(n_1534),
.B(n_1523),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1539),
.B(n_1277),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1562),
.B(n_1487),
.Y(n_1576)
);

OAI332xp33_ASAP7_75t_L g1577 ( 
.A1(n_1563),
.A2(n_1502),
.A3(n_1499),
.B1(n_1500),
.B2(n_1492),
.B3(n_1496),
.C1(n_1510),
.C2(n_1519),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_L g1578 ( 
.A(n_1560),
.B(n_1496),
.C(n_1492),
.Y(n_1578)
);

AOI22x1_ASAP7_75t_L g1579 ( 
.A1(n_1557),
.A2(n_1500),
.B1(n_1141),
.B2(n_1499),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1543),
.B(n_1467),
.Y(n_1580)
);

AOI221xp5_ASAP7_75t_L g1581 ( 
.A1(n_1557),
.A2(n_1519),
.B1(n_1524),
.B2(n_1526),
.C(n_1522),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1541),
.B(n_1544),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1533),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1551),
.B(n_1555),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1533),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1559),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1536),
.A2(n_1551),
.B1(n_1555),
.B2(n_1544),
.C(n_1548),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1547),
.A2(n_1483),
.B1(n_1438),
.B2(n_1524),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1546),
.Y(n_1589)
);

OAI31xp33_ASAP7_75t_L g1590 ( 
.A1(n_1534),
.A2(n_1483),
.A3(n_1526),
.B(n_1424),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1582),
.B(n_1548),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1568),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1566),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1576),
.B(n_1554),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1566),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1570),
.B(n_1550),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1576),
.B(n_1554),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1568),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1567),
.B(n_1550),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1587),
.B(n_1534),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1577),
.B(n_1534),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1586),
.B(n_1559),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1574),
.B(n_1559),
.Y(n_1603)
);

NAND2x1_ASAP7_75t_SL g1604 ( 
.A(n_1588),
.B(n_1553),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1575),
.B(n_1564),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1580),
.B(n_1552),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1578),
.B(n_1561),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1565),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1572),
.B(n_1553),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1571),
.B(n_1531),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1609),
.A2(n_1547),
.B1(n_1579),
.B2(n_1540),
.Y(n_1611)
);

NAND3xp33_ASAP7_75t_SL g1612 ( 
.A(n_1601),
.B(n_1569),
.C(n_1581),
.Y(n_1612)
);

NOR3xp33_ASAP7_75t_L g1613 ( 
.A(n_1605),
.B(n_1584),
.C(n_1583),
.Y(n_1613)
);

OAI21xp33_ASAP7_75t_L g1614 ( 
.A1(n_1604),
.A2(n_1584),
.B(n_1573),
.Y(n_1614)
);

OAI21xp33_ASAP7_75t_L g1615 ( 
.A1(n_1600),
.A2(n_1589),
.B(n_1585),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1610),
.A2(n_1607),
.B1(n_1597),
.B2(n_1594),
.Y(n_1616)
);

OAI211xp5_ASAP7_75t_L g1617 ( 
.A1(n_1610),
.A2(n_1590),
.B(n_1540),
.C(n_1549),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1595),
.Y(n_1618)
);

O2A1O1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1592),
.A2(n_1546),
.B(n_1549),
.C(n_1538),
.Y(n_1619)
);

NAND3xp33_ASAP7_75t_L g1620 ( 
.A(n_1598),
.B(n_1538),
.C(n_1531),
.Y(n_1620)
);

NAND5xp2_ASAP7_75t_L g1621 ( 
.A(n_1596),
.B(n_1558),
.C(n_1556),
.D(n_1552),
.E(n_1424),
.Y(n_1621)
);

AOI211x1_ASAP7_75t_L g1622 ( 
.A1(n_1602),
.A2(n_1558),
.B(n_1556),
.C(n_1424),
.Y(n_1622)
);

AOI221xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_1513),
.B2(n_1522),
.C(n_1516),
.Y(n_1623)
);

XNOR2xp5_ASAP7_75t_L g1624 ( 
.A(n_1616),
.B(n_1591),
.Y(n_1624)
);

NOR3x1_ASAP7_75t_L g1625 ( 
.A(n_1612),
.B(n_1593),
.C(n_1608),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1614),
.B(n_1603),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1618),
.B(n_1591),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1620),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1622),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1619),
.Y(n_1630)
);

NOR3xp33_ASAP7_75t_L g1631 ( 
.A(n_1613),
.B(n_1593),
.C(n_1595),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_L g1632 ( 
.A(n_1615),
.B(n_1606),
.C(n_1599),
.Y(n_1632)
);

NOR3x1_ASAP7_75t_L g1633 ( 
.A(n_1617),
.B(n_1611),
.C(n_1621),
.Y(n_1633)
);

NOR2x1_ASAP7_75t_L g1634 ( 
.A(n_1623),
.B(n_1599),
.Y(n_1634)
);

NAND3xp33_ASAP7_75t_L g1635 ( 
.A(n_1628),
.B(n_1606),
.C(n_1513),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1624),
.B(n_1632),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1627),
.Y(n_1637)
);

NAND3xp33_ASAP7_75t_SL g1638 ( 
.A(n_1631),
.B(n_1210),
.C(n_1537),
.Y(n_1638)
);

AOI21xp33_ASAP7_75t_L g1639 ( 
.A1(n_1632),
.A2(n_1516),
.B(n_1508),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_L g1640 ( 
.A(n_1630),
.B(n_1508),
.C(n_1537),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1636),
.A2(n_1629),
.B1(n_1626),
.B2(n_1634),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1637),
.Y(n_1642)
);

AOI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1638),
.A2(n_1635),
.B1(n_1640),
.B2(n_1639),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1637),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1637),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1636),
.A2(n_1625),
.B1(n_1633),
.B2(n_1483),
.Y(n_1646)
);

NAND4xp75_ASAP7_75t_L g1647 ( 
.A(n_1641),
.B(n_1545),
.C(n_1537),
.D(n_1528),
.Y(n_1647)
);

XNOR2xp5_ASAP7_75t_L g1648 ( 
.A(n_1646),
.B(n_1134),
.Y(n_1648)
);

NOR4xp25_ASAP7_75t_SL g1649 ( 
.A(n_1642),
.B(n_1545),
.C(n_1429),
.D(n_1423),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_L g1650 ( 
.A(n_1644),
.B(n_1545),
.Y(n_1650)
);

OAI211xp5_ASAP7_75t_L g1651 ( 
.A1(n_1643),
.A2(n_1189),
.B(n_1143),
.C(n_1191),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1650),
.B(n_1645),
.Y(n_1652)
);

XNOR2xp5_ASAP7_75t_L g1653 ( 
.A(n_1648),
.B(n_1201),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1647),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1652),
.Y(n_1655)
);

XNOR2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1655),
.B(n_1653),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1656),
.A2(n_1654),
.B(n_1651),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1656),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1657),
.A2(n_1649),
.B(n_1483),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1658),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1659),
.A2(n_1189),
.B1(n_1143),
.B2(n_1484),
.C(n_1467),
.Y(n_1661)
);

AO221x1_ASAP7_75t_L g1662 ( 
.A1(n_1660),
.A2(n_1189),
.B1(n_1143),
.B2(n_1408),
.C(n_1427),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1661),
.B(n_1662),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_L g1664 ( 
.A(n_1663),
.B(n_1189),
.C(n_1143),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1664),
.A2(n_1476),
.B1(n_1471),
.B2(n_1429),
.C(n_1423),
.Y(n_1665)
);

AOI211xp5_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1134),
.B(n_1139),
.C(n_1297),
.Y(n_1666)
);


endmodule