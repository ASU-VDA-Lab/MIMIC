module real_aes_7852_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g186 ( .A1(n_0), .A2(n_187), .B(n_188), .C(n_192), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_1), .B(n_182), .Y(n_193) );
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_3), .B(n_147), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_4), .A2(n_128), .B(n_476), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_5), .A2(n_133), .B(n_138), .C(n_512), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_6), .A2(n_128), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_7), .B(n_182), .Y(n_482) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_8), .A2(n_161), .B(n_211), .Y(n_210) );
AND2x6_ASAP7_75t_L g133 ( .A(n_9), .B(n_134), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_10), .A2(n_133), .B(n_138), .C(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g537 ( .A(n_11), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_12), .B(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_12), .B(n_41), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_13), .B(n_191), .Y(n_514) );
INVx1_ASAP7_75t_L g157 ( .A(n_14), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_15), .B(n_147), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_16), .A2(n_148), .B(n_522), .C(n_524), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_17), .B(n_182), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_18), .A2(n_100), .B1(n_112), .B2(n_744), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_19), .B(n_175), .Y(n_566) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_20), .A2(n_138), .B(n_169), .C(n_174), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_21), .A2(n_190), .B(n_205), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_22), .B(n_191), .Y(n_467) );
OAI222xp33_ASAP7_75t_L g447 ( .A1(n_23), .A2(n_448), .B1(n_730), .B2(n_731), .C1(n_737), .C2(n_741), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_23), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_24), .B(n_191), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_25), .Y(n_463) );
INVx1_ASAP7_75t_L g488 ( .A(n_26), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_27), .A2(n_138), .B(n_174), .C(n_214), .Y(n_213) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_28), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_29), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_30), .Y(n_741) );
INVx1_ASAP7_75t_L g564 ( .A(n_31), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_32), .A2(n_128), .B(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g131 ( .A(n_33), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_34), .A2(n_136), .B(n_141), .C(n_151), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_35), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_36), .A2(n_190), .B(n_479), .C(n_481), .Y(n_478) );
INVxp67_ASAP7_75t_L g565 ( .A(n_37), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_38), .B(n_216), .Y(n_215) );
CKINVDCx14_ASAP7_75t_R g477 ( .A(n_39), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_40), .A2(n_138), .B(n_174), .C(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g111 ( .A(n_41), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_42), .A2(n_192), .B(n_535), .C(n_536), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_43), .B(n_167), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_44), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_45), .B(n_147), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_46), .B(n_128), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_47), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_48), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_49), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_50), .A2(n_136), .B(n_151), .C(n_225), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_51), .A2(n_119), .B1(n_120), .B2(n_438), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_51), .Y(n_119) );
INVx1_ASAP7_75t_L g189 ( .A(n_52), .Y(n_189) );
INVx1_ASAP7_75t_L g226 ( .A(n_53), .Y(n_226) );
INVx1_ASAP7_75t_L g500 ( .A(n_54), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_55), .B(n_128), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_56), .Y(n_178) );
CKINVDCx14_ASAP7_75t_R g533 ( .A(n_57), .Y(n_533) );
INVx1_ASAP7_75t_L g134 ( .A(n_58), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_59), .B(n_128), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_60), .B(n_182), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_61), .A2(n_173), .B(n_236), .C(n_238), .Y(n_235) );
INVx1_ASAP7_75t_L g156 ( .A(n_62), .Y(n_156) );
INVx1_ASAP7_75t_SL g480 ( .A(n_63), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_64), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_65), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_66), .B(n_182), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_67), .B(n_148), .Y(n_202) );
INVx1_ASAP7_75t_L g466 ( .A(n_68), .Y(n_466) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_69), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_70), .B(n_144), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_71), .A2(n_138), .B(n_151), .C(n_262), .Y(n_261) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_72), .Y(n_234) );
INVx1_ASAP7_75t_L g108 ( .A(n_73), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_74), .A2(n_128), .B(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_75), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_76), .A2(n_128), .B(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_77), .A2(n_167), .B(n_560), .Y(n_559) );
CKINVDCx16_ASAP7_75t_R g485 ( .A(n_78), .Y(n_485) );
INVx1_ASAP7_75t_L g520 ( .A(n_79), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_80), .B(n_143), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_81), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_82), .A2(n_128), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g523 ( .A(n_83), .Y(n_523) );
INVx2_ASAP7_75t_L g154 ( .A(n_84), .Y(n_154) );
INVx1_ASAP7_75t_L g513 ( .A(n_85), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_86), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_87), .B(n_191), .Y(n_203) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_88), .B(n_105), .C(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g440 ( .A(n_88), .B(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g450 ( .A(n_88), .B(n_442), .Y(n_450) );
INVx2_ASAP7_75t_L g453 ( .A(n_88), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_89), .A2(n_138), .B(n_151), .C(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_90), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g142 ( .A(n_91), .Y(n_142) );
INVxp67_ASAP7_75t_L g239 ( .A(n_92), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_93), .B(n_161), .Y(n_538) );
INVx2_ASAP7_75t_L g503 ( .A(n_94), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_95), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g198 ( .A(n_96), .Y(n_198) );
INVx1_ASAP7_75t_L g263 ( .A(n_97), .Y(n_263) );
AND2x2_ASAP7_75t_L g228 ( .A(n_98), .B(n_153), .Y(n_228) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_SL g746 ( .A(n_102), .Y(n_746) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_109), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g442 ( .A(n_105), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI21x1_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_117), .B(n_446), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g743 ( .A(n_115), .Y(n_743) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_439), .B(n_444), .Y(n_117) );
INVx2_ASAP7_75t_L g438 ( .A(n_120), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_120), .A2(n_732), .B1(n_735), .B2(n_736), .Y(n_731) );
OR3x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_352), .C(n_395), .Y(n_120) );
NAND5xp2_ASAP7_75t_L g121 ( .A(n_122), .B(n_279), .C(n_309), .D(n_326), .E(n_341), .Y(n_121) );
AOI221xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_194), .B1(n_241), .B2(n_247), .C(n_251), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_163), .Y(n_123) );
OR2x2_ASAP7_75t_L g256 ( .A(n_124), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g296 ( .A(n_124), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g314 ( .A(n_124), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_124), .B(n_249), .Y(n_331) );
OR2x2_ASAP7_75t_L g343 ( .A(n_124), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_124), .B(n_302), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_124), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_124), .B(n_280), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_124), .B(n_288), .Y(n_394) );
AND2x2_ASAP7_75t_L g426 ( .A(n_124), .B(n_180), .Y(n_426) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_124), .Y(n_434) );
INVx5_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_125), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g253 ( .A(n_125), .B(n_229), .Y(n_253) );
BUFx2_ASAP7_75t_L g276 ( .A(n_125), .Y(n_276) );
AND2x2_ASAP7_75t_L g305 ( .A(n_125), .B(n_164), .Y(n_305) );
AND2x2_ASAP7_75t_L g360 ( .A(n_125), .B(n_257), .Y(n_360) );
OR2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_158), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_135), .B(n_153), .Y(n_126) );
BUFx2_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
NAND2x1p5_ASAP7_75t_L g199 ( .A(n_129), .B(n_133), .Y(n_199) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
INVx1_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g139 ( .A(n_131), .Y(n_139) );
INVx1_ASAP7_75t_L g206 ( .A(n_131), .Y(n_206) );
INVx1_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_132), .Y(n_145) );
INVx3_ASAP7_75t_L g148 ( .A(n_132), .Y(n_148) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_132), .Y(n_191) );
INVx1_ASAP7_75t_L g216 ( .A(n_132), .Y(n_216) );
INVx4_ASAP7_75t_SL g152 ( .A(n_133), .Y(n_152) );
BUFx3_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_SL g184 ( .A1(n_137), .A2(n_152), .B(n_185), .C(n_186), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_137), .A2(n_152), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_137), .A2(n_152), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g499 ( .A1(n_137), .A2(n_152), .B(n_500), .C(n_501), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_SL g519 ( .A1(n_137), .A2(n_152), .B(n_520), .C(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_137), .A2(n_152), .B(n_533), .C(n_534), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_SL g560 ( .A1(n_137), .A2(n_152), .B(n_561), .C(n_562), .Y(n_560) );
INVx5_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
BUFx3_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_139), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_146), .C(n_149), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_143), .A2(n_149), .B(n_226), .C(n_227), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_143), .A2(n_466), .B(n_467), .C(n_468), .Y(n_465) );
O2A1O1Ixp5_ASAP7_75t_L g512 ( .A1(n_143), .A2(n_468), .B(n_513), .C(n_514), .Y(n_512) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx4_ASAP7_75t_L g237 ( .A(n_145), .Y(n_237) );
INVx2_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_147), .B(n_239), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_147), .A2(n_172), .B(n_488), .C(n_489), .Y(n_487) );
OAI22xp33_ASAP7_75t_L g563 ( .A1(n_147), .A2(n_237), .B1(n_564), .B2(n_565), .Y(n_563) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_148), .B(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g192 ( .A(n_150), .Y(n_192) );
INVx1_ASAP7_75t_L g524 ( .A(n_150), .Y(n_524) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g176 ( .A(n_153), .Y(n_176) );
INVx1_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_153), .A2(n_223), .B(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_153), .A2(n_199), .B(n_485), .C(n_486), .Y(n_484) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_153), .A2(n_531), .B(n_538), .Y(n_530) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AND2x2_ASAP7_75t_L g162 ( .A(n_154), .B(n_155), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx3_ASAP7_75t_L g182 ( .A(n_160), .Y(n_182) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_160), .A2(n_197), .B(n_207), .Y(n_196) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_160), .A2(n_260), .B(n_268), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_160), .B(n_269), .Y(n_268) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_160), .A2(n_462), .B(n_469), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_160), .B(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_160), .B(n_516), .Y(n_515) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_161), .A2(n_212), .B(n_213), .Y(n_211) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_161), .Y(n_231) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_163), .B(n_314), .Y(n_323) );
OAI32xp33_ASAP7_75t_L g337 ( .A1(n_163), .A2(n_273), .A3(n_338), .B1(n_339), .B2(n_340), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_163), .B(n_339), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_163), .B(n_256), .Y(n_380) );
INVx1_ASAP7_75t_SL g409 ( .A(n_163), .Y(n_409) );
NAND4xp25_ASAP7_75t_L g418 ( .A(n_163), .B(n_196), .C(n_360), .D(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g163 ( .A(n_164), .B(n_180), .Y(n_163) );
INVx5_ASAP7_75t_L g250 ( .A(n_164), .Y(n_250) );
AND2x2_ASAP7_75t_L g280 ( .A(n_164), .B(n_181), .Y(n_280) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_164), .Y(n_359) );
AND2x2_ASAP7_75t_L g429 ( .A(n_164), .B(n_376), .Y(n_429) );
OR2x6_ASAP7_75t_L g164 ( .A(n_165), .B(n_177), .Y(n_164) );
AOI21xp5_ASAP7_75t_SL g165 ( .A1(n_166), .A2(n_168), .B(n_175), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_172), .Y(n_169) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_173), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_176), .B(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_179), .A2(n_509), .B(n_515), .Y(n_508) );
AND2x4_ASAP7_75t_L g302 ( .A(n_180), .B(n_250), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_180), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g336 ( .A(n_180), .B(n_257), .Y(n_336) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g249 ( .A(n_181), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g288 ( .A(n_181), .B(n_259), .Y(n_288) );
AND2x2_ASAP7_75t_L g297 ( .A(n_181), .B(n_258), .Y(n_297) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_193), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_190), .B(n_480), .Y(n_479) );
INVx4_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g535 ( .A(n_191), .Y(n_535) );
INVx2_ASAP7_75t_L g468 ( .A(n_192), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g365 ( .A1(n_194), .A2(n_366), .B1(n_368), .B2(n_370), .C1(n_373), .C2(n_374), .Y(n_365) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_218), .Y(n_194) );
AND2x2_ASAP7_75t_L g298 ( .A(n_195), .B(n_299), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g415 ( .A(n_195), .B(n_276), .C(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_210), .Y(n_195) );
INVx5_ASAP7_75t_SL g246 ( .A(n_196), .Y(n_246) );
OAI322xp33_ASAP7_75t_L g251 ( .A1(n_196), .A2(n_252), .A3(n_254), .B1(n_255), .B2(n_270), .C1(n_273), .C2(n_275), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_196), .B(n_244), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_196), .B(n_230), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_199), .A2(n_463), .B(n_464), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_199), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_204), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_204), .A2(n_215), .B(n_217), .Y(n_214) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
INVx2_ASAP7_75t_L g558 ( .A(n_209), .Y(n_558) );
INVx2_ASAP7_75t_L g244 ( .A(n_210), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_210), .B(n_220), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_218), .B(n_283), .Y(n_338) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g317 ( .A(n_219), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_229), .Y(n_219) );
OR2x2_ASAP7_75t_L g245 ( .A(n_220), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_220), .B(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g285 ( .A(n_220), .B(n_230), .Y(n_285) );
AND2x2_ASAP7_75t_L g308 ( .A(n_220), .B(n_244), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_220), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g324 ( .A(n_220), .B(n_283), .Y(n_324) );
AND2x2_ASAP7_75t_L g332 ( .A(n_220), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_220), .B(n_292), .Y(n_382) );
INVx5_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g272 ( .A(n_221), .B(n_246), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_221), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g299 ( .A(n_221), .B(n_230), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_221), .B(n_346), .Y(n_387) );
OR2x2_ASAP7_75t_L g403 ( .A(n_221), .B(n_347), .Y(n_403) );
AND2x2_ASAP7_75t_SL g410 ( .A(n_221), .B(n_364), .Y(n_410) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_221), .Y(n_417) );
OR2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_228), .Y(n_221) );
AND2x2_ASAP7_75t_L g271 ( .A(n_229), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g321 ( .A(n_229), .B(n_244), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_229), .B(n_246), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_229), .B(n_283), .Y(n_405) );
INVx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_230), .B(n_246), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_230), .B(n_244), .Y(n_293) );
OR2x2_ASAP7_75t_L g347 ( .A(n_230), .B(n_244), .Y(n_347) );
AND2x2_ASAP7_75t_L g364 ( .A(n_230), .B(n_243), .Y(n_364) );
INVxp67_ASAP7_75t_L g386 ( .A(n_230), .Y(n_386) );
AND2x2_ASAP7_75t_L g413 ( .A(n_230), .B(n_283), .Y(n_413) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_230), .Y(n_420) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_240), .Y(n_230) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_231), .A2(n_475), .B(n_482), .Y(n_474) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_231), .A2(n_498), .B(n_504), .Y(n_497) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_231), .A2(n_518), .B(n_525), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_236), .A2(n_263), .B(n_264), .C(n_265), .Y(n_262) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_237), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_237), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_245), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_243), .B(n_294), .Y(n_367) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g283 ( .A(n_244), .B(n_246), .Y(n_283) );
OR2x2_ASAP7_75t_L g350 ( .A(n_244), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g294 ( .A(n_245), .Y(n_294) );
OR2x2_ASAP7_75t_L g355 ( .A(n_245), .B(n_347), .Y(n_355) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g254 ( .A(n_249), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_249), .B(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g255 ( .A(n_250), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_250), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_250), .B(n_257), .Y(n_290) );
INVx2_ASAP7_75t_L g335 ( .A(n_250), .Y(n_335) );
AND2x2_ASAP7_75t_L g348 ( .A(n_250), .B(n_288), .Y(n_348) );
AND2x2_ASAP7_75t_L g373 ( .A(n_250), .B(n_297), .Y(n_373) );
INVx1_ASAP7_75t_L g325 ( .A(n_255), .Y(n_325) );
INVx2_ASAP7_75t_SL g312 ( .A(n_256), .Y(n_312) );
INVx1_ASAP7_75t_L g315 ( .A(n_257), .Y(n_315) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_258), .Y(n_278) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx2_ASAP7_75t_L g376 ( .A(n_259), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_267), .Y(n_260) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx3_ASAP7_75t_L g481 ( .A(n_266), .Y(n_481) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g345 ( .A(n_272), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g351 ( .A(n_272), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_272), .A2(n_354), .B1(n_356), .B2(n_361), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_272), .B(n_364), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_273), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g307 ( .A(n_274), .Y(n_307) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
OR2x2_ASAP7_75t_L g289 ( .A(n_276), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_276), .B(n_280), .Y(n_340) );
AND2x2_ASAP7_75t_L g363 ( .A(n_276), .B(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g339 ( .A(n_278), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B(n_286), .C(n_300), .Y(n_279) );
INVx1_ASAP7_75t_L g303 ( .A(n_280), .Y(n_303) );
OAI221xp5_ASAP7_75t_SL g411 ( .A1(n_280), .A2(n_412), .B1(n_414), .B2(n_415), .C(n_418), .Y(n_411) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g430 ( .A(n_283), .Y(n_430) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g379 ( .A(n_285), .B(n_318), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_289), .B(n_291), .C(n_295), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OAI32xp33_ASAP7_75t_L g404 ( .A1(n_293), .A2(n_294), .A3(n_357), .B1(n_394), .B2(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
AND2x2_ASAP7_75t_L g436 ( .A(n_296), .B(n_335), .Y(n_436) );
AND2x2_ASAP7_75t_L g383 ( .A(n_297), .B(n_335), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_297), .B(n_305), .Y(n_401) );
AOI31xp33_ASAP7_75t_SL g300 ( .A1(n_301), .A2(n_303), .A3(n_304), .B(n_306), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_302), .B(n_314), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_302), .B(n_312), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_302), .A2(n_332), .B1(n_422), .B2(n_425), .C(n_427), .Y(n_421) );
CKINVDCx16_ASAP7_75t_R g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
AND2x2_ASAP7_75t_L g327 ( .A(n_307), .B(n_328), .Y(n_327) );
AOI222xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_316), .B1(n_319), .B2(n_322), .C1(n_324), .C2(n_325), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g392 ( .A(n_311), .Y(n_392) );
INVx1_ASAP7_75t_L g414 ( .A(n_314), .Y(n_414) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_317), .A2(n_428), .B1(n_430), .B2(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g333 ( .A(n_318), .Y(n_333) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .B1(n_332), .B2(n_334), .C(n_337), .Y(n_326) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g371 ( .A(n_329), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g423 ( .A(n_329), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g398 ( .A(n_334), .Y(n_398) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g362 ( .A(n_335), .Y(n_362) );
INVx1_ASAP7_75t_L g344 ( .A(n_336), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_339), .B(n_426), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_345), .B1(n_348), .B2(n_349), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g435 ( .A(n_348), .Y(n_435) );
INVxp33_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_350), .B(n_394), .Y(n_393) );
OAI32xp33_ASAP7_75t_L g384 ( .A1(n_351), .A2(n_385), .A3(n_386), .B1(n_387), .B2(n_388), .Y(n_384) );
NAND4xp25_ASAP7_75t_L g352 ( .A(n_353), .B(n_365), .C(n_377), .D(n_389), .Y(n_352) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
NAND2xp33_ASAP7_75t_SL g356 ( .A(n_357), .B(n_358), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_360), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
CKINVDCx16_ASAP7_75t_R g370 ( .A(n_371), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_374), .A2(n_390), .B1(n_407), .B2(n_410), .C(n_411), .Y(n_406) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g425 ( .A(n_376), .B(n_426), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B1(n_381), .B2(n_383), .C(n_384), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_386), .B(n_417), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B(n_393), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND4xp25_ASAP7_75t_L g395 ( .A(n_396), .B(n_406), .C(n_421), .D(n_432), .Y(n_395) );
O2A1O1Ixp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .B(n_402), .C(n_404), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g437 ( .A(n_424), .Y(n_437) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_436), .B(n_437), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_438), .A2(n_449), .B1(n_451), .B2(n_454), .Y(n_448) );
NOR2xp33_ASAP7_75t_SL g444 ( .A(n_439), .B(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR2x2_ASAP7_75t_L g740 ( .A(n_441), .B(n_453), .Y(n_740) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g452 ( .A(n_442), .B(n_453), .Y(n_452) );
OAI21xp5_ASAP7_75t_SL g446 ( .A1(n_444), .A2(n_447), .B(n_742), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g734 ( .A(n_450), .Y(n_734) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx6_ASAP7_75t_L g735 ( .A(n_452), .Y(n_735) );
INVx3_ASAP7_75t_L g736 ( .A(n_454), .Y(n_736) );
AND2x2_ASAP7_75t_SL g454 ( .A(n_455), .B(n_685), .Y(n_454) );
NOR4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_622), .C(n_656), .D(n_672), .Y(n_455) );
NAND4xp25_ASAP7_75t_SL g456 ( .A(n_457), .B(n_551), .C(n_586), .D(n_602), .Y(n_456) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_492), .B1(n_526), .B2(n_539), .C1(n_544), .C2(n_550), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI31xp33_ASAP7_75t_L g718 ( .A1(n_459), .A2(n_719), .A3(n_720), .B(n_722), .Y(n_718) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .Y(n_459) );
AND2x2_ASAP7_75t_L g693 ( .A(n_460), .B(n_473), .Y(n_693) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_SL g543 ( .A(n_461), .Y(n_543) );
AND2x2_ASAP7_75t_L g550 ( .A(n_461), .B(n_483), .Y(n_550) );
AND2x2_ASAP7_75t_L g607 ( .A(n_461), .B(n_474), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_471), .B(n_637), .Y(n_636) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_472), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_472), .B(n_554), .Y(n_597) );
AND2x2_ASAP7_75t_L g690 ( .A(n_472), .B(n_630), .Y(n_690) );
OAI321xp33_ASAP7_75t_L g724 ( .A1(n_472), .A2(n_543), .A3(n_697), .B1(n_725), .B2(n_727), .C(n_728), .Y(n_724) );
NAND4xp25_ASAP7_75t_L g728 ( .A(n_472), .B(n_529), .C(n_637), .D(n_729), .Y(n_728) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_483), .Y(n_472) );
AND2x2_ASAP7_75t_L g592 ( .A(n_473), .B(n_541), .Y(n_592) );
AND2x2_ASAP7_75t_L g611 ( .A(n_473), .B(n_543), .Y(n_611) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g542 ( .A(n_474), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g567 ( .A(n_474), .B(n_483), .Y(n_567) );
AND2x2_ASAP7_75t_L g653 ( .A(n_474), .B(n_541), .Y(n_653) );
INVx3_ASAP7_75t_SL g541 ( .A(n_483), .Y(n_541) );
AND2x2_ASAP7_75t_L g585 ( .A(n_483), .B(n_572), .Y(n_585) );
OR2x2_ASAP7_75t_L g618 ( .A(n_483), .B(n_543), .Y(n_618) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_483), .Y(n_625) );
AND2x2_ASAP7_75t_L g654 ( .A(n_483), .B(n_542), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_483), .B(n_627), .Y(n_669) );
AND2x2_ASAP7_75t_L g701 ( .A(n_483), .B(n_693), .Y(n_701) );
AND2x2_ASAP7_75t_L g710 ( .A(n_483), .B(n_555), .Y(n_710) );
OR2x6_ASAP7_75t_L g483 ( .A(n_484), .B(n_490), .Y(n_483) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_505), .Y(n_493) );
INVx1_ASAP7_75t_SL g678 ( .A(n_494), .Y(n_678) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g546 ( .A(n_495), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g528 ( .A(n_496), .B(n_507), .Y(n_528) );
AND2x2_ASAP7_75t_L g614 ( .A(n_496), .B(n_530), .Y(n_614) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g584 ( .A(n_497), .B(n_517), .Y(n_584) );
OR2x2_ASAP7_75t_L g595 ( .A(n_497), .B(n_530), .Y(n_595) );
AND2x2_ASAP7_75t_L g621 ( .A(n_497), .B(n_530), .Y(n_621) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_497), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_505), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_505), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g594 ( .A(n_506), .B(n_595), .Y(n_594) );
AOI322xp5_ASAP7_75t_L g680 ( .A1(n_506), .A2(n_584), .A3(n_590), .B1(n_621), .B2(n_671), .C1(n_681), .C2(n_683), .Y(n_680) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_517), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_507), .B(n_529), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_507), .B(n_530), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_507), .B(n_547), .Y(n_601) );
AND2x2_ASAP7_75t_L g655 ( .A(n_507), .B(n_621), .Y(n_655) );
INVx1_ASAP7_75t_L g659 ( .A(n_507), .Y(n_659) );
AND2x2_ASAP7_75t_L g671 ( .A(n_507), .B(n_517), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_507), .B(n_546), .Y(n_703) );
INVx4_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g568 ( .A(n_508), .B(n_517), .Y(n_568) );
BUFx3_ASAP7_75t_L g582 ( .A(n_508), .Y(n_582) );
AND3x2_ASAP7_75t_L g664 ( .A(n_508), .B(n_644), .C(n_665), .Y(n_664) );
NAND3xp33_ASAP7_75t_L g527 ( .A(n_517), .B(n_528), .C(n_529), .Y(n_527) );
INVx1_ASAP7_75t_SL g547 ( .A(n_517), .Y(n_547) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_517), .Y(n_649) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g643 ( .A(n_528), .B(n_644), .Y(n_643) );
INVxp67_ASAP7_75t_L g650 ( .A(n_528), .Y(n_650) );
AND2x2_ASAP7_75t_L g688 ( .A(n_529), .B(n_666), .Y(n_688) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx3_ASAP7_75t_L g569 ( .A(n_530), .Y(n_569) );
AND2x2_ASAP7_75t_L g644 ( .A(n_530), .B(n_547), .Y(n_644) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
OR2x2_ASAP7_75t_L g588 ( .A(n_541), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g707 ( .A(n_541), .B(n_607), .Y(n_707) );
AND2x2_ASAP7_75t_L g721 ( .A(n_541), .B(n_543), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_542), .B(n_555), .Y(n_662) );
AND2x2_ASAP7_75t_L g709 ( .A(n_542), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g572 ( .A(n_543), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g589 ( .A(n_543), .B(n_555), .Y(n_589) );
INVx1_ASAP7_75t_L g599 ( .A(n_543), .Y(n_599) );
AND2x2_ASAP7_75t_L g630 ( .A(n_543), .B(n_555), .Y(n_630) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_545), .A2(n_673), .B1(n_677), .B2(n_679), .C(n_680), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_546), .B(n_548), .Y(n_545) );
AND2x2_ASAP7_75t_L g576 ( .A(n_546), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_549), .B(n_583), .Y(n_726) );
AOI322xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_568), .A3(n_569), .B1(n_570), .B2(n_576), .C1(n_578), .C2(n_585), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_567), .Y(n_553) );
NAND2x1p5_ASAP7_75t_L g606 ( .A(n_554), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_554), .B(n_617), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_554), .A2(n_567), .B(n_641), .C(n_642), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_554), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_554), .B(n_611), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_554), .B(n_693), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_554), .B(n_721), .Y(n_720) );
BUFx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_555), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_555), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g682 ( .A(n_555), .B(n_569), .Y(n_682) );
OA21x2_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_559), .B(n_566), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_557), .A2(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g574 ( .A(n_559), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_566), .Y(n_575) );
INVx1_ASAP7_75t_L g657 ( .A(n_567), .Y(n_657) );
OAI31xp33_ASAP7_75t_L g667 ( .A1(n_567), .A2(n_592), .A3(n_668), .B(n_670), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_567), .B(n_573), .Y(n_719) );
INVx1_ASAP7_75t_SL g580 ( .A(n_568), .Y(n_580) );
AND2x2_ASAP7_75t_L g613 ( .A(n_568), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g694 ( .A(n_568), .B(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g579 ( .A(n_569), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g604 ( .A(n_569), .Y(n_604) );
AND2x2_ASAP7_75t_L g631 ( .A(n_569), .B(n_584), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_569), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g723 ( .A(n_569), .B(n_671), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_571), .B(n_641), .Y(n_714) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g610 ( .A(n_573), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g628 ( .A(n_573), .Y(n_628) );
NAND2xp33_ASAP7_75t_SL g578 ( .A(n_579), .B(n_581), .Y(n_578) );
OAI211xp5_ASAP7_75t_SL g622 ( .A1(n_580), .A2(n_623), .B(n_629), .C(n_645), .Y(n_622) );
OR2x2_ASAP7_75t_L g697 ( .A(n_580), .B(n_678), .Y(n_697) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
CKINVDCx16_ASAP7_75t_R g634 ( .A(n_582), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_582), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g603 ( .A(n_584), .B(n_604), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_590), .B(n_593), .C(n_596), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_SL g637 ( .A(n_589), .Y(n_637) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_592), .B(n_630), .Y(n_635) );
INVx1_ASAP7_75t_L g641 ( .A(n_592), .Y(n_641) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g600 ( .A(n_595), .B(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g633 ( .A(n_595), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g695 ( .A(n_595), .Y(n_695) );
AOI21xp33_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_598), .B(n_600), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_598), .A2(n_609), .B(n_612), .Y(n_608) );
AOI211xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_605), .B(n_608), .C(n_615), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_603), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_606), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_SL g619 ( .A(n_607), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_609), .A2(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_614), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g639 ( .A(n_614), .Y(n_639) );
AOI21xp33_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_619), .B(n_620), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g670 ( .A(n_621), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_627), .B(n_653), .Y(n_679) );
AND2x2_ASAP7_75t_L g692 ( .A(n_627), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g706 ( .A(n_627), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g716 ( .A(n_627), .B(n_654), .Y(n_716) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AOI211xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B(n_632), .C(n_640), .Y(n_629) );
INVx1_ASAP7_75t_L g676 ( .A(n_630), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B1(n_636), .B2(n_638), .Y(n_632) );
OR2x2_ASAP7_75t_L g638 ( .A(n_634), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_634), .B(n_695), .Y(n_717) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g711 ( .A(n_644), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_651), .B1(n_654), .B2(n_655), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g729 ( .A(n_649), .Y(n_729) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g675 ( .A(n_653), .Y(n_675) );
OAI211xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_658), .B(n_660), .C(n_667), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx2_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_675), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NOR5xp2_ASAP7_75t_L g685 ( .A(n_686), .B(n_704), .C(n_712), .D(n_718), .E(n_724), .Y(n_685) );
OAI211xp5_ASAP7_75t_SL g686 ( .A1(n_687), .A2(n_689), .B(n_691), .C(n_698), .Y(n_686) );
INVxp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_694), .B(n_696), .Y(n_691) );
OAI21xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_701), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_708), .B(n_711), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g727 ( .A(n_707), .Y(n_727) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B(n_717), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
endmodule