module fake_ariane_1897_n_1859 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1859);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1859;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_699;
wire n_590;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_115),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_4),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_164),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_47),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_110),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_53),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_66),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_34),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_0),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_88),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_12),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_24),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_116),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_89),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_37),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_28),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_53),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_127),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_100),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_15),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_32),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_153),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_99),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_135),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_142),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_65),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_1),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_155),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_123),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_30),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_130),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_60),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_57),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_17),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_45),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_106),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_23),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_46),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_126),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_77),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_17),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_14),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_97),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_163),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_48),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_78),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_52),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_40),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_139),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_42),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_72),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_96),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_5),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_29),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_51),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_49),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_64),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_6),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_145),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_144),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_168),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_154),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_54),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_75),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_47),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_55),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_14),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_90),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_26),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_105),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_147),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_107),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_160),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_80),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_6),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_3),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_67),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_63),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_62),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_12),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_82),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_43),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_43),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_0),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_40),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_69),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_29),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_143),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_133),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_117),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_23),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_124),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_20),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_41),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_104),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_31),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_119),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_30),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_50),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_86),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_38),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_84),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_27),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_61),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_122),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_148),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_70),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_114),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_132),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_131),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_151),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_125),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_111),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_48),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_118),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_169),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_92),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_73),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_16),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_165),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_5),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_22),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_35),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_39),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_11),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_59),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_102),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_24),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_79),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_162),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_9),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_20),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_166),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_28),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_46),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_2),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_18),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_10),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_45),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_10),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_19),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_8),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_44),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_42),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_52),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_108),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_58),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_121),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_50),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_113),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_26),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_101),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_161),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_2),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_35),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_120),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_16),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_41),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_27),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_11),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_176),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_245),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_236),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_236),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_204),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_236),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_335),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_269),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_307),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_174),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_318),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_204),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_174),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_180),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_175),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_175),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_226),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_195),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_216),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_177),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_226),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_308),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_171),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_259),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_255),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_259),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_173),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_171),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_320),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_178),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_186),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_178),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_186),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_185),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_185),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_199),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_281),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_177),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_199),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_182),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g387 ( 
.A(n_214),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_214),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_182),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_170),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_281),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_222),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_222),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_173),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_234),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_234),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_264),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_264),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_337),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_265),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_265),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_267),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_337),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_267),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_338),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_338),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_188),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_193),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_196),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_273),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_183),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_273),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_274),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_200),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_274),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_317),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_317),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_183),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_194),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_194),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_205),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_206),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_205),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_220),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_334),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_209),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_220),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_228),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_373),
.Y(n_429)
);

NAND2x1p5_ASAP7_75t_L g430 ( 
.A(n_355),
.B(n_254),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_411),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_368),
.B(n_228),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_355),
.B(n_241),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_373),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_360),
.A2(n_189),
.B1(n_304),
.B2(n_314),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_424),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_409),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_373),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_386),
.B(n_389),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_377),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_377),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_386),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_368),
.B(n_238),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_359),
.B(n_211),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_424),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_390),
.B(n_241),
.Y(n_447)
);

NOR2x1_ASAP7_75t_L g448 ( 
.A(n_389),
.B(n_313),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_L g450 ( 
.A(n_345),
.B(n_221),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_342),
.A2(n_262),
.B1(n_221),
.B2(n_213),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_373),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_361),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_361),
.B(n_262),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_341),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_362),
.Y(n_456)
);

OA21x2_ASAP7_75t_L g457 ( 
.A1(n_362),
.A2(n_246),
.B(n_244),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_394),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_372),
.B(n_244),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_394),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_366),
.B(n_246),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_407),
.B(n_212),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_366),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_384),
.B(n_253),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_418),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_418),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_419),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_419),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_420),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_356),
.A2(n_334),
.B1(n_339),
.B2(n_217),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_420),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_364),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_421),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_368),
.B(n_238),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_349),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_344),
.B(n_271),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_345),
.B(n_253),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_423),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_423),
.B(n_427),
.Y(n_486)
);

AND2x2_ASAP7_75t_SL g487 ( 
.A(n_427),
.B(n_211),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_374),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_343),
.B(n_271),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_376),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_378),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_381),
.Y(n_492)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_369),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_385),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_383),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_352),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_392),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_399),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_393),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_396),
.B(n_215),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_346),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_395),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_397),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_493),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_475),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_475),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_475),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_484),
.B(n_407),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_475),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_475),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_475),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_448),
.B(n_261),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_502),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_478),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_478),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_471),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_435),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_471),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_471),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_467),
.B(n_350),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_447),
.B(n_408),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_478),
.Y(n_523)
);

NAND3xp33_ASAP7_75t_L g524 ( 
.A(n_449),
.B(n_363),
.C(n_358),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_477),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_478),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_493),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_443),
.B(n_493),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_443),
.B(n_358),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_455),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_502),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_477),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_451),
.A2(n_363),
.B1(n_367),
.B2(n_370),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_477),
.Y(n_534)
);

AND3x2_ASAP7_75t_L g535 ( 
.A(n_467),
.B(n_357),
.C(n_425),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_485),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_485),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_485),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_464),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_464),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_449),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_464),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_443),
.B(n_367),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_464),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_453),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_453),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_430),
.B(n_440),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_456),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_457),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_456),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_465),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_429),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_465),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_469),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_469),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_488),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_430),
.B(n_408),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_430),
.B(n_414),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_479),
.B(n_365),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_493),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_488),
.Y(n_561)
);

AND2x2_ASAP7_75t_SL g562 ( 
.A(n_487),
.B(n_252),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_472),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_493),
.B(n_370),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_472),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_429),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_429),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_502),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_487),
.B(n_347),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_439),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_487),
.B(n_348),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_439),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_440),
.B(n_351),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_439),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_458),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_458),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_440),
.B(n_414),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_458),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_473),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_440),
.B(n_422),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_474),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_459),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_459),
.Y(n_583)
);

OAI21xp33_ASAP7_75t_SL g584 ( 
.A1(n_486),
.A2(n_382),
.B(n_380),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_488),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_474),
.B(n_422),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_459),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_457),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_468),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_451),
.A2(n_463),
.B1(n_476),
.B2(n_403),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_448),
.B(n_398),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_468),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_428),
.Y(n_593)
);

BUFx6f_ASAP7_75t_SL g594 ( 
.A(n_454),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_480),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_480),
.B(n_426),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_454),
.B(n_400),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_431),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_431),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_434),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_434),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_454),
.B(n_353),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_437),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_428),
.B(n_401),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_468),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_437),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_446),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_470),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_470),
.Y(n_609)
);

BUFx6f_ASAP7_75t_SL g610 ( 
.A(n_454),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_483),
.B(n_402),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_499),
.B(n_399),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_499),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_446),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_432),
.B(n_444),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_501),
.B(n_403),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_483),
.Y(n_617)
);

NOR3xp33_ASAP7_75t_L g618 ( 
.A(n_476),
.B(n_406),
.C(n_405),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_470),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_488),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_457),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_457),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_450),
.B(n_405),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_501),
.B(n_406),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_486),
.B(n_404),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_488),
.Y(n_626)
);

NAND3xp33_ASAP7_75t_L g627 ( 
.A(n_488),
.B(n_270),
.C(n_261),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_457),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_492),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_492),
.Y(n_630)
);

AND2x2_ASAP7_75t_SL g631 ( 
.A(n_433),
.B(n_252),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_490),
.B(n_410),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_441),
.B(n_357),
.Y(n_633)
);

OAI22xp33_ASAP7_75t_L g634 ( 
.A1(n_441),
.A2(n_496),
.B1(n_442),
.B2(n_460),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_492),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_492),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_490),
.B(n_412),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_491),
.B(n_413),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_491),
.B(n_415),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_492),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_492),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_489),
.A2(n_312),
.B1(n_321),
.B2(n_319),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_494),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_494),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_442),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_496),
.B(n_379),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_494),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_433),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_435),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_435),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_462),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_SL g652 ( 
.A(n_462),
.B(n_391),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_466),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_435),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_432),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_517),
.Y(n_656)
);

A2O1A1Ixp33_ASAP7_75t_L g657 ( 
.A1(n_648),
.A2(n_466),
.B(n_503),
.C(n_500),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_648),
.B(n_495),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_613),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_651),
.B(n_653),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_623),
.B(n_524),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_517),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_613),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_645),
.B(n_438),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_651),
.B(n_495),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_645),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_564),
.B(n_498),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_653),
.B(n_504),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_591),
.B(n_504),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_591),
.B(n_444),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_562),
.B(n_270),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_521),
.B(n_438),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_559),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_541),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_562),
.A2(n_311),
.B1(n_276),
.B2(n_230),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_591),
.B(n_481),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_593),
.B(n_482),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_591),
.B(n_481),
.Y(n_678)
);

INVx8_ASAP7_75t_L g679 ( 
.A(n_594),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_580),
.B(n_489),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_505),
.B(n_489),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_631),
.A2(n_445),
.B1(n_289),
.B2(n_272),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_505),
.B(n_489),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_519),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_559),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_631),
.B(n_272),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_SL g687 ( 
.A(n_594),
.B(n_354),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_593),
.A2(n_436),
.B1(n_445),
.B2(n_321),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_541),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_521),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_527),
.B(n_285),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_535),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_527),
.B(n_285),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_527),
.B(n_516),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_560),
.B(n_445),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_529),
.B(n_225),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_545),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_520),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_527),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_516),
.B(n_286),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_514),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_545),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_617),
.B(n_445),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_520),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_546),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_525),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_543),
.B(n_227),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_586),
.A2(n_278),
.B1(n_256),
.B2(n_279),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_526),
.B(n_549),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_509),
.B(n_233),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_646),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_604),
.B(n_497),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_526),
.B(n_286),
.Y(n_713)
);

AO221x1_ASAP7_75t_L g714 ( 
.A1(n_533),
.A2(n_436),
.B1(n_300),
.B2(n_309),
.C(n_289),
.Y(n_714)
);

INVx8_ASAP7_75t_L g715 ( 
.A(n_610),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_514),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_530),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_525),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_655),
.B(n_445),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_596),
.B(n_235),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_655),
.B(n_445),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_532),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_597),
.B(n_445),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_549),
.B(n_290),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_532),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_547),
.B(n_243),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_546),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_537),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_597),
.B(n_445),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_548),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_621),
.A2(n_293),
.B(n_290),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_514),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_530),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_515),
.A2(n_277),
.B(n_215),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_SL g735 ( 
.A(n_522),
.B(n_247),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_537),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_534),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_534),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_536),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_536),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_604),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_531),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_597),
.B(n_327),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_597),
.B(n_615),
.Y(n_744)
);

AND2x2_ASAP7_75t_SL g745 ( 
.A(n_618),
.B(n_569),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_584),
.A2(n_319),
.B(n_315),
.C(n_283),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_507),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_610),
.A2(n_309),
.B1(n_293),
.B2(n_297),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_633),
.B(n_371),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_612),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_538),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_615),
.B(n_283),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_625),
.B(n_312),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_611),
.B(n_315),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_538),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_513),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_548),
.B(n_297),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_557),
.A2(n_300),
.B1(n_310),
.B2(n_328),
.Y(n_758)
);

OA22x2_ASAP7_75t_L g759 ( 
.A1(n_558),
.A2(n_577),
.B1(n_602),
.B2(n_573),
.Y(n_759)
);

NOR2x1p5_ASAP7_75t_L g760 ( 
.A(n_524),
.B(n_416),
.Y(n_760)
);

AND2x2_ASAP7_75t_SL g761 ( 
.A(n_571),
.B(n_258),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_507),
.B(n_249),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_550),
.B(n_310),
.Y(n_763)
);

OAI221xp5_ASAP7_75t_L g764 ( 
.A1(n_584),
.A2(n_263),
.B1(n_299),
.B2(n_340),
.C(n_302),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_550),
.B(n_328),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_513),
.A2(n_336),
.B1(n_277),
.B2(n_207),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_531),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_SL g768 ( 
.A1(n_634),
.A2(n_375),
.B1(n_305),
.B2(n_329),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_551),
.B(n_336),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_551),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_643),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_553),
.B(n_417),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_553),
.B(n_260),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_531),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_549),
.B(n_258),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_554),
.B(n_294),
.Y(n_776)
);

NAND2xp33_ASAP7_75t_L g777 ( 
.A(n_507),
.B(n_303),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_513),
.A2(n_284),
.B1(n_322),
.B2(n_325),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_554),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_644),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_568),
.B(n_316),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_555),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_568),
.B(n_323),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_513),
.A2(n_284),
.B1(n_331),
.B2(n_324),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_555),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_568),
.B(n_616),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_563),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_513),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_549),
.B(n_173),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_563),
.A2(n_3),
.B(n_4),
.C(n_7),
.Y(n_790)
);

NAND3x1_ASAP7_75t_L g791 ( 
.A(n_632),
.B(n_7),
.C(n_8),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_565),
.B(n_172),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_515),
.A2(n_461),
.B(n_452),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_513),
.A2(n_173),
.B1(n_268),
.B2(n_282),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_644),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_647),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_565),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_629),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_579),
.B(n_179),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_588),
.B(n_173),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_513),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_579),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_581),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_647),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_523),
.B(n_184),
.C(n_333),
.Y(n_805)
);

INVx8_ASAP7_75t_L g806 ( 
.A(n_507),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_624),
.B(n_9),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_528),
.B(n_523),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_588),
.B(n_268),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_629),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_652),
.B(n_13),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_629),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_581),
.B(n_181),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_637),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_595),
.B(n_13),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_595),
.B(n_187),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_598),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_588),
.B(n_268),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_598),
.B(n_190),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_663),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_741),
.B(n_638),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_664),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_714),
.A2(n_642),
.B1(n_599),
.B2(n_600),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_R g824 ( 
.A(n_687),
.B(n_556),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_817),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_656),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_666),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_659),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_690),
.B(n_639),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_656),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_701),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_711),
.B(n_599),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_817),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_733),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_660),
.B(n_667),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_677),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_667),
.B(n_600),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_806),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_674),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_672),
.B(n_601),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_712),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_814),
.B(n_744),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_689),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_697),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_679),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_806),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_679),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_720),
.A2(n_601),
.B1(n_607),
.B2(n_606),
.Y(n_848)
);

OR2x2_ASAP7_75t_SL g849 ( 
.A(n_685),
.B(n_749),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_679),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_702),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_715),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_705),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_727),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_709),
.A2(n_588),
.B(n_621),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_730),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_715),
.Y(n_857)
);

INVx5_ASAP7_75t_L g858 ( 
.A(n_715),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_770),
.B(n_603),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_662),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_662),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_717),
.B(n_603),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_806),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_692),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_779),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_670),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_782),
.B(n_606),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_785),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_671),
.A2(n_614),
.B1(n_607),
.B2(n_627),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_720),
.A2(n_614),
.B1(n_556),
.B2(n_585),
.Y(n_870)
);

CKINVDCx8_ASAP7_75t_R g871 ( 
.A(n_710),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_787),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_671),
.A2(n_627),
.B1(n_628),
.B2(n_622),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_797),
.B(n_622),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_745),
.A2(n_561),
.B1(n_585),
.B2(n_556),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_761),
.A2(n_628),
.B1(n_630),
.B2(n_626),
.Y(n_876)
);

AND3x2_ASAP7_75t_SL g877 ( 
.A(n_768),
.B(n_620),
.C(n_640),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_760),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_781),
.B(n_783),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_802),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_684),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_747),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_803),
.Y(n_883)
);

OR2x6_ASAP7_75t_L g884 ( 
.A(n_673),
.B(n_630),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_737),
.Y(n_885)
);

OAI21xp33_ASAP7_75t_SL g886 ( 
.A1(n_731),
.A2(n_506),
.B(n_508),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_658),
.B(n_510),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_752),
.B(n_539),
.Y(n_888)
);

AO22x1_ASAP7_75t_L g889 ( 
.A1(n_710),
.A2(n_242),
.B1(n_295),
.B2(n_292),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_737),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_767),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_676),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_750),
.B(n_561),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_665),
.B(n_510),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_668),
.B(n_510),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_781),
.B(n_511),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_657),
.B(n_506),
.Y(n_897)
);

NOR2x2_ASAP7_75t_L g898 ( 
.A(n_675),
.B(n_539),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_696),
.A2(n_585),
.B1(n_561),
.B2(n_636),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_684),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_767),
.B(n_678),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_657),
.B(n_508),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_696),
.B(n_512),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_738),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_807),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_815),
.A2(n_544),
.B1(n_542),
.B2(n_540),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_771),
.B(n_780),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_738),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_739),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_739),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_761),
.A2(n_620),
.B1(n_626),
.B2(n_641),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_698),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_716),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_759),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_SL g915 ( 
.A1(n_707),
.A2(n_649),
.B(n_540),
.C(n_542),
.Y(n_915)
);

OAI221xp5_ASAP7_75t_L g916 ( 
.A1(n_746),
.A2(n_635),
.B1(n_640),
.B2(n_641),
.C(n_544),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_707),
.A2(n_511),
.B1(n_291),
.B2(n_288),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_680),
.A2(n_511),
.B1(n_296),
.B2(n_287),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_SL g919 ( 
.A(n_699),
.B(n_649),
.Y(n_919)
);

NOR2x2_ASAP7_75t_L g920 ( 
.A(n_687),
.B(n_650),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_743),
.B(n_669),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_754),
.B(n_552),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_780),
.B(n_552),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_698),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_740),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_726),
.B(n_649),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_680),
.A2(n_203),
.B1(n_202),
.B2(n_201),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_716),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_704),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_704),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_759),
.Y(n_931)
);

AND2x6_ASAP7_75t_L g932 ( 
.A(n_742),
.B(n_566),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_795),
.B(n_566),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_783),
.B(n_654),
.Y(n_934)
);

NAND2x1p5_ASAP7_75t_L g935 ( 
.A(n_732),
.B(n_649),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_747),
.Y(n_936)
);

NAND2xp33_ASAP7_75t_L g937 ( 
.A(n_747),
.B(n_654),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_795),
.B(n_567),
.Y(n_938)
);

OR2x6_ASAP7_75t_L g939 ( 
.A(n_756),
.B(n_567),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_735),
.Y(n_940)
);

NOR2x1_ASAP7_75t_R g941 ( 
.A(n_773),
.B(n_191),
.Y(n_941)
);

AND3x1_ASAP7_75t_SL g942 ( 
.A(n_764),
.B(n_15),
.C(n_18),
.Y(n_942)
);

INVx5_ASAP7_75t_L g943 ( 
.A(n_747),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_776),
.B(n_570),
.Y(n_944)
);

AND2x6_ASAP7_75t_L g945 ( 
.A(n_742),
.B(n_774),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_740),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_732),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_708),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_788),
.B(n_570),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_SL g950 ( 
.A1(n_688),
.A2(n_208),
.B1(n_332),
.B2(n_330),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_706),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_706),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_751),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_812),
.Y(n_954)
);

BUFx4f_ASAP7_75t_L g955 ( 
.A(n_811),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_726),
.B(n_572),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_709),
.A2(n_650),
.B(n_582),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_812),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_786),
.B(n_807),
.Y(n_959)
);

OR2x6_ASAP7_75t_L g960 ( 
.A(n_801),
.B(n_572),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_723),
.B(n_574),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_718),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_796),
.B(n_574),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_786),
.A2(n_784),
.B1(n_778),
.B2(n_686),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_815),
.A2(n_589),
.B1(n_619),
.B2(n_609),
.Y(n_965)
);

INVx5_ASAP7_75t_L g966 ( 
.A(n_774),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_686),
.A2(n_589),
.B1(n_619),
.B2(n_609),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_796),
.B(n_804),
.Y(n_968)
);

NAND2xp33_ASAP7_75t_L g969 ( 
.A(n_694),
.B(n_654),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_804),
.B(n_575),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_753),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_718),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_766),
.A2(n_266),
.B1(n_197),
.B2(n_198),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_751),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_722),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_755),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_755),
.B(n_575),
.Y(n_977)
);

AO21x2_ASAP7_75t_L g978 ( 
.A1(n_789),
.A2(n_608),
.B(n_605),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_682),
.A2(n_608),
.B1(n_605),
.B2(n_592),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_808),
.B(n_576),
.Y(n_980)
);

NOR2xp67_ASAP7_75t_L g981 ( 
.A(n_748),
.B(n_578),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_772),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_729),
.B(n_578),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_722),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_746),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_798),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_725),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_725),
.Y(n_988)
);

NAND2x1p5_ASAP7_75t_L g989 ( 
.A(n_810),
.B(n_518),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_758),
.B(n_792),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_681),
.Y(n_991)
);

INVx5_ASAP7_75t_L g992 ( 
.A(n_728),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_728),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_736),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_808),
.B(n_583),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_838),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_835),
.A2(n_809),
.B(n_818),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_858),
.B(n_683),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_826),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_R g1000 ( 
.A(n_824),
.B(n_703),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_839),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_830),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_860),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_840),
.B(n_757),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_835),
.B(n_763),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_861),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_R g1007 ( 
.A(n_871),
.B(n_762),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_879),
.A2(n_790),
.B(n_816),
.C(n_813),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_828),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_837),
.A2(n_769),
.B1(n_765),
.B2(n_799),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_827),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_820),
.B(n_691),
.Y(n_1012)
);

OR2x6_ASAP7_75t_L g1013 ( 
.A(n_884),
.B(n_857),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_822),
.B(n_700),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_837),
.A2(n_700),
.B1(n_713),
.B2(n_724),
.Y(n_1015)
);

O2A1O1Ixp5_ASAP7_75t_L g1016 ( 
.A1(n_990),
.A2(n_818),
.B(n_809),
.C(n_789),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_834),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_832),
.B(n_819),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_843),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_R g1020 ( 
.A(n_858),
.B(n_777),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_858),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_L g1022 ( 
.A(n_948),
.B(n_805),
.C(n_713),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_866),
.B(n_736),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_844),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_858),
.B(n_694),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_905),
.B(n_691),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_827),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_959),
.A2(n_724),
.B(n_734),
.C(n_693),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_866),
.B(n_693),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_903),
.A2(n_800),
.B(n_775),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_980),
.A2(n_995),
.B(n_874),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_892),
.B(n_921),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_862),
.A2(n_721),
.B(n_719),
.C(n_800),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_980),
.A2(n_775),
.B(n_793),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_851),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_943),
.B(n_518),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_892),
.B(n_583),
.Y(n_1037)
);

INVx5_ASAP7_75t_L g1038 ( 
.A(n_838),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_841),
.B(n_587),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_955),
.A2(n_794),
.B1(n_695),
.B2(n_587),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_982),
.B(n_592),
.Y(n_1041)
);

OAI21xp33_ASAP7_75t_L g1042 ( 
.A1(n_927),
.A2(n_240),
.B(n_326),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_836),
.Y(n_1043)
);

INVx8_ASAP7_75t_L g1044 ( 
.A(n_945),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_829),
.B(n_955),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_859),
.A2(n_791),
.B1(n_518),
.B2(n_298),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_R g1047 ( 
.A(n_845),
.B(n_210),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_995),
.A2(n_874),
.B(n_937),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_884),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_838),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_846),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_881),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_853),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_926),
.A2(n_248),
.B(n_218),
.C(n_219),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_907),
.B(n_968),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_859),
.A2(n_192),
.B1(n_223),
.B2(n_224),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_846),
.B(n_257),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_842),
.B(n_229),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_907),
.B(n_19),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_847),
.B(n_21),
.Y(n_1060)
);

OA21x2_ASAP7_75t_L g1061 ( 
.A1(n_897),
.A2(n_231),
.B(n_232),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_SL g1062 ( 
.A(n_941),
.B(n_275),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_854),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_900),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_887),
.A2(n_237),
.B(n_239),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_856),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_SL g1067 ( 
.A1(n_915),
.A2(n_21),
.B(n_22),
.C(n_25),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_821),
.B(n_25),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_865),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_971),
.B(n_250),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_868),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_912),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_867),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_821),
.B(n_33),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_884),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_964),
.A2(n_280),
.B(n_251),
.C(n_282),
.Y(n_1076)
);

O2A1O1Ixp5_ASAP7_75t_L g1077 ( 
.A1(n_934),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_924),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_950),
.A2(n_282),
.B1(n_268),
.B2(n_435),
.Y(n_1079)
);

O2A1O1Ixp5_ASAP7_75t_L g1080 ( 
.A1(n_896),
.A2(n_39),
.B(n_44),
.C(n_49),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_968),
.B(n_51),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_867),
.B(n_825),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_864),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_929),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_957),
.A2(n_268),
.B(n_282),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_846),
.B(n_863),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_872),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_863),
.B(n_461),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_887),
.A2(n_895),
.B(n_894),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_SL g1090 ( 
.A1(n_848),
.A2(n_54),
.B(n_461),
.C(n_452),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_863),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_894),
.A2(n_282),
.B(n_452),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_878),
.B(n_461),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_833),
.B(n_461),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_991),
.B(n_452),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_919),
.A2(n_969),
.B(n_957),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_954),
.B(n_56),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_954),
.B(n_68),
.Y(n_1098)
);

OAI21xp33_ASAP7_75t_L g1099 ( 
.A1(n_973),
.A2(n_71),
.B(n_74),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_914),
.A2(n_76),
.B(n_85),
.C(n_91),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_885),
.B(n_93),
.Y(n_1101)
);

AO32x1_ASAP7_75t_L g1102 ( 
.A1(n_931),
.A2(n_94),
.A3(n_98),
.B1(n_103),
.B2(n_109),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_850),
.B(n_112),
.Y(n_1103)
);

AO32x2_ASAP7_75t_L g1104 ( 
.A1(n_965),
.A2(n_128),
.A3(n_129),
.B1(n_137),
.B2(n_141),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_852),
.B(n_149),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_890),
.B(n_150),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_849),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_904),
.B(n_152),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_908),
.B(n_158),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_893),
.B(n_159),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_954),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_880),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_901),
.Y(n_1113)
);

AND2x2_ASAP7_75t_SL g1114 ( 
.A(n_877),
.B(n_167),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_883),
.A2(n_985),
.B1(n_869),
.B2(n_902),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_SL g1116 ( 
.A1(n_855),
.A2(n_913),
.B(n_947),
.C(n_928),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_901),
.B(n_958),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_956),
.B(n_893),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_882),
.Y(n_1119)
);

INVxp67_ASAP7_75t_SL g1120 ( 
.A(n_882),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_958),
.B(n_943),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_882),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_898),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_943),
.B(n_831),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_906),
.A2(n_855),
.B(n_897),
.Y(n_1125)
);

BUFx4f_ASAP7_75t_L g1126 ( 
.A(n_936),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_991),
.B(n_823),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_920),
.Y(n_1128)
);

INVxp67_ASAP7_75t_L g1129 ( 
.A(n_986),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_923),
.A2(n_963),
.B(n_933),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_944),
.A2(n_888),
.B(n_886),
.C(n_925),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_940),
.B(n_889),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_909),
.A2(n_974),
.B(n_946),
.C(n_910),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_943),
.B(n_831),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_SL g1135 ( 
.A(n_917),
.B(n_918),
.C(n_875),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_953),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_891),
.B(n_976),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_933),
.A2(n_938),
.B(n_963),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_984),
.B(n_987),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_891),
.B(n_966),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_966),
.B(n_936),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_930),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_994),
.B(n_993),
.Y(n_1143)
);

AO21x2_ASAP7_75t_L g1144 ( 
.A1(n_978),
.A2(n_916),
.B(n_977),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_870),
.A2(n_899),
.B(n_981),
.C(n_983),
.Y(n_1145)
);

OAI22x1_ASAP7_75t_L g1146 ( 
.A1(n_877),
.A2(n_942),
.B1(n_992),
.B2(n_994),
.Y(n_1146)
);

NOR3xp33_ASAP7_75t_L g1147 ( 
.A(n_1018),
.B(n_928),
.C(n_913),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1004),
.B(n_966),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1027),
.B(n_966),
.Y(n_1149)
);

AOI211x1_ASAP7_75t_L g1150 ( 
.A1(n_1068),
.A2(n_938),
.B(n_970),
.C(n_873),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1032),
.B(n_975),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1027),
.B(n_952),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1045),
.B(n_951),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1073),
.A2(n_970),
.B1(n_911),
.B2(n_967),
.C(n_876),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1026),
.B(n_936),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_1011),
.B(n_922),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1096),
.A2(n_935),
.B(n_989),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1034),
.A2(n_962),
.B(n_988),
.Y(n_1158)
);

NOR2x1_ASAP7_75t_SL g1159 ( 
.A(n_1021),
.B(n_939),
.Y(n_1159)
);

O2A1O1Ixp5_ASAP7_75t_L g1160 ( 
.A1(n_1076),
.A2(n_1010),
.B(n_1016),
.C(n_1030),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1009),
.B(n_992),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1005),
.B(n_992),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1031),
.A2(n_978),
.B(n_992),
.Y(n_1163)
);

NAND3x1_ASAP7_75t_L g1164 ( 
.A(n_1132),
.B(n_945),
.C(n_932),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1005),
.B(n_972),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_996),
.B(n_983),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_1017),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_999),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1082),
.B(n_945),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_L g1170 ( 
.A(n_1044),
.B(n_945),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_1113),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1048),
.A2(n_939),
.B(n_949),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1126),
.Y(n_1173)
);

NAND2x1p5_ASAP7_75t_L g1174 ( 
.A(n_996),
.B(n_961),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_996),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1118),
.B(n_932),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1083),
.Y(n_1177)
);

BUFx10_ASAP7_75t_L g1178 ( 
.A(n_1060),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1125),
.A2(n_979),
.B(n_932),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1043),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1082),
.B(n_949),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1111),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1001),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1114),
.A2(n_960),
.B1(n_1062),
.B2(n_1022),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_1044),
.B(n_1013),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1092),
.A2(n_1130),
.B(n_1138),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1019),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_SL g1188 ( 
.A(n_996),
.B(n_1038),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1107),
.A2(n_1128),
.B1(n_1056),
.B2(n_1142),
.Y(n_1189)
);

AO21x1_ASAP7_75t_L g1190 ( 
.A1(n_1010),
.A2(n_1115),
.B(n_1046),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1113),
.B(n_1024),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1115),
.A2(n_1015),
.B1(n_1055),
.B2(n_1059),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1013),
.B(n_1038),
.Y(n_1193)
);

AOI21x1_ASAP7_75t_L g1194 ( 
.A1(n_997),
.A2(n_1061),
.B(n_1146),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1062),
.B(n_1070),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1014),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1035),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1074),
.B(n_1053),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1055),
.B(n_1023),
.Y(n_1199)
);

NAND3x1_ASAP7_75t_L g1200 ( 
.A(n_1058),
.B(n_1110),
.C(n_1112),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1099),
.A2(n_1131),
.B(n_1135),
.C(n_1145),
.Y(n_1201)
);

BUFx2_ASAP7_75t_SL g1202 ( 
.A(n_1038),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1063),
.B(n_1066),
.Y(n_1203)
);

OA21x2_ASAP7_75t_L g1204 ( 
.A1(n_1033),
.A2(n_1109),
.B(n_1108),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1056),
.A2(n_1090),
.B(n_1012),
.C(n_1015),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1059),
.A2(n_1081),
.B1(n_1071),
.B2(n_1087),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1060),
.B(n_1049),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1069),
.B(n_1029),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1136),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1075),
.B(n_1139),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1081),
.B(n_1137),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_1143),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1002),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1129),
.B(n_1007),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1111),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1116),
.A2(n_1028),
.B(n_1044),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_L g1217 ( 
.A(n_1054),
.B(n_1046),
.C(n_1077),
.Y(n_1217)
);

AO32x2_ASAP7_75t_L g1218 ( 
.A1(n_1104),
.A2(n_1144),
.A3(n_1067),
.B1(n_1021),
.B2(n_1061),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1101),
.A2(n_1108),
.A3(n_1109),
.B(n_1106),
.Y(n_1219)
);

NOR2x1_ASAP7_75t_SL g1220 ( 
.A(n_1121),
.B(n_1141),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1039),
.B(n_1013),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1003),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1037),
.B(n_1051),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1042),
.A2(n_1079),
.B(n_1133),
.C(n_1080),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1111),
.Y(n_1225)
);

AOI21xp33_ASAP7_75t_L g1226 ( 
.A1(n_1000),
.A2(n_1095),
.B(n_1143),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1093),
.B(n_1047),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1006),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1051),
.B(n_1091),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1101),
.A2(n_1094),
.B(n_1025),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1144),
.A2(n_1102),
.B(n_1041),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1050),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_1050),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1094),
.A2(n_1065),
.B(n_1041),
.Y(n_1234)
);

OAI22x1_ASAP7_75t_L g1235 ( 
.A1(n_1105),
.A2(n_1117),
.B1(n_1057),
.B2(n_1104),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1102),
.A2(n_1140),
.B(n_1134),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1091),
.B(n_1052),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1050),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1025),
.A2(n_1124),
.B(n_1036),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1100),
.A2(n_1097),
.B(n_1098),
.Y(n_1240)
);

NAND2xp33_ASAP7_75t_L g1241 ( 
.A(n_1020),
.B(n_1122),
.Y(n_1241)
);

NAND2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1140),
.B(n_998),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_L g1243 ( 
.A(n_1040),
.B(n_1119),
.C(n_1122),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1119),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1036),
.A2(n_1088),
.B(n_1064),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1105),
.B(n_998),
.Y(n_1246)
);

OR2x6_ASAP7_75t_L g1247 ( 
.A(n_1086),
.B(n_1103),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1072),
.A2(n_1078),
.B(n_1084),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1120),
.A2(n_711),
.B1(n_530),
.B2(n_948),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1104),
.B(n_1102),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1031),
.A2(n_835),
.B(n_1048),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1085),
.A2(n_1096),
.B(n_1034),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_999),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1045),
.B(n_690),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1031),
.A2(n_835),
.B(n_1048),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1031),
.A2(n_835),
.B(n_1048),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1004),
.B(n_840),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1004),
.B(n_840),
.Y(n_1258)
);

NAND2x1_ASAP7_75t_L g1259 ( 
.A(n_1021),
.B(n_945),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1044),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1001),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1085),
.A2(n_1096),
.B(n_1034),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1085),
.A2(n_1096),
.B(n_1034),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_996),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1004),
.A2(n_835),
.B1(n_1005),
.B2(n_837),
.Y(n_1265)
);

INVx5_ASAP7_75t_L g1266 ( 
.A(n_1044),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1085),
.A2(n_1096),
.B(n_1034),
.Y(n_1267)
);

AOI21xp33_ASAP7_75t_L g1268 ( 
.A1(n_1010),
.A2(n_1114),
.B(n_879),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1018),
.A2(n_661),
.B(n_905),
.C(n_879),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1031),
.A2(n_1089),
.A3(n_1125),
.B(n_1138),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1085),
.A2(n_1096),
.B(n_1034),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1085),
.A2(n_1096),
.B(n_1034),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1018),
.A2(n_661),
.B(n_905),
.C(n_879),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_SL g1274 ( 
.A1(n_1082),
.A2(n_1008),
.B(n_1005),
.Y(n_1274)
);

AOI221x1_ASAP7_75t_L g1275 ( 
.A1(n_1099),
.A2(n_1076),
.B1(n_1146),
.B2(n_1046),
.C(n_1010),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1005),
.B(n_835),
.Y(n_1276)
);

BUFx8_ASAP7_75t_L g1277 ( 
.A(n_1017),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1018),
.A2(n_711),
.B(n_879),
.C(n_509),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1125),
.A2(n_997),
.B(n_1030),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1005),
.B(n_835),
.Y(n_1280)
);

NOR2xp67_ASAP7_75t_L g1281 ( 
.A(n_996),
.B(n_717),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1031),
.A2(n_835),
.B(n_1048),
.Y(n_1282)
);

AOI221xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1073),
.A2(n_1010),
.B1(n_790),
.B2(n_879),
.C(n_1018),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1045),
.B(n_690),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1045),
.B(n_690),
.Y(n_1285)
);

INVxp67_ASAP7_75t_SL g1286 ( 
.A(n_1011),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1018),
.A2(n_661),
.B(n_905),
.C(n_879),
.Y(n_1287)
);

BUFx4f_ASAP7_75t_L g1288 ( 
.A(n_1044),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1004),
.B(n_840),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1031),
.A2(n_835),
.B(n_1048),
.Y(n_1290)
);

AO22x2_ASAP7_75t_L g1291 ( 
.A1(n_1115),
.A2(n_1127),
.B1(n_1010),
.B2(n_1046),
.Y(n_1291)
);

AOI21xp33_ASAP7_75t_L g1292 ( 
.A1(n_1010),
.A2(n_1114),
.B(n_879),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1031),
.A2(n_835),
.B(n_1048),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1004),
.B(n_840),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1045),
.B(n_690),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1031),
.A2(n_835),
.B(n_1048),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1004),
.B(n_840),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1031),
.A2(n_835),
.B(n_1048),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1001),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1031),
.A2(n_835),
.B(n_1048),
.Y(n_1300)
);

BUFx8_ASAP7_75t_L g1301 ( 
.A(n_1173),
.Y(n_1301)
);

INVx5_ASAP7_75t_L g1302 ( 
.A(n_1185),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1201),
.A2(n_1192),
.B(n_1268),
.Y(n_1303)
);

OA21x2_ASAP7_75t_L g1304 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1262),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1288),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1291),
.A2(n_1268),
.B1(n_1292),
.B2(n_1190),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1203),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1288),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1222),
.Y(n_1309)
);

INVx5_ASAP7_75t_L g1310 ( 
.A(n_1185),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1267),
.A2(n_1272),
.B(n_1271),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1183),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1279),
.A2(n_1186),
.B(n_1231),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1163),
.A2(n_1279),
.B(n_1230),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1257),
.B(n_1258),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1251),
.A2(n_1256),
.B(n_1255),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1187),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1277),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1277),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1197),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1270),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1167),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1282),
.A2(n_1293),
.B(n_1290),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1261),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1270),
.Y(n_1325)
);

BUFx4_ASAP7_75t_SL g1326 ( 
.A(n_1233),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1296),
.A2(n_1300),
.B(n_1298),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1158),
.A2(n_1172),
.B(n_1157),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1253),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_SL g1330 ( 
.A1(n_1292),
.A2(n_1280),
.B(n_1276),
.C(n_1289),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1265),
.A2(n_1294),
.B1(n_1297),
.B2(n_1276),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1210),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1265),
.A2(n_1280),
.B1(n_1192),
.B2(n_1291),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1195),
.A2(n_1200),
.B1(n_1184),
.B2(n_1249),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1160),
.A2(n_1216),
.B(n_1234),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1250),
.A2(n_1206),
.B1(n_1211),
.B2(n_1287),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1250),
.A2(n_1206),
.B1(n_1269),
.B2(n_1273),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1232),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1234),
.A2(n_1179),
.B(n_1236),
.Y(n_1339)
);

AND2x2_ASAP7_75t_SL g1340 ( 
.A(n_1170),
.B(n_1241),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1167),
.Y(n_1341)
);

NOR2xp67_ASAP7_75t_L g1342 ( 
.A(n_1214),
.B(n_1177),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_1196),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1217),
.A2(n_1199),
.B1(n_1205),
.B2(n_1286),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1182),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1179),
.A2(n_1204),
.B(n_1274),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1239),
.A2(n_1245),
.B(n_1240),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1299),
.Y(n_1348)
);

AOI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1275),
.A2(n_1235),
.B(n_1204),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1240),
.A2(n_1169),
.B(n_1162),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1283),
.A2(n_1278),
.B(n_1224),
.Y(n_1351)
);

NOR2x1_ASAP7_75t_SL g1352 ( 
.A(n_1202),
.B(n_1266),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1169),
.A2(n_1165),
.B(n_1181),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1199),
.B(n_1212),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1209),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1217),
.A2(n_1208),
.B1(n_1189),
.B2(n_1156),
.Y(n_1356)
);

AOI21xp33_ASAP7_75t_L g1357 ( 
.A1(n_1283),
.A2(n_1154),
.B(n_1243),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1198),
.A2(n_1151),
.B1(n_1191),
.B2(n_1152),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1165),
.A2(n_1164),
.B(n_1259),
.Y(n_1359)
);

INVx8_ASAP7_75t_L g1360 ( 
.A(n_1173),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1215),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1225),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_SL g1363 ( 
.A1(n_1220),
.A2(n_1159),
.B(n_1223),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1221),
.B(n_1171),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1148),
.A2(n_1149),
.B(n_1155),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1260),
.A2(n_1243),
.B(n_1242),
.Y(n_1366)
);

AOI22x1_ASAP7_75t_L g1367 ( 
.A1(n_1175),
.A2(n_1264),
.B1(n_1244),
.B2(n_1227),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1270),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1254),
.B(n_1295),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1173),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1213),
.Y(n_1371)
);

OR2x6_ASAP7_75t_L g1372 ( 
.A(n_1246),
.B(n_1242),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1260),
.A2(n_1237),
.B(n_1176),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1188),
.B(n_1175),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_SL g1375 ( 
.A1(n_1226),
.A2(n_1264),
.B(n_1238),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1229),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1244),
.Y(n_1377)
);

OAI22x1_ASAP7_75t_L g1378 ( 
.A1(n_1207),
.A2(n_1180),
.B1(n_1161),
.B2(n_1285),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1228),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1171),
.B(n_1284),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1166),
.A2(n_1174),
.B(n_1248),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1226),
.B(n_1178),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1248),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1150),
.A2(n_1281),
.B1(n_1147),
.B2(n_1153),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1178),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1247),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1247),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1166),
.A2(n_1174),
.B(n_1218),
.Y(n_1388)
);

OAI221xp5_ASAP7_75t_L g1389 ( 
.A1(n_1154),
.A2(n_871),
.B1(n_1268),
.B2(n_1292),
.C(n_1283),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1247),
.B(n_1219),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1219),
.B(n_1218),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1218),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1219),
.B(n_1265),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_SL g1394 ( 
.A1(n_1195),
.A2(n_871),
.B1(n_768),
.B2(n_711),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1262),
.Y(n_1395)
);

BUFx2_ASAP7_75t_R g1396 ( 
.A(n_1257),
.Y(n_1396)
);

AO21x2_ASAP7_75t_L g1397 ( 
.A1(n_1231),
.A2(n_1163),
.B(n_1194),
.Y(n_1397)
);

NOR2xp67_ASAP7_75t_L g1398 ( 
.A(n_1249),
.B(n_1214),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1265),
.B(n_1199),
.Y(n_1399)
);

AOI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1268),
.A2(n_1292),
.B1(n_1192),
.B2(n_1265),
.C(n_590),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1262),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1268),
.A2(n_1292),
.B(n_661),
.C(n_1201),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1203),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1288),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1262),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1203),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1265),
.B(n_1199),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1251),
.A2(n_1256),
.B(n_1255),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1168),
.Y(n_1409)
);

INVx5_ASAP7_75t_L g1410 ( 
.A(n_1185),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1173),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1265),
.B(n_1199),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1203),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1254),
.B(n_1284),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1268),
.B(n_1292),
.C(n_1195),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1265),
.A2(n_1258),
.B1(n_1289),
.B2(n_1257),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1262),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1201),
.A2(n_1192),
.B(n_1268),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1203),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1195),
.A2(n_948),
.B1(n_1114),
.B2(n_711),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1203),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1262),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1203),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1288),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1262),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1257),
.A2(n_1289),
.B1(n_1294),
.B2(n_1258),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1265),
.B(n_1199),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1257),
.B(n_1258),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1188),
.B(n_1266),
.Y(n_1429)
);

INVx2_ASAP7_75t_R g1430 ( 
.A(n_1266),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1262),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1262),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1201),
.A2(n_1192),
.B(n_1268),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1268),
.A2(n_1292),
.B(n_1265),
.C(n_879),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1262),
.Y(n_1435)
);

OAI22x1_ASAP7_75t_L g1436 ( 
.A1(n_1184),
.A2(n_1195),
.B1(n_1123),
.B2(n_559),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1203),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1185),
.B(n_1193),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1262),
.Y(n_1439)
);

AO21x2_ASAP7_75t_L g1440 ( 
.A1(n_1231),
.A2(n_1163),
.B(n_1194),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1203),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1426),
.B(n_1315),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1400),
.A2(n_1402),
.B(n_1434),
.Y(n_1443)
);

OA22x2_ASAP7_75t_L g1444 ( 
.A1(n_1334),
.A2(n_1420),
.B1(n_1436),
.B2(n_1378),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1332),
.B(n_1380),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1323),
.A2(n_1408),
.B(n_1346),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1335),
.A2(n_1346),
.B(n_1314),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1426),
.B(n_1315),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1323),
.A2(n_1408),
.B(n_1303),
.Y(n_1449)
);

BUFx10_ASAP7_75t_L g1450 ( 
.A(n_1319),
.Y(n_1450)
);

AOI221x1_ASAP7_75t_SL g1451 ( 
.A1(n_1416),
.A2(n_1331),
.B1(n_1333),
.B2(n_1336),
.C(n_1415),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1351),
.A2(n_1344),
.B(n_1352),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1344),
.A2(n_1416),
.B(n_1303),
.Y(n_1453)
);

AOI21x1_ASAP7_75t_SL g1454 ( 
.A1(n_1321),
.A2(n_1368),
.B(n_1325),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1418),
.A2(n_1433),
.B(n_1327),
.Y(n_1455)
);

AOI21x1_ASAP7_75t_SL g1456 ( 
.A1(n_1321),
.A2(n_1368),
.B(n_1325),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1332),
.B(n_1364),
.Y(n_1457)
);

O2A1O1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1418),
.A2(n_1433),
.B(n_1389),
.C(n_1330),
.Y(n_1458)
);

A2O1A1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1333),
.A2(n_1389),
.B(n_1306),
.C(n_1398),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1393),
.Y(n_1460)
);

INVx3_ASAP7_75t_SL g1461 ( 
.A(n_1322),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1341),
.B(n_1354),
.Y(n_1462)
);

AOI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1336),
.A2(n_1356),
.B1(n_1331),
.B2(n_1337),
.C(n_1357),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1365),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1306),
.A2(n_1394),
.B1(n_1407),
.B2(n_1412),
.Y(n_1465)
);

AOI21x1_ASAP7_75t_SL g1466 ( 
.A1(n_1393),
.A2(n_1427),
.B(n_1412),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1327),
.A2(n_1399),
.B(n_1427),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1391),
.A2(n_1339),
.B(n_1439),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1428),
.B(n_1362),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1428),
.B(n_1307),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1399),
.A2(n_1407),
.B1(n_1343),
.B2(n_1337),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1396),
.A2(n_1356),
.B1(n_1308),
.B2(n_1424),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1345),
.B(n_1361),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1311),
.A2(n_1395),
.B(n_1417),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1401),
.A2(n_1431),
.B(n_1435),
.Y(n_1475)
);

OR2x6_ASAP7_75t_L g1476 ( 
.A(n_1390),
.B(n_1388),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1392),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1403),
.B(n_1406),
.Y(n_1478)
);

INVxp33_ASAP7_75t_L g1479 ( 
.A(n_1342),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1301),
.Y(n_1480)
);

O2A1O1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1357),
.A2(n_1384),
.B(n_1382),
.C(n_1385),
.Y(n_1481)
);

BUFx4_ASAP7_75t_R g1482 ( 
.A(n_1338),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1317),
.B(n_1320),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1413),
.B(n_1419),
.Y(n_1484)
);

AOI221x1_ASAP7_75t_SL g1485 ( 
.A1(n_1324),
.A2(n_1355),
.B1(n_1348),
.B2(n_1437),
.C(n_1441),
.Y(n_1485)
);

AOI221x1_ASAP7_75t_SL g1486 ( 
.A1(n_1421),
.A2(n_1423),
.B1(n_1384),
.B2(n_1382),
.C(n_1326),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1326),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1371),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1313),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1376),
.B(n_1396),
.Y(n_1490)
);

NOR3xp33_ASAP7_75t_L g1491 ( 
.A(n_1349),
.B(n_1424),
.C(n_1404),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1373),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1379),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1305),
.A2(n_1404),
.B1(n_1308),
.B2(n_1340),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1316),
.A2(n_1405),
.B(n_1304),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1353),
.Y(n_1496)
);

O2A1O1Ixp5_ASAP7_75t_L g1497 ( 
.A1(n_1377),
.A2(n_1386),
.B(n_1387),
.C(n_1411),
.Y(n_1497)
);

O2A1O1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1305),
.A2(n_1375),
.B(n_1363),
.C(n_1318),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1422),
.A2(n_1425),
.B(n_1432),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1358),
.B(n_1438),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1301),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1359),
.A2(n_1340),
.B(n_1358),
.C(n_1366),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1397),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1309),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1329),
.B(n_1409),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1372),
.A2(n_1367),
.B1(n_1411),
.B2(n_1374),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1372),
.A2(n_1374),
.B1(n_1429),
.B2(n_1310),
.Y(n_1507)
);

A2O1A1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1350),
.A2(n_1370),
.B(n_1347),
.C(n_1360),
.Y(n_1508)
);

A2O1A1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1381),
.A2(n_1302),
.B(n_1410),
.C(n_1310),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1328),
.A2(n_1383),
.B(n_1440),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1372),
.B(n_1302),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1302),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1310),
.B(n_1410),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1410),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1430),
.B(n_1397),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1304),
.A2(n_1420),
.B1(n_1400),
.B2(n_1415),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1405),
.B(n_1426),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1369),
.B(n_1414),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1426),
.B(n_1315),
.Y(n_1519)
);

INVx5_ASAP7_75t_L g1520 ( 
.A(n_1372),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1426),
.B(n_1315),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1400),
.A2(n_1201),
.B(n_1265),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1426),
.B(n_1315),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1426),
.B(n_1315),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1338),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1326),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1312),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1321),
.Y(n_1528)
);

O2A1O1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1402),
.A2(n_1268),
.B(n_1292),
.C(n_1303),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1369),
.B(n_1414),
.Y(n_1530)
);

AND2x2_ASAP7_75t_SL g1531 ( 
.A(n_1340),
.B(n_1114),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1369),
.B(n_1414),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1488),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1531),
.A2(n_1465),
.B1(n_1471),
.B2(n_1463),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1493),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1476),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1510),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1460),
.B(n_1467),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1477),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1460),
.B(n_1467),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1496),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1455),
.B(n_1485),
.Y(n_1542)
);

OA21x2_ASAP7_75t_L g1543 ( 
.A1(n_1446),
.A2(n_1449),
.B(n_1495),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1527),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1483),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1517),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1489),
.B(n_1468),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1489),
.B(n_1449),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1476),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1446),
.B(n_1455),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1476),
.B(n_1464),
.Y(n_1551)
);

AO21x1_ASAP7_75t_SL g1552 ( 
.A1(n_1515),
.A2(n_1443),
.B(n_1453),
.Y(n_1552)
);

INVx6_ASAP7_75t_L g1553 ( 
.A(n_1520),
.Y(n_1553)
);

AO21x2_ASAP7_75t_L g1554 ( 
.A1(n_1491),
.A2(n_1503),
.B(n_1516),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1447),
.B(n_1503),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1447),
.B(n_1492),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_SL g1557 ( 
.A1(n_1459),
.A2(n_1458),
.B(n_1529),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1462),
.B(n_1528),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1492),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1473),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1478),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1522),
.A2(n_1502),
.B(n_1481),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1445),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1457),
.B(n_1442),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1497),
.A2(n_1508),
.B(n_1509),
.Y(n_1565)
);

AO21x2_ASAP7_75t_L g1566 ( 
.A1(n_1481),
.A2(n_1458),
.B(n_1511),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1474),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1484),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1504),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1505),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1451),
.B(n_1521),
.Y(n_1571)
);

AOI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1475),
.A2(n_1499),
.B(n_1506),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1475),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1518),
.B(n_1532),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1444),
.A2(n_1448),
.B1(n_1524),
.B2(n_1519),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1497),
.Y(n_1576)
);

INVxp67_ASAP7_75t_R g1577 ( 
.A(n_1507),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1514),
.Y(n_1578)
);

INVxp67_ASAP7_75t_R g1579 ( 
.A(n_1494),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1500),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1513),
.A2(n_1512),
.B(n_1523),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1470),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1486),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_1461),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1539),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1548),
.B(n_1530),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1548),
.B(n_1452),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1541),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1538),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1538),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1581),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1537),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1533),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1548),
.B(n_1540),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1540),
.B(n_1550),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1533),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1535),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1546),
.B(n_1466),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1540),
.B(n_1469),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1547),
.Y(n_1600)
);

NOR2x1_ASAP7_75t_L g1601 ( 
.A(n_1562),
.B(n_1498),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1537),
.Y(n_1602)
);

OAI21xp33_ASAP7_75t_L g1603 ( 
.A1(n_1534),
.A2(n_1444),
.B(n_1472),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1543),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1546),
.B(n_1498),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1558),
.B(n_1564),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1550),
.B(n_1547),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1550),
.B(n_1461),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1582),
.B(n_1479),
.Y(n_1609)
);

AO21x2_ASAP7_75t_L g1610 ( 
.A1(n_1542),
.A2(n_1454),
.B(n_1456),
.Y(n_1610)
);

INVx5_ASAP7_75t_L g1611 ( 
.A(n_1553),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1547),
.B(n_1525),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1555),
.B(n_1487),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1573),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1555),
.B(n_1526),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1593),
.Y(n_1616)
);

AOI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1605),
.A2(n_1567),
.B(n_1572),
.Y(n_1617)
);

NOR2x1_ASAP7_75t_SL g1618 ( 
.A(n_1587),
.B(n_1552),
.Y(n_1618)
);

OAI211xp5_ASAP7_75t_SL g1619 ( 
.A1(n_1598),
.A2(n_1571),
.B(n_1542),
.C(n_1534),
.Y(n_1619)
);

OAI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1591),
.A2(n_1583),
.B1(n_1577),
.B2(n_1571),
.Y(n_1620)
);

AO21x2_ASAP7_75t_L g1621 ( 
.A1(n_1592),
.A2(n_1572),
.B(n_1554),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1606),
.B(n_1558),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1587),
.B(n_1551),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1593),
.Y(n_1624)
);

AOI221x1_ASAP7_75t_L g1625 ( 
.A1(n_1603),
.A2(n_1557),
.B1(n_1576),
.B2(n_1582),
.C(n_1578),
.Y(n_1625)
);

OAI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1603),
.A2(n_1575),
.B1(n_1583),
.B2(n_1576),
.C(n_1564),
.Y(n_1626)
);

NOR2x1_ASAP7_75t_SL g1627 ( 
.A(n_1587),
.B(n_1552),
.Y(n_1627)
);

AOI211xp5_ASAP7_75t_L g1628 ( 
.A1(n_1591),
.A2(n_1579),
.B(n_1577),
.C(n_1564),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1593),
.Y(n_1629)
);

OAI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1591),
.A2(n_1577),
.B1(n_1579),
.B2(n_1565),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1612),
.Y(n_1631)
);

AOI222xp33_ASAP7_75t_L g1632 ( 
.A1(n_1591),
.A2(n_1575),
.B1(n_1580),
.B2(n_1563),
.C1(n_1569),
.C2(n_1570),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1596),
.Y(n_1633)
);

AOI221x1_ASAP7_75t_SL g1634 ( 
.A1(n_1589),
.A2(n_1544),
.B1(n_1545),
.B2(n_1568),
.C(n_1561),
.Y(n_1634)
);

BUFx2_ASAP7_75t_SL g1635 ( 
.A(n_1611),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_L g1636 ( 
.A(n_1601),
.B(n_1581),
.C(n_1559),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1594),
.B(n_1560),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1596),
.Y(n_1638)
);

INVxp67_ASAP7_75t_SL g1639 ( 
.A(n_1605),
.Y(n_1639)
);

A2O1A1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1601),
.A2(n_1552),
.B(n_1536),
.C(n_1549),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1596),
.Y(n_1641)
);

NAND4xp25_ASAP7_75t_L g1642 ( 
.A(n_1598),
.B(n_1567),
.C(n_1556),
.D(n_1559),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1601),
.A2(n_1579),
.B1(n_1599),
.B2(n_1606),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1611),
.B(n_1551),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1613),
.Y(n_1645)
);

AOI222xp33_ASAP7_75t_L g1646 ( 
.A1(n_1600),
.A2(n_1580),
.B1(n_1563),
.B2(n_1569),
.C1(n_1570),
.C2(n_1545),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1588),
.Y(n_1647)
);

AOI211xp5_ASAP7_75t_L g1648 ( 
.A1(n_1600),
.A2(n_1544),
.B(n_1562),
.C(n_1567),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1597),
.Y(n_1649)
);

OAI31xp33_ASAP7_75t_L g1650 ( 
.A1(n_1609),
.A2(n_1551),
.A3(n_1562),
.B(n_1490),
.Y(n_1650)
);

INVx4_ASAP7_75t_SL g1651 ( 
.A(n_1644),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1621),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1639),
.B(n_1606),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1616),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1624),
.Y(n_1655)
);

OA21x2_ASAP7_75t_L g1656 ( 
.A1(n_1625),
.A2(n_1636),
.B(n_1617),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1629),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1633),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1622),
.Y(n_1659)
);

CKINVDCx16_ASAP7_75t_R g1660 ( 
.A(n_1635),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1638),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1617),
.A2(n_1614),
.B(n_1602),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1621),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1641),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1649),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1622),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1637),
.B(n_1594),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1637),
.B(n_1594),
.Y(n_1668)
);

INVx4_ASAP7_75t_SL g1669 ( 
.A(n_1644),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1645),
.B(n_1595),
.Y(n_1670)
);

NOR2x1p5_ASAP7_75t_L g1671 ( 
.A(n_1642),
.B(n_1599),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1634),
.B(n_1589),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1645),
.Y(n_1673)
);

INVx4_ASAP7_75t_SL g1674 ( 
.A(n_1644),
.Y(n_1674)
);

BUFx8_ASAP7_75t_L g1675 ( 
.A(n_1623),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1647),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1646),
.B(n_1590),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1650),
.B(n_1608),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1672),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1672),
.B(n_1599),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1651),
.B(n_1595),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1653),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1656),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1654),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1656),
.B(n_1648),
.C(n_1619),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1651),
.B(n_1607),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1653),
.B(n_1659),
.Y(n_1687)
);

OAI21xp33_ASAP7_75t_L g1688 ( 
.A1(n_1678),
.A2(n_1626),
.B(n_1620),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1654),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1651),
.B(n_1607),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1651),
.B(n_1607),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1677),
.B(n_1590),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1666),
.B(n_1590),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1677),
.B(n_1586),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1669),
.B(n_1618),
.Y(n_1695)
);

OAI211xp5_ASAP7_75t_SL g1696 ( 
.A1(n_1673),
.A2(n_1628),
.B(n_1643),
.C(n_1630),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1656),
.B(n_1586),
.Y(n_1697)
);

NAND5xp2_ASAP7_75t_L g1698 ( 
.A(n_1670),
.B(n_1608),
.C(n_1613),
.D(n_1615),
.E(n_1632),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1656),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1655),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_SL g1701 ( 
.A(n_1675),
.B(n_1584),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1669),
.B(n_1618),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1669),
.B(n_1627),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1671),
.B(n_1586),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1671),
.A2(n_1562),
.B1(n_1566),
.B2(n_1554),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1655),
.B(n_1585),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1662),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1662),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1657),
.B(n_1585),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1652),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1673),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1667),
.B(n_1610),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1669),
.B(n_1627),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1657),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1667),
.B(n_1610),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1668),
.B(n_1610),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1658),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1669),
.B(n_1631),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1658),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1699),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1699),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1684),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1684),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_SL g1724 ( 
.A(n_1685),
.B(n_1625),
.C(n_1640),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1679),
.B(n_1668),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1680),
.B(n_1661),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1699),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1687),
.B(n_1661),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1682),
.B(n_1664),
.Y(n_1729)
);

INVxp67_ASAP7_75t_L g1730 ( 
.A(n_1701),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1685),
.A2(n_1562),
.B1(n_1554),
.B2(n_1566),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1713),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1687),
.B(n_1664),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1705),
.A2(n_1688),
.B1(n_1694),
.B2(n_1697),
.Y(n_1734)
);

NOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1683),
.B(n_1584),
.Y(n_1735)
);

INVxp67_ASAP7_75t_L g1736 ( 
.A(n_1701),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1692),
.B(n_1665),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1689),
.Y(n_1738)
);

INVxp67_ASAP7_75t_SL g1739 ( 
.A(n_1683),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1693),
.B(n_1665),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1711),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1711),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1707),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1689),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1688),
.B(n_1574),
.Y(n_1745)
);

O2A1O1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1698),
.A2(n_1696),
.B(n_1700),
.C(n_1717),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1713),
.B(n_1674),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1705),
.A2(n_1640),
.B(n_1609),
.Y(n_1748)
);

OA21x2_ASAP7_75t_L g1749 ( 
.A1(n_1710),
.A2(n_1663),
.B(n_1652),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1700),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1714),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1707),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1713),
.B(n_1674),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1714),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1693),
.B(n_1676),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1754),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1741),
.B(n_1704),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1742),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1721),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1721),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1738),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1730),
.B(n_1675),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1736),
.B(n_1675),
.Y(n_1763)
);

OAI21x1_ASAP7_75t_L g1764 ( 
.A1(n_1721),
.A2(n_1718),
.B(n_1708),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1738),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1745),
.B(n_1675),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1728),
.B(n_1706),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1747),
.B(n_1713),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1728),
.B(n_1733),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1747),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_1720),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1727),
.B(n_1717),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1727),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1744),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1744),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1753),
.B(n_1695),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1749),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1733),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_SL g1779 ( 
.A1(n_1734),
.A2(n_1604),
.B1(n_1718),
.B2(n_1690),
.Y(n_1779)
);

CKINVDCx16_ASAP7_75t_R g1780 ( 
.A(n_1724),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_1732),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1780),
.B(n_1746),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1768),
.B(n_1753),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1758),
.A2(n_1731),
.B(n_1739),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1780),
.B(n_1752),
.C(n_1743),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1771),
.B(n_1725),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1773),
.A2(n_1748),
.B1(n_1726),
.B2(n_1752),
.C(n_1743),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1768),
.B(n_1753),
.Y(n_1788)
);

O2A1O1Ixp33_ASAP7_75t_L g1789 ( 
.A1(n_1771),
.A2(n_1729),
.B(n_1737),
.C(n_1751),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1777),
.A2(n_1735),
.B1(n_1732),
.B2(n_1737),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1781),
.B(n_1778),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1769),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1781),
.B(n_1755),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_1770),
.Y(n_1794)
);

OAI21xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1779),
.A2(n_1776),
.B(n_1763),
.Y(n_1795)
);

OAI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1777),
.A2(n_1708),
.B1(n_1751),
.B2(n_1750),
.C(n_1712),
.Y(n_1796)
);

CKINVDCx14_ASAP7_75t_R g1797 ( 
.A(n_1762),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1769),
.B(n_1773),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1761),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1760),
.B(n_1755),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1760),
.B(n_1722),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1767),
.B(n_1723),
.Y(n_1802)
);

NOR2x1_ASAP7_75t_L g1803 ( 
.A(n_1782),
.B(n_1759),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1792),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1784),
.A2(n_1759),
.B1(n_1772),
.B2(n_1774),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1794),
.B(n_1798),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1800),
.B(n_1756),
.Y(n_1807)
);

NAND2x1_ASAP7_75t_L g1808 ( 
.A(n_1783),
.B(n_1776),
.Y(n_1808)
);

INVx1_ASAP7_75t_SL g1809 ( 
.A(n_1788),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1791),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1797),
.B(n_1766),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1799),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1793),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1802),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1805),
.A2(n_1785),
.B1(n_1784),
.B2(n_1787),
.Y(n_1815)
);

O2A1O1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1803),
.A2(n_1813),
.B(n_1805),
.C(n_1806),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1809),
.B(n_1814),
.Y(n_1817)
);

OAI221xp5_ASAP7_75t_SL g1818 ( 
.A1(n_1807),
.A2(n_1790),
.B1(n_1795),
.B2(n_1789),
.C(n_1796),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1808),
.A2(n_1786),
.B(n_1801),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1810),
.B(n_1756),
.Y(n_1820)
);

OAI221xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1804),
.A2(n_1757),
.B1(n_1767),
.B2(n_1774),
.C(n_1765),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1811),
.A2(n_1765),
.B(n_1761),
.Y(n_1822)
);

NAND3xp33_ASAP7_75t_L g1823 ( 
.A(n_1804),
.B(n_1775),
.C(n_1750),
.Y(n_1823)
);

NAND3xp33_ASAP7_75t_L g1824 ( 
.A(n_1812),
.B(n_1775),
.C(n_1740),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1817),
.Y(n_1825)
);

OAI21xp33_ASAP7_75t_L g1826 ( 
.A1(n_1815),
.A2(n_1812),
.B(n_1764),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1824),
.Y(n_1827)
);

OAI221xp5_ASAP7_75t_SL g1828 ( 
.A1(n_1816),
.A2(n_1764),
.B1(n_1740),
.B2(n_1702),
.C(n_1695),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1823),
.A2(n_1819),
.B1(n_1820),
.B2(n_1822),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1821),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1825),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1825),
.B(n_1686),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1827),
.B(n_1829),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1828),
.B(n_1818),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1826),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1830),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1825),
.Y(n_1837)
);

INVx1_ASAP7_75t_SL g1838 ( 
.A(n_1833),
.Y(n_1838)
);

NAND4xp25_ASAP7_75t_SL g1839 ( 
.A(n_1832),
.B(n_1703),
.C(n_1702),
.D(n_1681),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1831),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1837),
.Y(n_1841)
);

CKINVDCx16_ASAP7_75t_R g1842 ( 
.A(n_1834),
.Y(n_1842)
);

NOR3xp33_ASAP7_75t_L g1843 ( 
.A(n_1842),
.B(n_1836),
.C(n_1835),
.Y(n_1843)
);

OAI211xp5_ASAP7_75t_SL g1844 ( 
.A1(n_1840),
.A2(n_1836),
.B(n_1715),
.C(n_1716),
.Y(n_1844)
);

INVx1_ASAP7_75t_SL g1845 ( 
.A(n_1838),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1845),
.Y(n_1846)
);

O2A1O1Ixp5_ASAP7_75t_L g1847 ( 
.A1(n_1846),
.A2(n_1840),
.B(n_1841),
.C(n_1843),
.Y(n_1847)
);

OAI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1847),
.A2(n_1844),
.B(n_1839),
.Y(n_1848)
);

AND3x2_ASAP7_75t_L g1849 ( 
.A(n_1847),
.B(n_1480),
.C(n_1703),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1848),
.B(n_1686),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1849),
.A2(n_1749),
.B1(n_1710),
.B2(n_1450),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1851),
.A2(n_1450),
.B1(n_1501),
.B2(n_1482),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1850),
.A2(n_1749),
.B1(n_1719),
.B2(n_1691),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1853),
.B(n_1719),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1854),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1855),
.B(n_1852),
.Y(n_1856)
);

CKINVDCx20_ASAP7_75t_R g1857 ( 
.A(n_1856),
.Y(n_1857)
);

OAI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1709),
.B1(n_1706),
.B2(n_1660),
.Y(n_1858)
);

AOI211xp5_ASAP7_75t_L g1859 ( 
.A1(n_1858),
.A2(n_1690),
.B(n_1691),
.C(n_1681),
.Y(n_1859)
);


endmodule