module fake_aes_4562_n_33 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_13;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_6), .B(n_9), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_3), .B(n_8), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_4), .Y(n_14) );
OAI21x1_ASAP7_75t_L g15 ( .A1(n_2), .A2(n_1), .B(n_5), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
INVx2_ASAP7_75t_SL g18 ( .A(n_14), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
CKINVDCx16_ASAP7_75t_R g20 ( .A(n_18), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_16), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_19), .B(n_17), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_21), .B(n_19), .Y(n_23) );
INVx3_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_0), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_1), .Y(n_26) );
NOR2xp67_ASAP7_75t_L g27 ( .A(n_26), .B(n_7), .Y(n_27) );
NAND2x1p5_ASAP7_75t_L g28 ( .A(n_25), .B(n_12), .Y(n_28) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_27), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
NAND4xp75_ASAP7_75t_L g32 ( .A(n_30), .B(n_12), .C(n_13), .D(n_10), .Y(n_32) );
XNOR2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_32), .Y(n_33) );
endmodule