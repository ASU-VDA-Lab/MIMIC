module fake_jpeg_28582_n_367 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_367);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_367;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_20),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_22),
.B(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_0),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_0),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_94),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_44),
.C(n_36),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_41),
.C(n_28),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_43),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_43),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_30),
.B1(n_46),
.B2(n_42),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_96),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_34),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_47),
.B(n_27),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_99),
.Y(n_138)
);

OR2x4_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_26),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_28),
.B1(n_46),
.B2(n_42),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_106),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_67),
.B(n_18),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_109),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_56),
.A2(n_38),
.B1(n_29),
.B2(n_40),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_31),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_82),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_113),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_81),
.A2(n_38),
.B1(n_55),
.B2(n_60),
.Y(n_114)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_122),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_52),
.B1(n_53),
.B2(n_69),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_124),
.B1(n_76),
.B2(n_73),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_39),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_81),
.B(n_69),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_139),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_87),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_125),
.Y(n_154)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_39),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_131),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_34),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_134),
.B(n_78),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_96),
.B(n_41),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_72),
.B(n_68),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_74),
.C(n_98),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_31),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_68),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_83),
.B(n_40),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_116),
.Y(n_157)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_108),
.B1(n_79),
.B2(n_102),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_155),
.B1(n_120),
.B2(n_113),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_164),
.B1(n_168),
.B2(n_135),
.Y(n_175)
);

BUFx4f_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_102),
.B1(n_90),
.B2(n_79),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_166),
.C(n_134),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_90),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_162),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_95),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_165),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_76),
.B1(n_74),
.B2(n_98),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_54),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_110),
.B1(n_58),
.B2(n_60),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_145),
.B1(n_154),
.B2(n_125),
.Y(n_190)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_123),
.B1(n_154),
.B2(n_149),
.Y(n_197)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_178),
.Y(n_196)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_180),
.Y(n_199)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_153),
.B1(n_150),
.B2(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_182),
.B(n_185),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_186),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_111),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_143),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_162),
.C(n_163),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_202),
.C(n_136),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_198),
.B1(n_141),
.B2(n_165),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_192),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_182),
.B(n_160),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_194),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_201),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_184),
.A2(n_149),
.B1(n_143),
.B2(n_157),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_200),
.A2(n_202),
.B(n_171),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_146),
.B1(n_165),
.B2(n_163),
.Y(n_201)
);

AOI32xp33_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_146),
.A3(n_167),
.B1(n_143),
.B2(n_156),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_117),
.Y(n_223)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_187),
.A2(n_204),
.B(n_201),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_207),
.A2(n_213),
.B(n_214),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_187),
.B(n_185),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_216),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_156),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_221),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_211),
.A2(n_218),
.B1(n_208),
.B2(n_223),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_112),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_212),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_146),
.B(n_173),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_171),
.B(n_174),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_194),
.B(n_196),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_181),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_116),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_194),
.C(n_195),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_126),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_225),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_189),
.A2(n_147),
.B(n_180),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_228),
.B(n_240),
.Y(n_258)
);

A2O1A1O1Ixp25_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_215),
.B(n_205),
.C(n_218),
.D(n_214),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_196),
.B1(n_199),
.B2(n_170),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_238),
.B1(n_247),
.B2(n_217),
.Y(n_254)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_170),
.B1(n_150),
.B2(n_147),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_127),
.C(n_178),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_225),
.C(n_219),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_240),
.A2(n_152),
.B1(n_129),
.B2(n_86),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_127),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_211),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_216),
.Y(n_250)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

INVx11_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_205),
.A2(n_152),
.B1(n_128),
.B2(n_130),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_248),
.B(n_258),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_255),
.Y(n_273)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_257),
.C(n_260),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_213),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_253),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_242),
.B1(n_231),
.B2(n_245),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_213),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_212),
.C(n_128),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_132),
.C(n_140),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_142),
.C(n_121),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_129),
.C(n_65),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_SL g262 ( 
.A(n_227),
.B(n_176),
.C(n_152),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_126),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_176),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_137),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_229),
.A2(n_236),
.B1(n_246),
.B2(n_243),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_242),
.B1(n_245),
.B2(n_232),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_230),
.A2(n_121),
.B(n_78),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_247),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_229),
.B(n_19),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_269),
.A2(n_226),
.B1(n_179),
.B2(n_137),
.Y(n_285)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_179),
.Y(n_292)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_280),
.B(n_283),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_256),
.B(n_232),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_285),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_237),
.B1(n_238),
.B2(n_235),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_253),
.A2(n_226),
.B1(n_244),
.B2(n_103),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_287),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_249),
.B(n_261),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_248),
.B(n_258),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_255),
.B(n_115),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_290),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_115),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_259),
.Y(n_307)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_269),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_0),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_257),
.C(n_260),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_290),
.C(n_279),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_274),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_301),
.B(n_309),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_307),
.Y(n_322)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_270),
.B(n_266),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_306),
.A2(n_291),
.B(n_278),
.Y(n_316)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_276),
.Y(n_308)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_281),
.B(n_20),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_296),
.A2(n_288),
.B1(n_273),
.B2(n_266),
.Y(n_310)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_314),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_273),
.B(n_287),
.Y(n_313)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_313),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_295),
.A2(n_305),
.B1(n_299),
.B2(n_298),
.Y(n_314)
);

AOI221xp5_ASAP7_75t_L g328 ( 
.A1(n_316),
.A2(n_297),
.B1(n_18),
.B2(n_4),
.C(n_5),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_300),
.A2(n_279),
.B1(n_289),
.B2(n_179),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_319),
.Y(n_333)
);

AOI21x1_ASAP7_75t_SL g321 ( 
.A1(n_304),
.A2(n_115),
.B(n_97),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_54),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_65),
.C(n_86),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_323),
.B(n_75),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_304),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_332),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_302),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_327),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_297),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_328),
.A2(n_333),
.B1(n_329),
.B2(n_324),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_1),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_331),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_323),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_3),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_3),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_342),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_338),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_330),
.A2(n_320),
.B1(n_313),
.B2(n_321),
.Y(n_340)
);

AOI21x1_ASAP7_75t_L g341 ( 
.A1(n_328),
.A2(n_316),
.B(n_310),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_322),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_311),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_344),
.B(n_345),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_318),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_3),
.C(n_5),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_348),
.B(n_351),
.Y(n_355)
);

OAI321xp33_ASAP7_75t_L g349 ( 
.A1(n_346),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_349)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_349),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_339),
.A2(n_7),
.B(n_8),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_343),
.A2(n_7),
.B1(n_9),
.B2(n_12),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_352),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_9),
.C(n_12),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_353),
.B(n_12),
.C(n_13),
.Y(n_358)
);

NOR3xp33_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_47),
.C(n_27),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_357),
.B(n_358),
.Y(n_361)
);

MAJx2_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_347),
.C(n_354),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_360),
.B(n_362),
.C(n_355),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_356),
.B(n_350),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_363),
.B(n_361),
.C(n_51),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_27),
.C(n_14),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_17),
.C(n_13),
.Y(n_366)
);

OAI21xp33_ASAP7_75t_L g367 ( 
.A1(n_366),
.A2(n_15),
.B(n_17),
.Y(n_367)
);


endmodule