module real_jpeg_2659_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_39;
wire n_36;
wire n_40;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_48;
wire n_26;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_2),
.A2(n_12),
.B1(n_20),
.B2(n_41),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_4),
.A2(n_12),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_4),
.A2(n_19),
.B1(n_46),
.B2(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_16),
.Y(n_15)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_21),
.B1(n_46),
.B2(n_48),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_12),
.C(n_31),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_6),
.A2(n_12),
.B1(n_20),
.B2(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_34),
.Y(n_8)
);

AOI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_24),
.B(n_33),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_17),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_15),
.Y(n_11)
);

INVx3_ASAP7_75t_SL g20 ( 
.A(n_12),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_12),
.A2(n_20),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_17)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_18),
.B1(n_22),
.B2(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_23),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_28),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_44)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_50),
.Y(n_49)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_32),
.B1(n_46),
.B2(n_48),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_55),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_42),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_52),
.B2(n_54),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx6p67_ASAP7_75t_R g48 ( 
.A(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_52),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);


endmodule