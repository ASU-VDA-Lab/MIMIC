module fake_jpeg_2331_n_539 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_539);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_52),
.Y(n_145)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_53),
.Y(n_136)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g120 ( 
.A(n_57),
.Y(n_120)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_68),
.Y(n_108)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_25),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_78),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_25),
.B(n_47),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_69),
.Y(n_160)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_73),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_74),
.Y(n_165)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_51),
.B(n_17),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_41),
.B(n_16),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_97),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_100),
.Y(n_131)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_43),
.B(n_46),
.Y(n_123)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_99),
.B(n_104),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_38),
.A2(n_0),
.B(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_102),
.B(n_0),
.Y(n_144)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_49),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_38),
.B(n_0),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_67),
.B(n_47),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_117),
.B(n_129),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_50),
.B1(n_34),
.B2(n_46),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_119),
.A2(n_161),
.B1(n_162),
.B2(n_6),
.Y(n_224)
);

NAND2x1_ASAP7_75t_SL g204 ( 
.A(n_123),
.B(n_42),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_77),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_66),
.A2(n_49),
.B1(n_44),
.B2(n_32),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_142),
.B1(n_146),
.B2(n_162),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_78),
.A2(n_85),
.B1(n_87),
.B2(n_94),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_74),
.B1(n_80),
.B2(n_88),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_55),
.A2(n_24),
.B1(n_34),
.B2(n_20),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_144),
.B(n_164),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_60),
.A2(n_24),
.B1(n_44),
.B2(n_32),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_146),
.A2(n_142),
.B1(n_161),
.B2(n_119),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_52),
.B(n_69),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_151),
.B(n_152),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_37),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_86),
.B(n_37),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_158),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_96),
.B(n_33),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_57),
.A2(n_33),
.B1(n_27),
.B2(n_22),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_91),
.A2(n_27),
.B1(n_22),
.B2(n_20),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_72),
.B(n_49),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_167),
.B(n_184),
.Y(n_251)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_168),
.B(n_173),
.Y(n_271)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_171),
.A2(n_201),
.B1(n_206),
.B2(n_213),
.Y(n_249)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_150),
.C(n_110),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_174),
.B(n_136),
.C(n_113),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_135),
.A2(n_57),
.B1(n_64),
.B2(n_100),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_175),
.A2(n_189),
.B1(n_200),
.B2(n_207),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx11_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_177),
.A2(n_182),
.B1(n_134),
.B2(n_165),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_178),
.Y(n_254)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_179),
.Y(n_262)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_93),
.B1(n_79),
.B2(n_75),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_183),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_120),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_185),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_186),
.B(n_188),
.Y(n_258)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_123),
.A2(n_64),
.B1(n_70),
.B2(n_56),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_114),
.B(n_101),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_190),
.B(n_191),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_153),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_192),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_108),
.B(n_1),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_194),
.B(n_198),
.Y(n_241)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_195),
.B(n_209),
.Y(n_274)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_196),
.Y(n_245)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

INVx13_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_127),
.A2(n_43),
.A3(n_42),
.B1(n_73),
.B2(n_5),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_122),
.A2(n_43),
.B1(n_2),
.B2(n_3),
.Y(n_200)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_204),
.B(n_212),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_137),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_159),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_145),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_210),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_159),
.A2(n_42),
.B1(n_3),
.B2(n_5),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_211),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_275)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_112),
.Y(n_212)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_214),
.Y(n_273)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_215),
.Y(n_264)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_132),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_226),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_149),
.B(n_2),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_219),
.Y(n_237)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_218),
.A2(n_220),
.B1(n_222),
.B2(n_224),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_139),
.B(n_6),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_165),
.Y(n_234)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_120),
.Y(n_223)
);

NAND2xp33_ASAP7_75t_SL g242 ( 
.A(n_223),
.B(n_160),
.Y(n_242)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_166),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_160),
.B1(n_113),
.B2(n_121),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_107),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_147),
.B(n_6),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_227),
.B(n_136),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_177),
.A2(n_106),
.B1(n_125),
.B2(n_132),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_231),
.A2(n_249),
.B1(n_255),
.B2(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_240),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_242),
.B(n_226),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_201),
.A2(n_121),
.B1(n_107),
.B2(n_125),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_243),
.A2(n_244),
.B1(n_266),
.B2(n_260),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_179),
.B1(n_224),
.B2(n_172),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_196),
.C(n_214),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_169),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_174),
.B(n_155),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_269),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_189),
.A2(n_155),
.B1(n_137),
.B2(n_106),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_204),
.A2(n_15),
.B1(n_8),
.B2(n_9),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_260),
.A2(n_267),
.B1(n_270),
.B2(n_276),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_224),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_175),
.A2(n_193),
.B1(n_205),
.B2(n_182),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_208),
.B(n_15),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_198),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_270)
);

OA22x2_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_207),
.B1(n_200),
.B2(n_203),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_194),
.B(n_11),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_250),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_277),
.B(n_312),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_271),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_278),
.B(n_287),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_280),
.B(n_295),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_281),
.B(n_236),
.C(n_238),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_282),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_284),
.B(n_319),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_224),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_299),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_225),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_286),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_271),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_249),
.A2(n_215),
.B1(n_183),
.B2(n_221),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_288),
.A2(n_290),
.B1(n_297),
.B2(n_298),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_222),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_289),
.B(n_296),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_241),
.A2(n_199),
.B1(n_178),
.B2(n_185),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_220),
.C(n_210),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_228),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_259),
.A2(n_202),
.B1(n_218),
.B2(n_181),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_294),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_176),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_176),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_241),
.A2(n_197),
.B1(n_14),
.B2(n_15),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_241),
.A2(n_267),
.B1(n_235),
.B2(n_270),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_237),
.B(n_15),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_237),
.B(n_268),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_308),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_242),
.A2(n_251),
.B(n_248),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_301),
.A2(n_263),
.B(n_300),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_302),
.B(n_297),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_255),
.A2(n_234),
.B1(n_233),
.B2(n_229),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_256),
.Y(n_304)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_304),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_229),
.A2(n_264),
.B1(n_253),
.B2(n_246),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_229),
.A2(n_264),
.B1(n_253),
.B2(n_246),
.Y(n_306)
);

AND2x4_ASAP7_75t_SL g307 ( 
.A(n_256),
.B(n_257),
.Y(n_307)
);

BUFx8_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_257),
.B(n_274),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_232),
.Y(n_311)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_261),
.B(n_239),
.Y(n_312)
);

BUFx8_ASAP7_75t_L g313 ( 
.A(n_238),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_313),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_232),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_315),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_261),
.B(n_239),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_316),
.Y(n_353)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_232),
.Y(n_317)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_317),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_230),
.A2(n_262),
.B1(n_272),
.B2(n_273),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_318),
.A2(n_320),
.B1(n_247),
.B2(n_245),
.Y(n_324)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_262),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_262),
.A2(n_230),
.B1(n_245),
.B2(n_273),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_285),
.A2(n_310),
.B(n_282),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_321),
.A2(n_320),
.B(n_314),
.Y(n_374)
);

O2A1O1Ixp33_ASAP7_75t_L g322 ( 
.A1(n_298),
.A2(n_306),
.B(n_305),
.C(n_310),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_322),
.B(n_328),
.Y(n_363)
);

INVxp33_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

AO22x1_ASAP7_75t_SL g328 ( 
.A1(n_288),
.A2(n_247),
.B1(n_254),
.B2(n_238),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_291),
.C(n_301),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_292),
.A2(n_254),
.B1(n_263),
.B2(n_236),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_332),
.A2(n_350),
.B1(n_359),
.B2(n_290),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_335),
.B(n_295),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_293),
.B(n_254),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_336),
.B(n_342),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_293),
.B(n_284),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_343),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_283),
.B(n_228),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_263),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_344),
.B(n_346),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_307),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_352),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_292),
.A2(n_302),
.B1(n_303),
.B2(n_278),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_307),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_287),
.B(n_299),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_354),
.B(n_341),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_281),
.B(n_308),
.Y(n_356)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_356),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_307),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_352),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_362),
.C(n_389),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_361),
.A2(n_375),
.B1(n_376),
.B2(n_379),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_291),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_347),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_366),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_353),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_326),
.A2(n_295),
.B1(n_282),
.B2(n_280),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_368),
.A2(n_351),
.B1(n_346),
.B2(n_322),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_304),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_370),
.B(n_372),
.Y(n_409)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_323),
.Y(n_371)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_341),
.B(n_311),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_323),
.Y(n_373)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_373),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_374),
.A2(n_383),
.B(n_386),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_326),
.A2(n_280),
.B1(n_319),
.B2(n_317),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_350),
.A2(n_280),
.B1(n_309),
.B2(n_316),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_380),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_331),
.A2(n_313),
.B1(n_359),
.B2(n_338),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_354),
.B(n_313),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_331),
.A2(n_313),
.B1(n_338),
.B2(n_332),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_381),
.A2(n_390),
.B1(n_392),
.B2(n_355),
.Y(n_413)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_382),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_336),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_384),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_334),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_385),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_342),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_358),
.Y(n_387)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_387),
.Y(n_416)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_388),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_335),
.B(n_344),
.C(n_337),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_333),
.B(n_345),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_338),
.A2(n_322),
.B1(n_321),
.B2(n_329),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_357),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_393),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_383),
.A2(n_349),
.B(n_346),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_394),
.A2(n_403),
.B(n_420),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_396),
.A2(n_422),
.B1(n_386),
.B2(n_384),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_376),
.A2(n_325),
.B1(n_327),
.B2(n_329),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_400),
.B(n_405),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_330),
.C(n_333),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_406),
.C(n_408),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_387),
.A2(n_351),
.B(n_325),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_379),
.A2(n_345),
.B1(n_328),
.B2(n_357),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_362),
.B(n_340),
.C(n_339),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_340),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_339),
.C(n_353),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_417),
.C(n_423),
.Y(n_431)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_413),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_414),
.B(n_415),
.Y(n_447)
);

MAJx2_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_324),
.C(n_355),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_367),
.B(n_328),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_383),
.A2(n_328),
.B(n_364),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_363),
.A2(n_375),
.B1(n_368),
.B2(n_361),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_389),
.B(n_364),
.C(n_382),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_363),
.A2(n_392),
.B1(n_381),
.B2(n_388),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_424),
.B(n_365),
.Y(n_450)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_419),
.Y(n_425)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_425),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_395),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_426),
.B(n_433),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_424),
.Y(n_471)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_395),
.Y(n_430)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_404),
.Y(n_432)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_432),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_421),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_434),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_397),
.B(n_385),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_435),
.B(n_436),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_397),
.B(n_366),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_420),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_439),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_409),
.B(n_377),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_438),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_422),
.A2(n_411),
.B1(n_396),
.B2(n_402),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_378),
.C(n_374),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_440),
.B(n_442),
.C(n_444),
.Y(n_452)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_404),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_441),
.B(n_448),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_378),
.C(n_393),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_401),
.B(n_371),
.C(n_373),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_380),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_445),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_406),
.B(n_391),
.C(n_365),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_410),
.C(n_415),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_418),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_400),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_414),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_451),
.B(n_459),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_428),
.A2(n_449),
.B1(n_450),
.B2(n_437),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_457),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_417),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_408),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_464),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_462),
.B(n_469),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_431),
.B(n_398),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_431),
.B(n_398),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_447),
.Y(n_485)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_468),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_428),
.A2(n_418),
.B1(n_416),
.B2(n_412),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_471),
.A2(n_449),
.B(n_429),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_426),
.B(n_407),
.Y(n_472)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_472),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_454),
.Y(n_473)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_473),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_479),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_442),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_477),
.B(n_483),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_453),
.A2(n_444),
.B(n_443),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_446),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_471),
.A2(n_433),
.B1(n_434),
.B2(n_443),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_484),
.A2(n_469),
.B1(n_457),
.B2(n_463),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_485),
.B(n_453),
.C(n_459),
.Y(n_493)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_458),
.Y(n_486)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_486),
.Y(n_503)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_466),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_487),
.B(n_488),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_439),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_458),
.Y(n_489)
);

NOR3xp33_ASAP7_75t_L g495 ( 
.A(n_489),
.B(n_461),
.C(n_472),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_490),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_467),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_494),
.A2(n_495),
.B(n_500),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_484),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_482),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_452),
.C(n_451),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_497),
.B(n_452),
.C(n_481),
.Y(n_506)
);

XNOR2x1_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_488),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_475),
.B(n_467),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_478),
.A2(n_456),
.B1(n_463),
.B2(n_425),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_501),
.A2(n_502),
.B1(n_504),
.B2(n_430),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_476),
.A2(n_468),
.B1(n_455),
.B2(n_471),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_474),
.A2(n_416),
.B(n_462),
.Y(n_504)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_505),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_508),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_507),
.A2(n_515),
.B1(n_491),
.B2(n_494),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_466),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_483),
.C(n_481),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_511),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_480),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_512),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_491),
.B(n_490),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_480),
.C(n_485),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_513),
.B(n_498),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_516),
.B(n_518),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_514),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_511),
.A2(n_503),
.B1(n_499),
.B2(n_500),
.Y(n_521)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_521),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_523),
.B(n_505),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_522),
.A2(n_509),
.B(n_512),
.Y(n_524)
);

AOI21xp33_ASAP7_75t_L g530 ( 
.A1(n_524),
.A2(n_527),
.B(n_516),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_517),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_520),
.A2(n_510),
.B(n_470),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_530),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_526),
.B(n_517),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_519),
.C(n_528),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_523),
.B(n_448),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_532),
.B1(n_432),
.B2(n_441),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_535),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_407),
.B(n_405),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_403),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_538),
.A2(n_394),
.B(n_447),
.Y(n_539)
);


endmodule