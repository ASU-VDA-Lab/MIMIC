module fake_aes_8704_n_17 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_17);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_17;
wire n_11;
wire n_16;
wire n_13;
wire n_12;
wire n_9;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
AND2x6_ASAP7_75t_L g7 ( .A(n_5), .B(n_1), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_3), .Y(n_8) );
BUFx6f_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
AO21x2_ASAP7_75t_L g11 ( .A1(n_8), .A2(n_0), .B(n_1), .Y(n_11) );
OR2x2_ASAP7_75t_L g12 ( .A(n_10), .B(n_0), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
OR2x2_ASAP7_75t_L g14 ( .A(n_12), .B(n_11), .Y(n_14) );
AOI221xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_13), .B1(n_11), .B2(n_9), .C(n_7), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
AOI222xp33_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_2), .B1(n_4), .B2(n_7), .C1(n_9), .C2(n_15), .Y(n_17) );
endmodule