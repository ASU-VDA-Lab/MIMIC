module fake_jpeg_9418_n_276 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_11),
.B(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_39),
.Y(n_50)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_0),
.C(n_1),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_31),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_65),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_48),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

OR2x2_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_27),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_58),
.B(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_53),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_63),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_20),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_19),
.B1(n_33),
.B2(n_17),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_37),
.B1(n_34),
.B2(n_38),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_77),
.B1(n_86),
.B2(n_60),
.Y(n_102)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_37),
.B1(n_34),
.B2(n_33),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_61),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_37),
.B1(n_34),
.B2(n_19),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_42),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_50),
.C(n_20),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_90),
.B(n_97),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_51),
.B(n_56),
.C(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_92),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_64),
.B(n_50),
.C(n_33),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_98),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_85),
.B(n_89),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_107),
.B1(n_84),
.B2(n_74),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_109),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_60),
.B1(n_54),
.B2(n_17),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_81),
.B(n_83),
.C(n_72),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_103),
.B1(n_68),
.B2(n_81),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_20),
.A3(n_29),
.B1(n_26),
.B2(n_25),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_19),
.B1(n_54),
.B2(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_72),
.B(n_54),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_74),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_23),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_23),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_123),
.B1(n_107),
.B2(n_23),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_80),
.C(n_82),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_98),
.C(n_93),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_137),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_129),
.B1(n_103),
.B2(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_68),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_132),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_80),
.B(n_49),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_80),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_75),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_130),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_91),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_90),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_159),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_95),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_149),
.C(n_151),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_22),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_102),
.B1(n_99),
.B2(n_97),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_95),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_29),
.A3(n_21),
.B1(n_26),
.B2(n_25),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_114),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_155),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_114),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_157),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_104),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_92),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_163),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_92),
.C(n_84),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_16),
.C(n_22),
.Y(n_182)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_164),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_28),
.Y(n_165)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_122),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_107),
.B1(n_30),
.B2(n_28),
.Y(n_167)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_153),
.A2(n_119),
.B1(n_135),
.B2(n_127),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_176),
.B1(n_154),
.B2(n_163),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_174),
.A2(n_186),
.B1(n_189),
.B2(n_191),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_129),
.B1(n_122),
.B2(n_117),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_126),
.B(n_117),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_180),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_24),
.B(n_30),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_185),
.C(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_48),
.C(n_45),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_3),
.B(n_4),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_152),
.C(n_142),
.Y(n_194)
);

AO22x1_ASAP7_75t_SL g189 ( 
.A1(n_159),
.A2(n_46),
.B1(n_48),
.B2(n_45),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_145),
.B(n_29),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_148),
.A2(n_16),
.B1(n_46),
.B2(n_26),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_199),
.C(n_189),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_196),
.B(n_193),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_155),
.Y(n_197)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_181),
.B1(n_173),
.B2(n_180),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_206),
.B1(n_171),
.B2(n_170),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_151),
.C(n_144),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_190),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_203),
.C(n_210),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_205),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_164),
.B1(n_146),
.B2(n_156),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_156),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_208),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_141),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_212),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_141),
.C(n_144),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_159),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_169),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_3),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_172),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_216),
.C(n_222),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_6),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_182),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_224),
.Y(n_232)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_191),
.B(n_169),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_49),
.B(n_26),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_186),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_199),
.B(n_169),
.Y(n_224)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_3),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_192),
.B1(n_210),
.B2(n_200),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_229),
.A2(n_200),
.B1(n_203),
.B2(n_201),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_214),
.A2(n_46),
.B1(n_49),
.B2(n_25),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_25),
.B1(n_21),
.B2(n_5),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_238),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_4),
.C(n_5),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_225),
.C(n_220),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_4),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_6),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_6),
.B(n_7),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_7),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_251),
.C(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_252),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_237),
.B(n_223),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_250),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_227),
.C(n_213),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_216),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_257),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_231),
.C(n_240),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_258),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_246),
.A2(n_224),
.B1(n_239),
.B2(n_232),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_232),
.C(n_222),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_235),
.B(n_217),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_244),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_260),
.A2(n_243),
.B(n_8),
.C(n_9),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_265),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_7),
.CI(n_9),
.CON(n_265),
.SN(n_265)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_266),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.C(n_263),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_254),
.C(n_11),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_272),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_10),
.C(n_12),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_268),
.B(n_12),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_14),
.Y(n_276)
);


endmodule