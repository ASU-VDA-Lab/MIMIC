module fake_jpeg_27071_n_23 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_23);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_23;

wire n_13;
wire n_21;
wire n_10;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_9),
.B(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_15),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_12),
.A2(n_4),
.B1(n_7),
.B2(n_5),
.Y(n_15)
);

AND2x6_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_8),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_16),
.B(n_10),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_18),
.B(n_11),
.Y(n_19)
);

AOI31xp67_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_20),
.A3(n_12),
.B(n_1),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_21),
.A2(n_0),
.B(n_2),
.Y(n_22)
);

AOI21x1_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_0),
.B(n_3),
.Y(n_23)
);


endmodule