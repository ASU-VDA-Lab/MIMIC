module fake_jpeg_20138_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_3),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_1),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_34),
.B(n_30),
.C(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_19),
.B1(n_21),
.B2(n_17),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_49),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_25),
.B1(n_18),
.B2(n_21),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_50),
.B1(n_22),
.B2(n_31),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_27),
.B1(n_16),
.B2(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_29),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_26),
.B(n_25),
.C(n_14),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_22),
.B1(n_20),
.B2(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_56),
.B(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_14),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_9),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_41),
.B1(n_38),
.B2(n_49),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_8),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx10_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_24),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_55),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_75),
.B1(n_52),
.B2(n_66),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_5),
.B1(n_6),
.B2(n_28),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_28),
.B(n_6),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_28),
.Y(n_91)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_52),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_90),
.C(n_94),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_57),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_81),
.B(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_93),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_56),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_97),
.A2(n_72),
.B1(n_85),
.B2(n_83),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_82),
.B1(n_94),
.B2(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_98),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_80),
.B(n_75),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_11),
.B(n_8),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_104),
.B(n_74),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_80),
.C(n_84),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_74),
.C(n_68),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_83),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_110),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_59),
.B(n_9),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_112),
.B(n_10),
.Y(n_115)
);

OAI31xp33_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_99),
.A3(n_11),
.B(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_101),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_118),
.B(n_113),
.C(n_111),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_107),
.C(n_102),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_121),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_118),
.B1(n_111),
.B2(n_116),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_125),
.B(n_98),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_119),
.C(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_127),
.Y(n_129)
);


endmodule