module fake_jpeg_31770_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_39),
.Y(n_79)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_14),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_55),
.Y(n_76)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_46),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_52),
.Y(n_84)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_17),
.B(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_13),
.Y(n_87)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_60),
.B1(n_61),
.B2(n_32),
.Y(n_82)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_24),
.B1(n_30),
.B2(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_62),
.A2(n_64),
.B1(n_67),
.B2(n_69),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_87),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_24),
.B1(n_20),
.B2(n_30),
.Y(n_69)
);

AO22x1_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_28),
.B1(n_30),
.B2(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_71),
.B(n_89),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_78),
.B1(n_91),
.B2(n_52),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_53),
.B(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_86),
.Y(n_100)
);

CKINVDCx9p33_ASAP7_75t_R g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_40),
.A2(n_24),
.B1(n_32),
.B2(n_25),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_83),
.A2(n_94),
.B1(n_28),
.B2(n_45),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_36),
.B(n_26),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_26),
.B(n_28),
.C(n_12),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_42),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_47),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_49),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_28),
.B1(n_12),
.B2(n_3),
.Y(n_94)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_35),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_98),
.B(n_125),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_92),
.B(n_48),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_68),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_111),
.B1(n_134),
.B2(n_72),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_104),
.B(n_109),
.Y(n_161)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_76),
.B(n_89),
.C(n_80),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_84),
.B(n_88),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_49),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_56),
.B1(n_47),
.B2(n_37),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_57),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_51),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_118),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_117),
.A2(n_119),
.B1(n_66),
.B2(n_90),
.Y(n_168)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_45),
.B1(n_44),
.B2(n_27),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_123),
.Y(n_159)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_74),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_74),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_126),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_87),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_1),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_131),
.B1(n_132),
.B2(n_72),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_68),
.Y(n_129)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_74),
.Y(n_130)
);

INVx2_ASAP7_75t_R g142 ( 
.A(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_1),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_1),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_65),
.A2(n_27),
.B1(n_45),
.B2(n_12),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_84),
.B(n_63),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_135),
.A2(n_143),
.B(n_164),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_138),
.B(n_139),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_103),
.B1(n_124),
.B2(n_107),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_148),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_63),
.B(n_88),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_144),
.A2(n_167),
.B1(n_129),
.B2(n_102),
.Y(n_192)
);

BUFx4f_ASAP7_75t_SL g145 ( 
.A(n_114),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_145),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_115),
.A2(n_68),
.B1(n_90),
.B2(n_85),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_111),
.B1(n_99),
.B2(n_134),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_125),
.Y(n_170)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_122),
.A2(n_95),
.B(n_2),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_166),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_90),
.B1(n_85),
.B2(n_95),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_129),
.B(n_106),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_171),
.B(n_202),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_175),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_174),
.A2(n_196),
.B1(n_197),
.B2(n_144),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_98),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_100),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_184),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_142),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_100),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_99),
.C(n_109),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_205),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_116),
.B1(n_99),
.B2(n_104),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_192),
.B1(n_153),
.B2(n_136),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_131),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_191),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_146),
.B(n_127),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_188),
.B(n_204),
.Y(n_220)
);

AO21x2_ASAP7_75t_L g190 ( 
.A1(n_142),
.A2(n_106),
.B(n_130),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_194),
.B(n_145),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_108),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_105),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_139),
.A2(n_108),
.B1(n_113),
.B2(n_123),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_143),
.A2(n_110),
.B1(n_118),
.B2(n_126),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_132),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_133),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_148),
.B(n_112),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_101),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_101),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_189),
.A2(n_135),
.B(n_138),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_206),
.A2(n_217),
.B(n_223),
.Y(n_244)
);

NAND2xp33_ASAP7_75t_SL g207 ( 
.A(n_193),
.B(n_135),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_218),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_219),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_189),
.A2(n_167),
.B1(n_161),
.B2(n_156),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_145),
.B1(n_159),
.B2(n_158),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_214),
.A2(n_230),
.B(n_190),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_172),
.A2(n_145),
.B(n_166),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_172),
.A2(n_153),
.B1(n_158),
.B2(n_165),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_171),
.B1(n_186),
.B2(n_187),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_233),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_171),
.A2(n_147),
.B(n_150),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_228),
.B(n_204),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_172),
.A2(n_136),
.B1(n_66),
.B2(n_150),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_175),
.B(n_136),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_191),
.B(n_199),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_147),
.B(n_66),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_200),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_236),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_173),
.A2(n_202),
.B(n_190),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_140),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_231),
.B(n_190),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_147),
.B1(n_152),
.B2(n_140),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_170),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_197),
.B1(n_185),
.B2(n_181),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_176),
.Y(n_263)
);

BUFx12_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_255),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_240),
.A2(n_247),
.B(n_265),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_178),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_263),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_177),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_177),
.Y(n_246)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_178),
.C(n_194),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_250),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_236),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_252),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_182),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_188),
.C(n_190),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_260),
.C(n_264),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_237),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_190),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_256),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_208),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_259),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_198),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_195),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_183),
.C(n_180),
.Y(n_260)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_217),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_262),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_176),
.C(n_179),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_230),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_266),
.A2(n_221),
.B1(n_211),
.B2(n_235),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_209),
.B1(n_213),
.B2(n_244),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_277),
.B1(n_279),
.B2(n_240),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_206),
.C(n_219),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_244),
.A2(n_214),
.B1(n_210),
.B2(n_207),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_223),
.B1(n_222),
.B2(n_228),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_245),
.A2(n_201),
.B(n_215),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_283),
.B(n_243),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_234),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_245),
.A2(n_201),
.B(n_212),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_245),
.B1(n_251),
.B2(n_249),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_274),
.B1(n_201),
.B2(n_239),
.Y(n_307)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_290),
.Y(n_306)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_242),
.B(n_246),
.C(n_258),
.D(n_256),
.Y(n_291)
);

BUFx12_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_276),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_249),
.B(n_256),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_272),
.B(n_284),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_257),
.C(n_254),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_298),
.C(n_268),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_296),
.Y(n_301)
);

AOI221xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_261),
.B1(n_232),
.B2(n_212),
.C(n_208),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_279),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_268),
.C(n_282),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_304),
.Y(n_309)
);

O2A1O1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_285),
.B(n_271),
.C(n_277),
.Y(n_303)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_286),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_307),
.A2(n_162),
.B1(n_160),
.B2(n_149),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_312),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_298),
.B(n_140),
.Y(n_312)
);

AND2x6_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_162),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_306),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_308),
.B1(n_316),
.B2(n_315),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_SL g315 ( 
.A1(n_305),
.A2(n_152),
.B(n_160),
.C(n_149),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_152),
.B1(n_27),
.B2(n_6),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_322),
.B(n_311),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_320),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_321),
.A2(n_2),
.B(n_6),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_318),
.C(n_319),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_322),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_328),
.B1(n_329),
.B2(n_324),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_7),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_330),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_9),
.B(n_10),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);


endmodule