module fake_jpeg_17234_n_185 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NAND2x1_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_2),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_28),
.Y(n_61)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_44),
.Y(n_56)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_53),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_25),
.B1(n_19),
.B2(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_60),
.B1(n_66),
.B2(n_4),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_32),
.A2(n_25),
.B1(n_24),
.B2(n_31),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_15),
.B1(n_29),
.B2(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_32),
.B(n_16),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_15),
.B1(n_30),
.B2(n_22),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_22),
.B1(n_23),
.B2(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_24),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_75),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_36),
.C(n_26),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_56),
.C(n_66),
.Y(n_100)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_77),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_46),
.B1(n_51),
.B2(n_58),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_86),
.B1(n_67),
.B2(n_48),
.Y(n_106)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_37),
.A3(n_27),
.B1(n_26),
.B2(n_18),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_91),
.B(n_8),
.Y(n_113)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_14),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_26),
.B1(n_5),
.B2(n_6),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_14),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_93),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_37),
.B1(n_5),
.B2(n_6),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_81),
.B1(n_49),
.B2(n_68),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_66),
.B1(n_50),
.B2(n_63),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_57),
.A2(n_4),
.B(n_7),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_115),
.B1(n_84),
.B2(n_74),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_55),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_101),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_70),
.C(n_86),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_56),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_110),
.Y(n_120)
);

XOR2x1_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_108),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_84),
.C(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_69),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_8),
.B(n_9),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_66),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_113),
.A2(n_91),
.B(n_94),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_89),
.B1(n_92),
.B2(n_71),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_50),
.B1(n_63),
.B2(n_12),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_126),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_131),
.B(n_132),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_122),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_82),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_105),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_106),
.C(n_110),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_93),
.B(n_77),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_93),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_127),
.C(n_98),
.Y(n_138)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_101),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_139),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_SL g155 ( 
.A1(n_138),
.A2(n_144),
.A3(n_119),
.B1(n_131),
.B2(n_111),
.C1(n_130),
.C2(n_10),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_114),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_146),
.B(n_132),
.Y(n_153)
);

AOI322xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_102),
.A3(n_113),
.B1(n_115),
.B2(n_111),
.C1(n_12),
.C2(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_145),
.B(n_121),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_111),
.Y(n_146)
);

BUFx12f_ASAP7_75t_SL g149 ( 
.A(n_136),
.Y(n_149)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_153),
.B(n_155),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_128),
.B1(n_126),
.B2(n_125),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_146),
.B1(n_140),
.B2(n_135),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_157),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_82),
.B1(n_124),
.B2(n_87),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_142),
.B(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_147),
.B(n_117),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_117),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_95),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_147),
.A3(n_146),
.B1(n_139),
.B2(n_135),
.C1(n_140),
.C2(n_142),
.Y(n_159)
);

AOI31xp67_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_165),
.A3(n_157),
.B(n_150),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_160),
.A2(n_148),
.B1(n_150),
.B2(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_141),
.A3(n_73),
.B1(n_85),
.B2(n_95),
.C1(n_103),
.C2(n_80),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_162),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_73),
.B1(n_85),
.B2(n_87),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_168),
.B(n_172),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_164),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_171),
.A2(n_160),
.B1(n_164),
.B2(n_11),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_163),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_11),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_166),
.C(n_167),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_176),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_11),
.A3(n_170),
.B1(n_171),
.B2(n_174),
.C1(n_175),
.C2(n_176),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_177),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_179),
.B(n_180),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_178),
.B(n_180),
.Y(n_182)
);

BUFx24_ASAP7_75t_SL g184 ( 
.A(n_182),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_183),
.Y(n_185)
);


endmodule