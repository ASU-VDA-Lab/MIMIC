module fake_jpeg_29866_n_265 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_60),
.Y(n_72)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_24),
.B(n_39),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_24),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_17),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_18),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_21),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_2),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_64),
.Y(n_73)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_66),
.Y(n_79)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_70),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_74),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_77),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_30),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_31),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_99),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_36),
.C(n_34),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_9),
.C(n_14),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_88),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_36),
.B1(n_34),
.B2(n_26),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_83),
.A2(n_6),
.B1(n_9),
.B2(n_12),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_27),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_27),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_92),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_41),
.B(n_11),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_62),
.B(n_12),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_25),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_20),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_6),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_51),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_120),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_79),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_114),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_53),
.B1(n_67),
.B2(n_49),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_104),
.B1(n_91),
.B2(n_102),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_72),
.Y(n_114)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_84),
.B1(n_71),
.B2(n_90),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_3),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

AO21x2_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_4),
.B(n_5),
.Y(n_124)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_127),
.B1(n_90),
.B2(n_87),
.Y(n_158)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_83),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_135),
.Y(n_155)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_84),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_69),
.B1(n_17),
.B2(n_15),
.Y(n_141)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_87),
.Y(n_157)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_141),
.A2(n_135),
.B1(n_128),
.B2(n_112),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_113),
.B1(n_130),
.B2(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_68),
.B(n_81),
.C(n_74),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_160),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_158),
.B1(n_128),
.B2(n_111),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_101),
.B1(n_90),
.B2(n_71),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_98),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_98),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_120),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_102),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_115),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_165),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_106),
.B(n_138),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_161),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_124),
.B(n_127),
.C(n_133),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_151),
.B(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_138),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_175),
.B(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_178),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_107),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_107),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_184),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_141),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_160),
.B(n_139),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_150),
.C(n_162),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_152),
.B1(n_159),
.B2(n_166),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_158),
.A2(n_124),
.B1(n_118),
.B2(n_125),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_143),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_144),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_190),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_147),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_191),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_193),
.A2(n_174),
.B1(n_178),
.B2(n_188),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_186),
.B1(n_183),
.B2(n_161),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_124),
.C(n_139),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_204),
.A2(n_176),
.B(n_180),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_108),
.B(n_148),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_189),
.B(n_170),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_166),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_207),
.B(n_177),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_167),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_213),
.B(n_216),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_169),
.B1(n_168),
.B2(n_187),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_215),
.C(n_224),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_182),
.C(n_185),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_182),
.B(n_169),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_197),
.B(n_172),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_223),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_183),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_221),
.A2(n_206),
.B1(n_196),
.B2(n_195),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_200),
.B(n_146),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_146),
.Y(n_224)
);

OAI321xp33_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_199),
.A3(n_202),
.B1(n_204),
.B2(n_208),
.C(n_195),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_227),
.A2(n_233),
.B1(n_219),
.B2(n_225),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_224),
.B(n_208),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_230),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_220),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_206),
.C(n_196),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_215),
.C(n_225),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_210),
.B(n_216),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_234),
.B(n_235),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_211),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_213),
.C(n_218),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_244),
.C(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_221),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_245),
.A2(n_218),
.B1(n_232),
.B2(n_203),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_248),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_240),
.B(n_242),
.Y(n_254)
);

OAI31xp33_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_233),
.A3(n_194),
.B(n_134),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_194),
.B(n_108),
.Y(n_255)
);

AOI21x1_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_252),
.B(n_250),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_255),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_238),
.B(n_241),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_257),
.B(n_126),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_244),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_258),
.A2(n_259),
.B(n_137),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_252),
.C(n_148),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_261),
.B(n_142),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_262),
.A2(n_263),
.B(n_260),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_142),
.Y(n_265)
);


endmodule