module real_aes_6482_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_1), .A2(n_150), .B(n_162), .C(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g269 ( .A(n_2), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_3), .A2(n_177), .B(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_4), .B(n_173), .Y(n_506) );
AOI21xp33_ASAP7_75t_L g176 ( .A1(n_5), .A2(n_177), .B(n_178), .Y(n_176) );
AND2x6_ASAP7_75t_L g150 ( .A(n_6), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_7), .A2(n_245), .B(n_246), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_8), .B(n_42), .Y(n_114) );
INVx1_ASAP7_75t_L g477 ( .A(n_9), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_10), .B(n_183), .Y(n_465) );
INVx1_ASAP7_75t_L g185 ( .A(n_11), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_12), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g147 ( .A(n_13), .Y(n_147) );
INVx1_ASAP7_75t_L g251 ( .A(n_14), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_15), .A2(n_186), .B(n_252), .C(n_486), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_16), .A2(n_128), .B1(n_129), .B2(n_130), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_16), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_17), .B(n_173), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_18), .A2(n_104), .B1(n_115), .B2(n_737), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_19), .B(n_196), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_20), .B(n_177), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_21), .B(n_519), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_22), .A2(n_153), .B(n_237), .C(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_23), .B(n_173), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_24), .B(n_183), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_25), .A2(n_249), .B(n_250), .C(n_252), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_26), .B(n_183), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_27), .Y(n_536) );
INVx1_ASAP7_75t_L g526 ( .A(n_28), .Y(n_526) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_29), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_30), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_31), .B(n_183), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_32), .A2(n_66), .B1(n_733), .B2(n_734), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_32), .Y(n_734) );
INVx1_ASAP7_75t_L g515 ( .A(n_33), .Y(n_515) );
INVx1_ASAP7_75t_L g161 ( .A(n_34), .Y(n_161) );
INVx2_ASAP7_75t_L g155 ( .A(n_35), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_36), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_37), .A2(n_187), .B(n_237), .C(n_504), .Y(n_503) );
INVxp67_ASAP7_75t_L g516 ( .A(n_38), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_39), .A2(n_150), .B(n_162), .C(n_207), .Y(n_206) );
CKINVDCx14_ASAP7_75t_R g502 ( .A(n_40), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_41), .A2(n_162), .B(n_525), .C(n_529), .Y(n_524) );
INVx1_ASAP7_75t_L g159 ( .A(n_43), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_44), .A2(n_182), .B(n_212), .C(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_45), .B(n_183), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_46), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_47), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_48), .Y(n_512) );
INVx1_ASAP7_75t_L g492 ( .A(n_49), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_50), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_51), .B(n_177), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_52), .A2(n_153), .B1(n_156), .B2(n_162), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_53), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g266 ( .A(n_54), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_55), .A2(n_182), .B(n_184), .C(n_187), .Y(n_181) );
CKINVDCx14_ASAP7_75t_R g474 ( .A(n_56), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_57), .Y(n_226) );
INVx1_ASAP7_75t_L g179 ( .A(n_58), .Y(n_179) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_59), .A2(n_731), .B1(n_732), .B2(n_735), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_59), .Y(n_735) );
INVx1_ASAP7_75t_L g151 ( .A(n_60), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_61), .A2(n_77), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_61), .Y(n_132) );
INVx1_ASAP7_75t_L g146 ( .A(n_62), .Y(n_146) );
INVx1_ASAP7_75t_SL g505 ( .A(n_63), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_64), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_65), .B(n_173), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_66), .Y(n_733) );
INVx1_ASAP7_75t_L g539 ( .A(n_67), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_SL g195 ( .A1(n_68), .A2(n_187), .B(n_196), .C(n_197), .Y(n_195) );
INVxp67_ASAP7_75t_L g198 ( .A(n_69), .Y(n_198) );
INVx1_ASAP7_75t_L g108 ( .A(n_70), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_71), .A2(n_177), .B(n_473), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_72), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_73), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_74), .A2(n_177), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g219 ( .A(n_75), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_76), .A2(n_245), .B(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_77), .Y(n_131) );
INVx1_ASAP7_75t_L g484 ( .A(n_78), .Y(n_484) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_79), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_80), .A2(n_150), .B(n_162), .C(n_221), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_81), .A2(n_177), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g487 ( .A(n_82), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_83), .B(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
INVx1_ASAP7_75t_L g463 ( .A(n_85), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_86), .B(n_196), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_87), .A2(n_150), .B(n_162), .C(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g110 ( .A(n_88), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g450 ( .A(n_88), .Y(n_450) );
OR2x2_ASAP7_75t_L g718 ( .A(n_88), .B(n_112), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_89), .A2(n_162), .B(n_538), .C(n_541), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_90), .B(n_190), .Y(n_189) );
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_91), .A2(n_126), .B1(n_127), .B2(n_133), .C1(n_719), .C2(n_723), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_92), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_93), .A2(n_150), .B(n_162), .C(n_234), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_94), .Y(n_241) );
INVx1_ASAP7_75t_L g194 ( .A(n_95), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_96), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_97), .B(n_209), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_98), .B(n_175), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_99), .B(n_175), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_100), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_101), .A2(n_177), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g495 ( .A(n_102), .Y(n_495) );
INVx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g738 ( .A(n_105), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_110), .Y(n_123) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_110), .Y(n_736) );
NOR2x2_ASAP7_75t_L g725 ( .A(n_111), .B(n_450), .Y(n_725) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g449 ( .A(n_112), .B(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_125), .B1(n_726), .B2(n_727), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_SL g726 ( .A(n_120), .Y(n_726) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_122), .A2(n_728), .B(n_736), .Y(n_727) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
CKINVDCx14_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_447), .B1(n_451), .B2(n_718), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g719 ( .A1(n_135), .A2(n_447), .B1(n_720), .B2(n_721), .Y(n_719) );
AND3x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_372), .C(n_421), .Y(n_135) );
NOR3xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_279), .C(n_317), .Y(n_136) );
OAI222xp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_200), .B1(n_254), .B2(n_260), .C1(n_274), .C2(n_277), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_171), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_139), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_139), .B(n_322), .Y(n_413) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g290 ( .A(n_140), .B(n_191), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_140), .B(n_172), .Y(n_298) );
AND2x2_ASAP7_75t_L g333 ( .A(n_140), .B(n_310), .Y(n_333) );
OR2x2_ASAP7_75t_L g357 ( .A(n_140), .B(n_172), .Y(n_357) );
OR2x2_ASAP7_75t_L g365 ( .A(n_140), .B(n_264), .Y(n_365) );
AND2x2_ASAP7_75t_L g368 ( .A(n_140), .B(n_191), .Y(n_368) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g262 ( .A(n_141), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g276 ( .A(n_141), .B(n_191), .Y(n_276) );
AND2x2_ASAP7_75t_L g326 ( .A(n_141), .B(n_264), .Y(n_326) );
AND2x2_ASAP7_75t_L g339 ( .A(n_141), .B(n_172), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_141), .B(n_425), .Y(n_446) );
AO21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_148), .B(n_169), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_142), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g214 ( .A(n_142), .Y(n_214) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_142), .A2(n_265), .B(n_272), .Y(n_264) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_143), .Y(n_175) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_144), .B(n_145), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .B1(n_165), .B2(n_166), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_149), .A2(n_179), .B(n_180), .C(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_149), .A2(n_180), .B(n_194), .C(n_195), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_149), .A2(n_180), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_SL g473 ( .A1(n_149), .A2(n_180), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_SL g483 ( .A1(n_149), .A2(n_180), .B(n_484), .C(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_SL g491 ( .A1(n_149), .A2(n_180), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_149), .A2(n_180), .B(n_502), .C(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_SL g511 ( .A1(n_149), .A2(n_180), .B(n_512), .C(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g541 ( .A(n_149), .Y(n_541) );
INVx4_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_150), .B(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g177 ( .A(n_150), .B(n_167), .Y(n_177) );
BUFx3_ASAP7_75t_L g529 ( .A(n_150), .Y(n_529) );
INVx2_ASAP7_75t_L g271 ( .A(n_153), .Y(n_271) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
INVx1_ASAP7_75t_L g168 ( .A(n_155), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g156 ( .A1(n_157), .A2(n_159), .B1(n_160), .B2(n_161), .Y(n_156) );
INVx2_ASAP7_75t_L g160 ( .A(n_157), .Y(n_160) );
INVx4_ASAP7_75t_L g249 ( .A(n_157), .Y(n_249) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
AND2x2_ASAP7_75t_L g167 ( .A(n_158), .B(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
INVx3_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
INVx1_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
INVx2_ASAP7_75t_L g464 ( .A(n_160), .Y(n_464) );
INVx5_ASAP7_75t_L g180 ( .A(n_162), .Y(n_180) );
AND2x6_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
BUFx3_ASAP7_75t_L g213 ( .A(n_163), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_166), .A2(n_219), .B(n_220), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_166), .A2(n_266), .B(n_267), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_166), .A2(n_460), .B(n_461), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_166), .A2(n_190), .B(n_523), .C(n_524), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_166), .A2(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g517 ( .A(n_168), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g364 ( .A1(n_171), .A2(n_365), .B(n_366), .C(n_369), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_171), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_171), .B(n_309), .Y(n_431) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_191), .Y(n_171) );
AND2x2_ASAP7_75t_SL g275 ( .A(n_172), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g289 ( .A(n_172), .Y(n_289) );
AND2x2_ASAP7_75t_L g316 ( .A(n_172), .B(n_310), .Y(n_316) );
INVx1_ASAP7_75t_SL g324 ( .A(n_172), .Y(n_324) );
AND2x2_ASAP7_75t_L g347 ( .A(n_172), .B(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g425 ( .A(n_172), .Y(n_425) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B(n_189), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_SL g215 ( .A(n_174), .B(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_174), .B(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_174), .B(n_531), .Y(n_530) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_174), .A2(n_535), .B(n_542), .Y(n_534) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_175), .A2(n_192), .B(n_199), .Y(n_191) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_175), .Y(n_481) );
BUFx2_ASAP7_75t_L g245 ( .A(n_177), .Y(n_245) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx4_ASAP7_75t_L g237 ( .A(n_183), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_186), .B(n_198), .Y(n_197) );
INVx5_ASAP7_75t_L g209 ( .A(n_186), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_186), .B(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_188), .Y(n_238) );
INVx1_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
INVx2_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_190), .A2(n_244), .B(n_253), .Y(n_243) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_190), .A2(n_472), .B(n_478), .Y(n_471) );
BUFx2_ASAP7_75t_L g261 ( .A(n_191), .Y(n_261) );
INVx1_ASAP7_75t_L g323 ( .A(n_191), .Y(n_323) );
INVx3_ASAP7_75t_L g348 ( .A(n_191), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_200), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_228), .Y(n_200) );
INVx1_ASAP7_75t_L g344 ( .A(n_201), .Y(n_344) );
OAI32xp33_ASAP7_75t_L g350 ( .A1(n_201), .A2(n_289), .A3(n_351), .B1(n_352), .B2(n_353), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_201), .A2(n_355), .B1(n_358), .B2(n_363), .Y(n_354) );
INVx4_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g292 ( .A(n_202), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g370 ( .A(n_202), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g440 ( .A(n_202), .B(n_386), .Y(n_440) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_217), .Y(n_202) );
AND2x2_ASAP7_75t_L g255 ( .A(n_203), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g285 ( .A(n_203), .Y(n_285) );
INVx1_ASAP7_75t_L g304 ( .A(n_203), .Y(n_304) );
OR2x2_ASAP7_75t_L g312 ( .A(n_203), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g319 ( .A(n_203), .B(n_293), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_203), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g340 ( .A(n_203), .B(n_258), .Y(n_340) );
INVx3_ASAP7_75t_L g362 ( .A(n_203), .Y(n_362) );
AND2x2_ASAP7_75t_L g387 ( .A(n_203), .B(n_259), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_203), .B(n_352), .Y(n_435) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_215), .Y(n_203) );
AOI21xp5_ASAP7_75t_SL g204 ( .A1(n_205), .A2(n_206), .B(n_214), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_210), .B(n_211), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_209), .A2(n_269), .B(n_270), .C(n_271), .Y(n_268) );
OAI22xp33_ASAP7_75t_L g514 ( .A1(n_209), .A2(n_249), .B1(n_515), .B2(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_209), .A2(n_526), .B(n_527), .C(n_528), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_211), .A2(n_222), .B(n_223), .Y(n_221) );
O2A1O1Ixp5_ASAP7_75t_L g462 ( .A1(n_211), .A2(n_463), .B(n_464), .C(n_465), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g538 ( .A1(n_211), .A2(n_464), .B(n_539), .C(n_540), .Y(n_538) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g252 ( .A(n_213), .Y(n_252) );
INVx1_ASAP7_75t_L g224 ( .A(n_214), .Y(n_224) );
INVx2_ASAP7_75t_L g259 ( .A(n_217), .Y(n_259) );
AND2x2_ASAP7_75t_L g391 ( .A(n_217), .B(n_229), .Y(n_391) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_224), .B(n_225), .Y(n_217) );
INVx1_ASAP7_75t_L g509 ( .A(n_224), .Y(n_509) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_224), .A2(n_562), .B(n_563), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_227), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_227), .B(n_273), .Y(n_272) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_227), .A2(n_459), .B(n_466), .Y(n_458) );
INVx2_ASAP7_75t_L g433 ( .A(n_228), .Y(n_433) );
OR2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_242), .Y(n_228) );
INVx1_ASAP7_75t_L g278 ( .A(n_229), .Y(n_278) );
AND2x2_ASAP7_75t_L g305 ( .A(n_229), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_229), .B(n_259), .Y(n_313) );
AND2x2_ASAP7_75t_L g371 ( .A(n_229), .B(n_294), .Y(n_371) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g257 ( .A(n_230), .Y(n_257) );
AND2x2_ASAP7_75t_L g284 ( .A(n_230), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g293 ( .A(n_230), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_230), .B(n_259), .Y(n_359) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_240), .Y(n_230) );
INVx1_ASAP7_75t_L g519 ( .A(n_231), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_231), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_239), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_238), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_237), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_242), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_242), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_242), .B(n_259), .Y(n_352) );
AND2x2_ASAP7_75t_L g361 ( .A(n_242), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g386 ( .A(n_242), .Y(n_386) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g258 ( .A(n_243), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g294 ( .A(n_243), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_249), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_249), .B(n_487), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_249), .B(n_495), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_254), .A2(n_264), .B1(n_423), .B2(n_426), .Y(n_422) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
OAI21xp5_ASAP7_75t_SL g445 ( .A1(n_256), .A2(n_367), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_257), .B(n_362), .Y(n_379) );
INVx1_ASAP7_75t_L g404 ( .A(n_257), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_258), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g331 ( .A(n_258), .B(n_284), .Y(n_331) );
INVx2_ASAP7_75t_L g287 ( .A(n_259), .Y(n_287) );
INVx1_ASAP7_75t_L g337 ( .A(n_259), .Y(n_337) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_260), .A2(n_412), .B1(n_429), .B2(n_432), .C(n_434), .Y(n_428) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g299 ( .A(n_261), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_261), .B(n_310), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_262), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g353 ( .A(n_262), .B(n_299), .Y(n_353) );
INVx3_ASAP7_75t_SL g394 ( .A(n_262), .Y(n_394) );
AND2x2_ASAP7_75t_L g338 ( .A(n_263), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g367 ( .A(n_263), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_263), .B(n_276), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_263), .B(n_322), .Y(n_408) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx3_ASAP7_75t_L g310 ( .A(n_264), .Y(n_310) );
OAI322xp33_ASAP7_75t_L g405 ( .A1(n_264), .A2(n_336), .A3(n_358), .B1(n_406), .B2(n_408), .C1(n_409), .C2(n_410), .Y(n_405) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI21xp33_ASAP7_75t_L g429 ( .A1(n_275), .A2(n_278), .B(n_430), .Y(n_429) );
NOR2xp33_ASAP7_75t_SL g355 ( .A(n_276), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g377 ( .A(n_276), .B(n_289), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_276), .B(n_316), .Y(n_392) );
INVxp67_ASAP7_75t_L g343 ( .A(n_278), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g349 ( .A1(n_278), .A2(n_350), .B(n_354), .C(n_364), .Y(n_349) );
OAI221xp5_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_288), .B1(n_291), .B2(n_295), .C(n_300), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g303 ( .A(n_287), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g420 ( .A(n_287), .Y(n_420) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_288), .A2(n_437), .B1(n_442), .B2(n_443), .C(n_445), .Y(n_436) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_289), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g336 ( .A(n_289), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_289), .B(n_367), .Y(n_374) );
AND2x2_ASAP7_75t_L g416 ( .A(n_289), .B(n_394), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_290), .B(n_315), .Y(n_314) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_290), .A2(n_302), .B1(n_412), .B2(n_413), .Y(n_411) );
OR2x2_ASAP7_75t_L g442 ( .A(n_290), .B(n_310), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g419 ( .A(n_293), .Y(n_419) );
AND2x2_ASAP7_75t_L g444 ( .A(n_293), .B(n_387), .Y(n_444) );
INVxp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_SL g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g308 ( .A(n_298), .B(n_309), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_307), .B1(n_311), .B2(n_314), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g375 ( .A(n_303), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_303), .B(n_343), .Y(n_410) );
AOI322xp5_ASAP7_75t_L g334 ( .A1(n_305), .A2(n_335), .A3(n_337), .B1(n_338), .B2(n_340), .C1(n_341), .C2(n_345), .Y(n_334) );
INVxp67_ASAP7_75t_L g328 ( .A(n_306), .Y(n_328) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_308), .A2(n_313), .B1(n_330), .B2(n_332), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_309), .B(n_322), .Y(n_409) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_310), .B(n_348), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_310), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g406 ( .A(n_312), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
NAND3xp33_ASAP7_75t_SL g317 ( .A(n_318), .B(n_334), .C(n_349), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B1(n_325), .B2(n_327), .C(n_329), .Y(n_318) );
AND2x2_ASAP7_75t_L g325 ( .A(n_321), .B(n_326), .Y(n_325) );
INVx3_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g335 ( .A(n_326), .B(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_328), .Y(n_407) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_333), .B(n_347), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_336), .B(n_394), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_337), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g412 ( .A(n_340), .Y(n_412) );
AND2x2_ASAP7_75t_L g427 ( .A(n_340), .B(n_404), .Y(n_427) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI211xp5_ASAP7_75t_L g421 ( .A1(n_351), .A2(n_422), .B(n_428), .C(n_436), .Y(n_421) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g390 ( .A(n_361), .B(n_391), .Y(n_390) );
NAND2x1_ASAP7_75t_SL g432 ( .A(n_362), .B(n_433), .Y(n_432) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_365), .Y(n_402) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g397 ( .A(n_371), .Y(n_397) );
AND2x2_ASAP7_75t_L g401 ( .A(n_371), .B(n_387), .Y(n_401) );
NOR5xp2_ASAP7_75t_L g372 ( .A(n_373), .B(n_388), .C(n_405), .D(n_411), .E(n_414), .Y(n_372) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_376), .B2(n_378), .C(n_380), .Y(n_373) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_377), .B(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g403 ( .A(n_387), .B(n_404), .Y(n_403) );
OAI221xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_392), .B1(n_393), .B2(n_395), .C(n_398), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g441 ( .A(n_401), .Y(n_441) );
AOI211xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_417), .B(n_419), .C(n_420), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
CKINVDCx14_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g720 ( .A(n_451), .Y(n_720) );
XNOR2xp5_ASAP7_75t_L g729 ( .A(n_451), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_SL g451 ( .A(n_452), .B(n_673), .Y(n_451) );
NAND5xp2_ASAP7_75t_L g452 ( .A(n_453), .B(n_585), .C(n_623), .D(n_644), .E(n_661), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_557), .C(n_578), .Y(n_453) );
OAI221xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_497), .B1(n_520), .B2(n_544), .C(n_548), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_468), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_457), .B(n_546), .Y(n_565) );
OR2x2_ASAP7_75t_L g592 ( .A(n_457), .B(n_480), .Y(n_592) );
AND2x2_ASAP7_75t_L g606 ( .A(n_457), .B(n_480), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_457), .B(n_471), .Y(n_620) );
AND2x2_ASAP7_75t_L g658 ( .A(n_457), .B(n_622), .Y(n_658) );
AND2x2_ASAP7_75t_L g687 ( .A(n_457), .B(n_597), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_457), .B(n_569), .Y(n_704) );
INVx4_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g584 ( .A(n_458), .B(n_479), .Y(n_584) );
BUFx3_ASAP7_75t_L g609 ( .A(n_458), .Y(n_609) );
AND2x2_ASAP7_75t_L g638 ( .A(n_458), .B(n_480), .Y(n_638) );
AND3x2_ASAP7_75t_L g651 ( .A(n_458), .B(n_652), .C(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g574 ( .A(n_468), .Y(n_574) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_479), .Y(n_468) );
AOI32xp33_ASAP7_75t_L g629 ( .A1(n_469), .A2(n_581), .A3(n_630), .B1(n_633), .B2(n_634), .Y(n_629) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g556 ( .A(n_470), .B(n_479), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_470), .B(n_584), .Y(n_627) );
AND2x2_ASAP7_75t_L g634 ( .A(n_470), .B(n_606), .Y(n_634) );
OR2x2_ASAP7_75t_L g640 ( .A(n_470), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_470), .B(n_595), .Y(n_665) );
OR2x2_ASAP7_75t_L g683 ( .A(n_470), .B(n_508), .Y(n_683) );
BUFx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g547 ( .A(n_471), .B(n_489), .Y(n_547) );
INVx2_ASAP7_75t_L g569 ( .A(n_471), .Y(n_569) );
OR2x2_ASAP7_75t_L g591 ( .A(n_471), .B(n_489), .Y(n_591) );
AND2x2_ASAP7_75t_L g596 ( .A(n_471), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_471), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g652 ( .A(n_471), .B(n_546), .Y(n_652) );
INVx1_ASAP7_75t_SL g703 ( .A(n_479), .Y(n_703) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_489), .Y(n_479) );
INVx1_ASAP7_75t_SL g546 ( .A(n_480), .Y(n_546) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_480), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_480), .B(n_632), .Y(n_631) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_480), .B(n_569), .C(n_687), .Y(n_698) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_488), .Y(n_480) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_481), .A2(n_490), .B(n_496), .Y(n_489) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_481), .A2(n_500), .B(n_506), .Y(n_499) );
INVx2_ASAP7_75t_L g597 ( .A(n_489), .Y(n_597) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_489), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
INVx1_ASAP7_75t_L g633 ( .A(n_498), .Y(n_633) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g551 ( .A(n_499), .B(n_533), .Y(n_551) );
INVx2_ASAP7_75t_L g568 ( .A(n_499), .Y(n_568) );
AND2x2_ASAP7_75t_L g573 ( .A(n_499), .B(n_534), .Y(n_573) );
AND2x2_ASAP7_75t_L g588 ( .A(n_499), .B(n_521), .Y(n_588) );
AND2x2_ASAP7_75t_L g600 ( .A(n_499), .B(n_572), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_507), .B(n_616), .Y(n_615) );
NAND2x1p5_ASAP7_75t_L g672 ( .A(n_507), .B(n_573), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_507), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_507), .B(n_567), .Y(n_695) );
BUFx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g532 ( .A(n_508), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_508), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g577 ( .A(n_508), .B(n_521), .Y(n_577) );
AND2x2_ASAP7_75t_L g603 ( .A(n_508), .B(n_533), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_508), .B(n_643), .Y(n_642) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_518), .Y(n_508) );
INVx1_ASAP7_75t_L g562 ( .A(n_510), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_514), .B(n_517), .Y(n_513) );
INVx2_ASAP7_75t_L g528 ( .A(n_517), .Y(n_528) );
INVx1_ASAP7_75t_L g563 ( .A(n_518), .Y(n_563) );
OR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_532), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_521), .B(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g567 ( .A(n_521), .B(n_568), .Y(n_567) );
INVx3_ASAP7_75t_SL g572 ( .A(n_521), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_521), .B(n_559), .Y(n_625) );
OR2x2_ASAP7_75t_L g635 ( .A(n_521), .B(n_561), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_521), .B(n_603), .Y(n_663) );
OR2x2_ASAP7_75t_L g693 ( .A(n_521), .B(n_533), .Y(n_693) );
AND2x2_ASAP7_75t_L g697 ( .A(n_521), .B(n_534), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_521), .B(n_573), .Y(n_710) );
AND2x2_ASAP7_75t_L g717 ( .A(n_521), .B(n_599), .Y(n_717) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_530), .Y(n_521) );
INVx1_ASAP7_75t_SL g660 ( .A(n_532), .Y(n_660) );
AND2x2_ASAP7_75t_L g599 ( .A(n_533), .B(n_561), .Y(n_599) );
AND2x2_ASAP7_75t_L g613 ( .A(n_533), .B(n_568), .Y(n_613) );
AND2x2_ASAP7_75t_L g616 ( .A(n_533), .B(n_572), .Y(n_616) );
INVx1_ASAP7_75t_L g643 ( .A(n_533), .Y(n_643) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_L g555 ( .A(n_534), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g714 ( .A1(n_545), .A2(n_591), .B(n_715), .C(n_716), .Y(n_714) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g621 ( .A(n_546), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_547), .B(n_564), .Y(n_579) );
AND2x2_ASAP7_75t_L g605 ( .A(n_547), .B(n_606), .Y(n_605) );
OAI21xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_552), .B(n_556), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_550), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g576 ( .A(n_551), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_551), .B(n_572), .Y(n_617) );
AND2x2_ASAP7_75t_L g708 ( .A(n_551), .B(n_559), .Y(n_708) );
INVxp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g581 ( .A(n_555), .B(n_568), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_555), .B(n_566), .Y(n_582) );
OAI322xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_565), .A3(n_566), .B1(n_569), .B2(n_570), .C1(n_574), .C2(n_575), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_564), .Y(n_558) );
AND2x2_ASAP7_75t_L g669 ( .A(n_559), .B(n_581), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_559), .B(n_633), .Y(n_715) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g612 ( .A(n_561), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g678 ( .A(n_565), .B(n_591), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_566), .B(n_660), .Y(n_659) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_567), .B(n_599), .Y(n_656) );
AND2x2_ASAP7_75t_L g602 ( .A(n_568), .B(n_572), .Y(n_602) );
AND2x2_ASAP7_75t_L g610 ( .A(n_569), .B(n_611), .Y(n_610) );
A2O1A1Ixp33_ASAP7_75t_L g707 ( .A1(n_569), .A2(n_648), .B(n_708), .C(n_709), .Y(n_707) );
AOI21xp33_ASAP7_75t_L g680 ( .A1(n_570), .A2(n_583), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_572), .B(n_599), .Y(n_639) );
AND2x2_ASAP7_75t_L g645 ( .A(n_572), .B(n_613), .Y(n_645) );
AND2x2_ASAP7_75t_L g679 ( .A(n_572), .B(n_581), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_573), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_SL g689 ( .A(n_573), .Y(n_689) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_577), .A2(n_605), .B1(n_607), .B2(n_612), .Y(n_604) );
OAI22xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_580), .B1(n_582), .B2(n_583), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g614 ( .A1(n_579), .A2(n_615), .B1(n_617), .B2(n_618), .Y(n_614) );
INVxp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_584), .A2(n_686), .B1(n_688), .B2(n_690), .C(n_694), .Y(n_685) );
AOI211xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_589), .B(n_593), .C(n_614), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
OR2x2_ASAP7_75t_L g655 ( .A(n_591), .B(n_608), .Y(n_655) );
INVx1_ASAP7_75t_L g706 ( .A(n_591), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_592), .A2(n_594), .B1(n_598), .B2(n_601), .C(n_604), .Y(n_593) );
INVx2_ASAP7_75t_SL g648 ( .A(n_592), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g713 ( .A(n_595), .Y(n_713) );
AND2x2_ASAP7_75t_L g637 ( .A(n_596), .B(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g622 ( .A(n_597), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g684 ( .A(n_600), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_608), .B(n_710), .Y(n_709) );
CKINVDCx16_ASAP7_75t_R g608 ( .A(n_609), .Y(n_608) );
INVxp67_ASAP7_75t_L g653 ( .A(n_611), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_612), .A2(n_624), .B(n_626), .C(n_628), .Y(n_623) );
INVx1_ASAP7_75t_L g701 ( .A(n_615), .Y(n_701) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_619), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g632 ( .A(n_622), .Y(n_632) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI222xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_635), .B1(n_636), .B2(n_639), .C1(n_640), .C2(n_642), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g668 ( .A(n_632), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_635), .B(n_689), .Y(n_688) );
NAND2xp33_ASAP7_75t_SL g666 ( .A(n_636), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g641 ( .A(n_638), .Y(n_641) );
AND2x2_ASAP7_75t_L g705 ( .A(n_638), .B(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g671 ( .A(n_641), .B(n_668), .Y(n_671) );
INVx1_ASAP7_75t_L g700 ( .A(n_642), .Y(n_700) );
AOI211xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B(n_649), .C(n_654), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_648), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
AOI322xp5_ASAP7_75t_L g699 ( .A1(n_651), .A2(n_679), .A3(n_684), .B1(n_700), .B2(n_701), .C1(n_702), .C2(n_705), .Y(n_699) );
AND2x2_ASAP7_75t_L g686 ( .A(n_652), .B(n_687), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B1(n_657), .B2(n_659), .Y(n_654) );
INVxp33_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_664), .B1(n_666), .B2(n_669), .C(n_670), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
NAND5xp2_ASAP7_75t_L g673 ( .A(n_674), .B(n_685), .C(n_699), .D(n_707), .E(n_711), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_679), .B(n_680), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVxp33_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g711 ( .A1(n_687), .A2(n_712), .B(n_713), .C(n_714), .Y(n_711) );
AOI31xp33_ASAP7_75t_L g694 ( .A1(n_689), .A2(n_695), .A3(n_696), .B(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g712 ( .A(n_710), .Y(n_712) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g722 ( .A(n_718), .Y(n_722) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
endmodule