module fake_netlist_1_4674_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
OA21x2_ASAP7_75t_L g12 ( .A1(n_3), .A2(n_0), .B(n_7), .Y(n_12) );
OR2x6_ASAP7_75t_L g13 ( .A(n_9), .B(n_1), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_13), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_13), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_18) );
OAI21x1_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_12), .B(n_11), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
BUFx3_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
HB1xp67_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_20), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_22), .B1(n_21), .B2(n_20), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
NOR2xp33_ASAP7_75t_L g27 ( .A(n_26), .B(n_17), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_14), .B1(n_13), .B2(n_12), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_28), .B(n_2), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_27), .B(n_14), .Y(n_30) );
OAI22xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_21), .B1(n_12), .B2(n_11), .Y(n_31) );
OAI22xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_11), .B1(n_19), .B2(n_10), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
OAI221xp5_ASAP7_75t_R g34 ( .A1(n_33), .A2(n_11), .B1(n_32), .B2(n_5), .C(n_8), .Y(n_34) );
endmodule