module fake_netlist_6_978_n_33 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_8, n_33);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_8;

output n_33;

wire n_16;
wire n_21;
wire n_24;
wire n_10;
wire n_18;
wire n_15;
wire n_27;
wire n_14;
wire n_32;
wire n_22;
wire n_26;
wire n_13;
wire n_11;
wire n_28;
wire n_23;
wire n_17;
wire n_12;
wire n_20;
wire n_30;
wire n_19;
wire n_29;
wire n_31;
wire n_25;

CKINVDCx5p33_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_6),
.B(n_2),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_16),
.A2(n_0),
.B(n_3),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_21),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

AOI222xp33_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_15),
.B1(n_10),
.B2(n_17),
.C1(n_25),
.C2(n_5),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_28),
.A2(n_19),
.B(n_18),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_29),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_15),
.B1(n_27),
.B2(n_5),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_31),
.B1(n_0),
.B2(n_3),
.Y(n_33)
);


endmodule