module fake_jpeg_6393_n_190 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_1),
.B(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_34),
.A2(n_38),
.B1(n_29),
.B2(n_31),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_1),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_2),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_42),
.B(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_45),
.Y(n_65)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_39),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_14),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_44)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_20),
.B1(n_5),
.B2(n_8),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_58),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_55),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_17),
.B1(n_15),
.B2(n_25),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_54),
.A2(n_57),
.B1(n_59),
.B2(n_64),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_44),
.B(n_41),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_17),
.B1(n_15),
.B2(n_25),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_26),
.B1(n_23),
.B2(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_69),
.Y(n_84)
);

CKINVDCx6p67_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_34),
.A2(n_26),
.B1(n_18),
.B2(n_28),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_72),
.B1(n_73),
.B2(n_78),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_20),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_76),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_38),
.A2(n_28),
.B1(n_27),
.B2(n_21),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_38),
.A2(n_20),
.B1(n_32),
.B2(n_29),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_36),
.A2(n_27),
.B1(n_21),
.B2(n_16),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_64),
.B1(n_55),
.B2(n_52),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_20),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_36),
.A2(n_32),
.B1(n_20),
.B2(n_19),
.Y(n_78)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_40),
.Y(n_97)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_48),
.B(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_93),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_48),
.B(n_19),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_62),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_4),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_99),
.B1(n_104),
.B2(n_73),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_67),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_20),
.B1(n_22),
.B2(n_9),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_22),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_22),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_4),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_49),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_22),
.B1(n_9),
.B2(n_10),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_106),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_82),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_101),
.B1(n_89),
.B2(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_111),
.Y(n_133)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_62),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_83),
.B(n_95),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_69),
.C(n_58),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_80),
.C(n_96),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_103),
.A2(n_73),
.B1(n_78),
.B2(n_53),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_116),
.B1(n_83),
.B2(n_95),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_71),
.B1(n_66),
.B2(n_56),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_56),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_94),
.Y(n_128)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_124),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_65),
.B(n_22),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_91),
.B(n_87),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_127),
.C(n_128),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_94),
.C(n_90),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_81),
.B(n_88),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_143),
.C(n_118),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_137),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_89),
.B1(n_104),
.B2(n_75),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_70),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_109),
.C(n_106),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_70),
.C(n_79),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_116),
.B1(n_115),
.B2(n_119),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_138),
.B(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_146),
.B(n_133),
.Y(n_163)
);

AO22x2_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_110),
.B1(n_123),
.B2(n_108),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_149),
.A2(n_126),
.B(n_129),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_121),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_105),
.C(n_117),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_147),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_127),
.C(n_130),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_160),
.A2(n_161),
.B(n_162),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_149),
.B(n_135),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_167),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_141),
.B(n_137),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_166),
.A2(n_151),
.B(n_148),
.Y(n_174)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_159),
.C(n_161),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_149),
.B1(n_142),
.B2(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_111),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_174),
.B(n_162),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_176),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_164),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_177),
.A2(n_140),
.B(n_111),
.C(n_125),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_180),
.B(n_172),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_140),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_175),
.B(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

AOI31xp67_ASAP7_75t_SL g183 ( 
.A1(n_177),
.A2(n_179),
.A3(n_176),
.B(n_125),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_13),
.B(n_8),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_186),
.A2(n_187),
.B(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_189),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_185),
.A2(n_13),
.B(n_8),
.Y(n_189)
);


endmodule