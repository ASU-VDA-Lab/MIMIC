module fake_jpeg_15023_n_196 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_196);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_39),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_31),
.B1(n_33),
.B2(n_21),
.Y(n_58)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_2),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_21),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_4),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_27),
.Y(n_68)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_45),
.B(n_46),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_5),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_5),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_49),
.Y(n_70)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_7),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_54),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

HAxp5_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_43),
.CON(n_69),
.SN(n_69)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_31),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_8),
.B(n_10),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_58),
.A2(n_60),
.B1(n_82),
.B2(n_75),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_29),
.B1(n_24),
.B2(n_20),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_26),
.B1(n_27),
.B2(n_25),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_20),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_24),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_17),
.B1(n_33),
.B2(n_22),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_66),
.B1(n_83),
.B2(n_13),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_17),
.B(n_10),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_87),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_34),
.B(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_78),
.B(n_63),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_80),
.Y(n_109)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_23),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_36),
.A2(n_47),
.B1(n_41),
.B2(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_23),
.Y(n_85)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_16),
.Y(n_86)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_52),
.B(n_25),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_66),
.B1(n_64),
.B2(n_80),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_26),
.B1(n_52),
.B2(n_54),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_103),
.B1(n_66),
.B2(n_86),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_109),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_11),
.C(n_12),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_95),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_11),
.C(n_12),
.Y(n_95)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_13),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_104),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_82),
.B1(n_74),
.B2(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_64),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_110),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_71),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_62),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_115),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_78),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_64),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_78),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_106),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_136),
.Y(n_140)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_66),
.A3(n_87),
.B1(n_83),
.B2(n_64),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_107),
.Y(n_146)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_129),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_126),
.A2(n_107),
.B1(n_114),
.B2(n_97),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_107),
.B(n_89),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_81),
.Y(n_129)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_135),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_91),
.A2(n_74),
.B1(n_83),
.B2(n_57),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_96),
.B(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_57),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_89),
.C(n_112),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_147),
.C(n_148),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_139),
.A2(n_127),
.B(n_117),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_135),
.B1(n_133),
.B2(n_127),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_145),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_120),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_97),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_108),
.C(n_100),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_108),
.C(n_100),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_153),
.C(n_137),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_116),
.C(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_101),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_155),
.B(n_119),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_149),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_101),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_162),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_129),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_126),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_165),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_166),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_148),
.C(n_153),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_168),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_93),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_141),
.B(n_144),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_171),
.B(n_163),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_152),
.B(n_139),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_147),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_176),
.C(n_159),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_154),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_97),
.C(n_94),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_179),
.A2(n_177),
.B(n_174),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_181),
.C(n_185),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_166),
.C(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_183),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_145),
.B1(n_134),
.B2(n_95),
.Y(n_183)
);

AO21x1_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_94),
.B(n_81),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_SL g188 ( 
.A1(n_184),
.A2(n_182),
.B(n_174),
.C(n_83),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_83),
.C(n_122),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_186),
.A2(n_188),
.B(n_189),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_170),
.B(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

OAI221xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_193),
.B1(n_187),
.B2(n_130),
.C(n_84),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_170),
.B1(n_142),
.B2(n_132),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_195),
.Y(n_196)
);

AOI321xp33_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_84),
.A3(n_88),
.B1(n_92),
.B2(n_130),
.C(n_191),
.Y(n_195)
);


endmodule