module fake_jpeg_11191_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_1),
.B(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_12),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_19),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_29),
.B1(n_21),
.B2(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_24),
.B1(n_15),
.B2(n_30),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_18),
.B1(n_28),
.B2(n_19),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_26),
.B1(n_38),
.B2(n_25),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_21),
.B1(n_23),
.B2(n_20),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_36),
.B1(n_29),
.B2(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_65),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_40),
.B1(n_18),
.B2(n_28),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_45),
.B1(n_38),
.B2(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_63),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_34),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_68),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_26),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_76),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_97),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_79),
.B(n_63),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_52),
.C(n_48),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_67),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_51),
.B1(n_38),
.B2(n_20),
.Y(n_116)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_65),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_20),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_65),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_68),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_114),
.C(n_83),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_20),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_73),
.B(n_75),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_57),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_76),
.B1(n_78),
.B2(n_45),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_116),
.B1(n_95),
.B2(n_91),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_66),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_1),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_123),
.B(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_89),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_133),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_101),
.B1(n_108),
.B2(n_85),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_82),
.B1(n_95),
.B2(n_91),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_84),
.B1(n_113),
.B2(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_98),
.B(n_94),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_134),
.B(n_93),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_86),
.C(n_99),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_98),
.B(n_94),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_138),
.Y(n_151)
);

OAI322xp33_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_88),
.A3(n_107),
.B1(n_112),
.B2(n_114),
.C1(n_104),
.C2(n_116),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_132),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_120),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_90),
.B1(n_100),
.B2(n_87),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_119),
.B(n_138),
.C(n_121),
.D(n_143),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_103),
.B1(n_25),
.B2(n_16),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_144),
.A2(n_145),
.B(n_134),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_120),
.Y(n_145)
);

XOR2x2_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_133),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_148),
.C(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_150),
.B(n_152),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_13),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_146),
.B1(n_144),
.B2(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_119),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_158),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_159),
.B(n_10),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_127),
.C(n_142),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_161),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_151),
.C(n_121),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_141),
.B(n_140),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_162),
.A2(n_103),
.B(n_25),
.C(n_3),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_149),
.B1(n_124),
.B2(n_122),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_1),
.B(n_2),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_165),
.A2(n_167),
.B1(n_10),
.B2(n_9),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_156),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.Y(n_172)
);

AOI21x1_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_167),
.B(n_9),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_5),
.B(n_6),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_173),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_176),
.B(n_172),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_6),
.A3(n_7),
.B1(n_16),
.B2(n_17),
.C1(n_154),
.C2(n_159),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_7),
.Y(n_179)
);


endmodule