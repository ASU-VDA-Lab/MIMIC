module fake_aes_6694_n_948 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_948);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_948;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_622;
wire n_549;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_14), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_60), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_91), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_34), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_5), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_19), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_67), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_71), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_57), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_101), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_103), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_72), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_26), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_48), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_80), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_40), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_85), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_66), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_45), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_99), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_47), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_59), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_95), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_90), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_83), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_89), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_35), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_31), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_22), .Y(n_139) );
INVx1_ASAP7_75t_SL g140 ( .A(n_6), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_17), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_96), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_55), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_4), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_69), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_100), .Y(n_146) );
NOR2xp67_ASAP7_75t_L g147 ( .A(n_33), .B(n_43), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_0), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_78), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_65), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_41), .Y(n_151) );
INVx5_ASAP7_75t_L g152 ( .A(n_136), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_115), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_136), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_136), .B(n_0), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_127), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g157 ( .A1(n_110), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_125), .B(n_1), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_127), .B(n_2), .Y(n_159) );
BUFx12f_ASAP7_75t_L g160 ( .A(n_111), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_139), .Y(n_162) );
INVxp67_ASAP7_75t_L g163 ( .A(n_114), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_113), .B(n_23), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_110), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_127), .Y(n_166) );
BUFx12f_ASAP7_75t_L g167 ( .A(n_111), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_113), .B(n_3), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_144), .B(n_4), .Y(n_169) );
AND2x6_ASAP7_75t_L g170 ( .A(n_112), .B(n_24), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_142), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_144), .B(n_5), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_127), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_127), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_142), .B(n_6), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_165), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_162), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_160), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_160), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_152), .B(n_149), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_167), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_155), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_167), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_171), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
NOR2xp33_ASAP7_75t_R g188 ( .A(n_175), .B(n_149), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_168), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_168), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_175), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_163), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_169), .Y(n_194) );
NOR2xp33_ASAP7_75t_R g195 ( .A(n_152), .B(n_151), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_168), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_172), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_158), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_168), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_152), .B(n_116), .Y(n_201) );
NOR2xp67_ASAP7_75t_L g202 ( .A(n_152), .B(n_128), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_157), .Y(n_203) );
NAND2xp33_ASAP7_75t_R g204 ( .A(n_153), .B(n_141), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_157), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_174), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_153), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_161), .Y(n_208) );
INVxp67_ASAP7_75t_L g209 ( .A(n_161), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_154), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_159), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_154), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_154), .Y(n_213) );
NOR2xp33_ASAP7_75t_R g214 ( .A(n_170), .B(n_151), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_174), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_170), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_170), .B(n_140), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_174), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_170), .Y(n_219) );
AOI21x1_ASAP7_75t_L g220 ( .A1(n_164), .A2(n_150), .B(n_146), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_156), .Y(n_221) );
CKINVDCx16_ASAP7_75t_R g222 ( .A(n_170), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_173), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_170), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_170), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_164), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_208), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_222), .B(n_130), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_184), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_199), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_199), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_199), .Y(n_232) );
INVxp33_ASAP7_75t_L g233 ( .A(n_188), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_219), .B(n_143), .Y(n_234) );
INVxp67_ASAP7_75t_L g235 ( .A(n_192), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_176), .B(n_145), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_210), .B(n_117), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_193), .Y(n_238) );
INVx2_ASAP7_75t_SL g239 ( .A(n_184), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_194), .B(n_118), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_197), .B(n_119), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_198), .B(n_120), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_214), .B(n_147), .Y(n_243) );
NOR3xp33_ASAP7_75t_L g244 ( .A(n_205), .B(n_121), .C(n_122), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_212), .B(n_148), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_213), .B(n_123), .Y(n_246) );
INVxp67_ASAP7_75t_L g247 ( .A(n_204), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_207), .B(n_124), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_209), .B(n_126), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_189), .B(n_190), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_186), .Y(n_251) );
INVx2_ASAP7_75t_SL g252 ( .A(n_180), .Y(n_252) );
INVx1_ASAP7_75t_SL g253 ( .A(n_186), .Y(n_253) );
NOR3xp33_ASAP7_75t_L g254 ( .A(n_191), .B(n_129), .C(n_131), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_196), .B(n_132), .Y(n_255) );
INVxp67_ASAP7_75t_L g256 ( .A(n_177), .Y(n_256) );
INVxp67_ASAP7_75t_L g257 ( .A(n_183), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_193), .Y(n_258) );
NOR3xp33_ASAP7_75t_L g259 ( .A(n_198), .B(n_133), .C(n_134), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_180), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_180), .B(n_135), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_225), .B(n_137), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_182), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_187), .B(n_138), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_201), .B(n_164), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_201), .B(n_164), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_201), .B(n_164), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_200), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_211), .B(n_164), .Y(n_269) );
NOR3xp33_ASAP7_75t_L g270 ( .A(n_183), .B(n_164), .C(n_8), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_195), .B(n_173), .Y(n_271) );
INVxp67_ASAP7_75t_SL g272 ( .A(n_216), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_217), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_217), .B(n_156), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_202), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_211), .B(n_25), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_185), .B(n_7), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_206), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_206), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_226), .B(n_156), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_181), .B(n_27), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_216), .A2(n_166), .B(n_156), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_224), .B(n_156), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_215), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_224), .B(n_173), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_185), .B(n_173), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_218), .Y(n_287) );
AO221x1_ASAP7_75t_L g288 ( .A1(n_203), .A2(n_173), .B1(n_166), .B2(n_156), .C(n_10), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_220), .B(n_166), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_178), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_278), .Y(n_291) );
O2A1O1Ixp33_ASAP7_75t_L g292 ( .A1(n_273), .A2(n_203), .B(n_223), .C(n_179), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_229), .B(n_166), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_236), .B(n_7), .Y(n_294) );
NAND2xp33_ASAP7_75t_L g295 ( .A(n_239), .B(n_166), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_278), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_227), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_269), .A2(n_166), .B1(n_223), .B2(n_221), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_251), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_260), .Y(n_300) );
BUFx8_ASAP7_75t_L g301 ( .A(n_245), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_236), .B(n_8), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_263), .B(n_9), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_250), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_229), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_229), .B(n_221), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_279), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_242), .A2(n_221), .B1(n_12), .B2(n_13), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_240), .B(n_11), .Y(n_310) );
INVx4_ASAP7_75t_SL g311 ( .A(n_229), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_241), .B(n_12), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_251), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_287), .Y(n_314) );
AND2x6_ASAP7_75t_L g315 ( .A(n_265), .B(n_221), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_239), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_230), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_248), .B(n_13), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_245), .A2(n_221), .B1(n_15), .B2(n_16), .C(n_17), .Y(n_319) );
INVx5_ASAP7_75t_L g320 ( .A(n_252), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_252), .B(n_109), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_287), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_238), .Y(n_323) );
NAND2x1p5_ASAP7_75t_L g324 ( .A(n_268), .B(n_14), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_231), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_235), .B(n_15), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_237), .B(n_16), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_246), .B(n_18), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_232), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_253), .B(n_18), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_256), .Y(n_331) );
NOR2x1p5_ASAP7_75t_L g332 ( .A(n_277), .B(n_19), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_257), .Y(n_333) );
O2A1O1Ixp5_ASAP7_75t_L g334 ( .A1(n_243), .A2(n_64), .B(n_107), .C(n_28), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_247), .B(n_20), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_238), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_233), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_284), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_233), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_254), .B(n_20), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_259), .B(n_21), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_297), .B(n_228), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_333), .B(n_272), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_314), .Y(n_344) );
AND2x6_ASAP7_75t_L g345 ( .A(n_316), .B(n_266), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_291), .A2(n_267), .B(n_274), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_307), .A2(n_289), .B(n_282), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_291), .A2(n_274), .B(n_234), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_331), .B(n_244), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_338), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_333), .B(n_290), .Y(n_351) );
INVx1_ASAP7_75t_SL g352 ( .A(n_299), .Y(n_352) );
NOR3xp33_ASAP7_75t_L g353 ( .A(n_292), .B(n_276), .C(n_228), .Y(n_353) );
AOI21x1_ASAP7_75t_L g354 ( .A1(n_321), .A2(n_243), .B(n_271), .Y(n_354) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_303), .A2(n_270), .B(n_275), .C(n_255), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_322), .Y(n_356) );
NAND3xp33_ASAP7_75t_SL g357 ( .A(n_319), .B(n_286), .C(n_249), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_314), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_313), .B(n_264), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g360 ( .A1(n_296), .A2(n_234), .B(n_258), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_301), .Y(n_361) );
XNOR2xp5_ASAP7_75t_L g362 ( .A(n_332), .B(n_262), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_300), .B(n_258), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_322), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_296), .A2(n_280), .B(n_261), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_317), .B(n_283), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_337), .B(n_283), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_294), .A2(n_285), .B1(n_262), .B2(n_280), .Y(n_368) );
OAI21xp33_ASAP7_75t_L g369 ( .A1(n_302), .A2(n_281), .B(n_288), .Y(n_369) );
AO32x2_ASAP7_75t_L g370 ( .A1(n_304), .A2(n_324), .A3(n_309), .B1(n_334), .B2(n_335), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_295), .A2(n_68), .B(n_29), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_325), .B(n_21), .Y(n_372) );
O2A1O1Ixp33_ASAP7_75t_L g373 ( .A1(n_341), .A2(n_30), .B(n_32), .C(n_36), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_356), .Y(n_374) );
AO21x2_ASAP7_75t_L g375 ( .A1(n_369), .A2(n_321), .B(n_327), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_356), .Y(n_376) );
AO21x2_ASAP7_75t_L g377 ( .A1(n_354), .A2(n_328), .B(n_318), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_363), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_350), .B(n_342), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_347), .A2(n_307), .B(n_293), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_344), .Y(n_381) );
NOR2xp67_ASAP7_75t_SL g382 ( .A(n_356), .B(n_322), .Y(n_382) );
AO21x2_ASAP7_75t_L g383 ( .A1(n_357), .A2(n_298), .B(n_293), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_358), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_364), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_361), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_349), .B(n_301), .Y(n_387) );
INVx1_ASAP7_75t_SL g388 ( .A(n_352), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_362), .Y(n_389) );
OAI21x1_ASAP7_75t_L g390 ( .A1(n_371), .A2(n_324), .B(n_310), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_363), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_364), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_366), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_366), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g395 ( .A1(n_355), .A2(n_305), .B(n_308), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_364), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_360), .B(n_311), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_345), .Y(n_398) );
NOR2x1_ASAP7_75t_SL g399 ( .A(n_372), .B(n_322), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_372), .Y(n_400) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_370), .Y(n_401) );
BUFx2_ASAP7_75t_SL g402 ( .A(n_345), .Y(n_402) );
OAI21x1_ASAP7_75t_L g403 ( .A1(n_371), .A2(n_312), .B(n_323), .Y(n_403) );
OAI21x1_ASAP7_75t_L g404 ( .A1(n_373), .A2(n_323), .B(n_305), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_386), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_379), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_376), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_404), .A2(n_365), .B(n_346), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_379), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_374), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_388), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_378), .Y(n_412) );
BUFx8_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_391), .A2(n_340), .B1(n_342), .B2(n_367), .Y(n_414) );
NAND2x1p5_ASAP7_75t_L g415 ( .A(n_382), .B(n_320), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_391), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_381), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_388), .B(n_340), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_398), .B(n_311), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_381), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_384), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_400), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_400), .A2(n_340), .B1(n_353), .B2(n_330), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_384), .B(n_308), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_393), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_387), .A2(n_301), .B1(n_335), .B2(n_359), .Y(n_426) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_382), .B(n_374), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_400), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_393), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_400), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_394), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_394), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_386), .Y(n_433) );
INVx1_ASAP7_75t_SL g434 ( .A(n_387), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_376), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_395), .B(n_370), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
INVx6_ASAP7_75t_L g438 ( .A(n_374), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_399), .Y(n_439) );
AOI21x1_ASAP7_75t_L g440 ( .A1(n_404), .A2(n_368), .B(n_348), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_389), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_399), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_374), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_385), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_402), .A2(n_343), .B1(n_316), .B2(n_326), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_380), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_402), .A2(n_351), .B1(n_339), .B2(n_329), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_390), .Y(n_448) );
CKINVDCx11_ASAP7_75t_R g449 ( .A(n_396), .Y(n_449) );
OAI21x1_ASAP7_75t_SL g450 ( .A1(n_398), .A2(n_370), .B(n_345), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_397), .A2(n_345), .B1(n_315), .B2(n_306), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_390), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_417), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_406), .B(n_390), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g455 ( .A(n_405), .Y(n_455) );
NOR2xp33_ASAP7_75t_R g456 ( .A(n_413), .B(n_398), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_413), .A2(n_401), .B1(n_402), .B2(n_375), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_422), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_420), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_405), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_434), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_411), .B(n_396), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_424), .B(n_392), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_424), .B(n_392), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_412), .Y(n_465) );
INVx4_ASAP7_75t_L g466 ( .A(n_449), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_422), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_421), .Y(n_468) );
INVxp33_ASAP7_75t_SL g469 ( .A(n_441), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_428), .Y(n_470) );
NOR2xp33_ASAP7_75t_R g471 ( .A(n_413), .B(n_392), .Y(n_471) );
AO31x2_ASAP7_75t_L g472 ( .A1(n_448), .A2(n_375), .A3(n_401), .B(n_377), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_412), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_423), .A2(n_403), .B(n_380), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_428), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_414), .A2(n_401), .B1(n_397), .B2(n_375), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_416), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_433), .B(n_392), .Y(n_478) );
BUFx10_ASAP7_75t_L g479 ( .A(n_441), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_409), .B(n_401), .Y(n_480) );
NAND2xp33_ASAP7_75t_R g481 ( .A(n_407), .B(n_397), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_415), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_449), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_418), .B(n_392), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_416), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_425), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_430), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_407), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_435), .B(n_397), .Y(n_489) );
AO32x2_ASAP7_75t_L g490 ( .A1(n_445), .A2(n_401), .A3(n_375), .B1(n_377), .B2(n_404), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_429), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_430), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_435), .Y(n_493) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_410), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_431), .B(n_385), .Y(n_495) );
INVxp33_ASAP7_75t_SL g496 ( .A(n_426), .Y(n_496) );
OR2x6_ASAP7_75t_L g497 ( .A(n_427), .B(n_397), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_432), .B(n_401), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_447), .B(n_401), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_446), .Y(n_500) );
NOR2xp33_ASAP7_75t_R g501 ( .A(n_443), .B(n_385), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_443), .B(n_401), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_439), .B(n_442), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_419), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_446), .Y(n_505) );
AOI21xp33_ASAP7_75t_L g506 ( .A1(n_452), .A2(n_375), .B(n_377), .Y(n_506) );
NOR2xp33_ASAP7_75t_R g507 ( .A(n_443), .B(n_385), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_451), .A2(n_320), .B1(n_306), .B2(n_323), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_438), .Y(n_509) );
NAND2x1_ASAP7_75t_L g510 ( .A(n_438), .B(n_382), .Y(n_510) );
NAND2xp33_ASAP7_75t_R g511 ( .A(n_436), .B(n_403), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_437), .A2(n_383), .B1(n_377), .B2(n_345), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_438), .Y(n_513) );
NOR2xp33_ASAP7_75t_R g514 ( .A(n_438), .B(n_320), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_410), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_436), .B(n_377), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_419), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_419), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_415), .Y(n_519) );
AO31x2_ASAP7_75t_L g520 ( .A1(n_440), .A2(n_403), .A3(n_380), .B(n_383), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_410), .B(n_311), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_410), .B(n_383), .Y(n_522) );
OR2x6_ASAP7_75t_L g523 ( .A(n_427), .B(n_336), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_440), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_410), .B(n_383), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_444), .B(n_383), .Y(n_526) );
NAND2xp33_ASAP7_75t_R g527 ( .A(n_450), .B(n_37), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_444), .B(n_336), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_415), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_408), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_444), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_427), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_500), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_516), .B(n_444), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_473), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_497), .B(n_444), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_497), .B(n_502), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_453), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_459), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_468), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_485), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_500), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_505), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_486), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_497), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_480), .B(n_408), .Y(n_546) );
OAI21x1_ASAP7_75t_L g547 ( .A1(n_524), .A2(n_450), .B(n_315), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_532), .B(n_38), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_491), .B(n_315), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_488), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_458), .B(n_39), .Y(n_551) );
INVx4_ASAP7_75t_L g552 ( .A(n_504), .Y(n_552) );
BUFx2_ASAP7_75t_SL g553 ( .A(n_466), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_493), .B(n_315), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_465), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_458), .B(n_42), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_462), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_477), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_467), .B(n_44), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_505), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_467), .B(n_46), .Y(n_561) );
OAI321xp33_ASAP7_75t_L g562 ( .A1(n_457), .A2(n_336), .A3(n_50), .B1(n_51), .B2(n_52), .C(n_53), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_496), .A2(n_295), .B(n_315), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_470), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_503), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_503), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_470), .B(n_49), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_495), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_494), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_475), .B(n_54), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_475), .B(n_56), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_454), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_525), .B(n_58), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_498), .B(n_61), .Y(n_574) );
AND2x4_ASAP7_75t_SL g575 ( .A(n_466), .B(n_336), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_487), .B(n_62), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_478), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_484), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_492), .B(n_63), .Y(n_579) );
OA21x2_ASAP7_75t_L g580 ( .A1(n_506), .A2(n_70), .B(n_73), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_463), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_464), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_461), .B(n_320), .Y(n_583) );
AND2x4_ASAP7_75t_SL g584 ( .A(n_482), .B(n_320), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_524), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_476), .B(n_74), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_501), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_476), .B(n_75), .Y(n_588) );
AO21x2_ASAP7_75t_L g589 ( .A1(n_474), .A2(n_76), .B(n_77), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_513), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_472), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_518), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_472), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_472), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_501), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_512), .B(n_79), .Y(n_596) );
BUFx2_ASAP7_75t_L g597 ( .A(n_507), .Y(n_597) );
NOR2xp33_ASAP7_75t_SL g598 ( .A(n_455), .B(n_81), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_509), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_489), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_472), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_507), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_512), .B(n_82), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_499), .B(n_84), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_517), .B(n_86), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_489), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_522), .B(n_87), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_515), .B(n_92), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_529), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_530), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_482), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_531), .B(n_93), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_519), .Y(n_613) );
OAI33xp33_ASAP7_75t_L g614 ( .A1(n_483), .A2(n_94), .A3(n_97), .B1(n_98), .B2(n_102), .B3(n_104), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_519), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_520), .B(n_105), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_526), .Y(n_617) );
NOR2x1_ASAP7_75t_L g618 ( .A(n_510), .B(n_106), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_520), .B(n_108), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_520), .B(n_457), .Y(n_620) );
AND2x4_ASAP7_75t_L g621 ( .A(n_494), .B(n_530), .Y(n_621) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_494), .Y(n_622) );
OA21x2_ASAP7_75t_L g623 ( .A1(n_528), .A2(n_490), .B(n_511), .Y(n_623) );
BUFx3_ASAP7_75t_L g624 ( .A(n_521), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_471), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_494), .Y(n_626) );
BUFx5_ASAP7_75t_L g627 ( .A(n_514), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_520), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_481), .A2(n_527), .B1(n_460), .B2(n_469), .Y(n_629) );
INVx2_ASAP7_75t_SL g630 ( .A(n_471), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_490), .B(n_523), .Y(n_631) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_481), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_523), .B(n_508), .Y(n_633) );
NOR2x1_ASAP7_75t_SL g634 ( .A(n_523), .B(n_456), .Y(n_634) );
INVx3_ASAP7_75t_L g635 ( .A(n_527), .Y(n_635) );
AO31x2_ASAP7_75t_L g636 ( .A1(n_490), .A2(n_511), .A3(n_514), .B(n_456), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_490), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_479), .A2(n_461), .B1(n_496), .B2(n_504), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_572), .B(n_479), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_544), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_557), .B(n_534), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_538), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_597), .Y(n_643) );
INVx3_ASAP7_75t_L g644 ( .A(n_552), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_572), .B(n_535), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_534), .B(n_565), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_578), .B(n_581), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_539), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_582), .B(n_568), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_535), .B(n_541), .Y(n_650) );
AND2x2_ASAP7_75t_SL g651 ( .A(n_552), .B(n_597), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_577), .B(n_540), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_537), .B(n_552), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_566), .B(n_638), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_541), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_537), .B(n_550), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_553), .B(n_583), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_592), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_632), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_564), .Y(n_660) );
NAND2xp67_ASAP7_75t_L g661 ( .A(n_575), .B(n_586), .Y(n_661) );
AND2x4_ASAP7_75t_SL g662 ( .A(n_630), .B(n_587), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_617), .B(n_555), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_564), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_590), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_537), .B(n_599), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_558), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_609), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_631), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_624), .B(n_602), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_600), .B(n_606), .Y(n_671) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_533), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_545), .B(n_602), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_533), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_634), .B(n_545), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_542), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_542), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_620), .B(n_591), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_543), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_543), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_624), .B(n_573), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_573), .B(n_545), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_634), .B(n_636), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_560), .Y(n_684) );
AND2x2_ASAP7_75t_SL g685 ( .A(n_629), .B(n_575), .Y(n_685) );
BUFx2_ASAP7_75t_L g686 ( .A(n_627), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_636), .B(n_595), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_620), .B(n_601), .Y(n_688) );
AND2x4_ASAP7_75t_L g689 ( .A(n_636), .B(n_595), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_560), .Y(n_690) );
NOR2x1_ASAP7_75t_L g691 ( .A(n_553), .B(n_618), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_591), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_536), .B(n_625), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_593), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_593), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_594), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_546), .B(n_630), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_546), .B(n_636), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_594), .Y(n_699) );
BUFx2_ASAP7_75t_SL g700 ( .A(n_627), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_601), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_631), .B(n_635), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_536), .B(n_613), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_636), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_536), .B(n_607), .Y(n_705) );
INVx3_ASAP7_75t_L g706 ( .A(n_627), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_611), .B(n_615), .Y(n_707) );
AND2x4_ASAP7_75t_SL g708 ( .A(n_548), .B(n_635), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_627), .B(n_635), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_627), .B(n_588), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_627), .B(n_588), .Y(n_711) );
AND2x4_ASAP7_75t_SL g712 ( .A(n_548), .B(n_627), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_637), .B(n_619), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_637), .B(n_619), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_585), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_586), .B(n_623), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_616), .B(n_585), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_616), .B(n_628), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_610), .Y(n_719) );
AND2x4_ASAP7_75t_L g720 ( .A(n_633), .B(n_621), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_614), .B(n_598), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_607), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_610), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_626), .Y(n_724) );
INVxp67_ASAP7_75t_SL g725 ( .A(n_628), .Y(n_725) );
INVx5_ASAP7_75t_L g726 ( .A(n_622), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_551), .Y(n_727) );
INVx2_ASAP7_75t_SL g728 ( .A(n_584), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_623), .B(n_604), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_551), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_623), .B(n_604), .Y(n_731) );
BUFx2_ASAP7_75t_L g732 ( .A(n_548), .Y(n_732) );
NOR3xp33_ASAP7_75t_SL g733 ( .A(n_563), .B(n_562), .C(n_554), .Y(n_733) );
AND2x4_ASAP7_75t_L g734 ( .A(n_633), .B(n_621), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_556), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_556), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_559), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_596), .B(n_603), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_559), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_626), .B(n_574), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_561), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_561), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_596), .B(n_603), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_621), .B(n_574), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_569), .B(n_549), .Y(n_745) );
BUFx2_ASAP7_75t_L g746 ( .A(n_651), .Y(n_746) );
INVx3_ASAP7_75t_L g747 ( .A(n_683), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_645), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_694), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_645), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_646), .B(n_729), .Y(n_751) );
AND2x4_ASAP7_75t_L g752 ( .A(n_683), .B(n_569), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_716), .B(n_569), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_640), .Y(n_754) );
OR2x2_ASAP7_75t_L g755 ( .A(n_678), .B(n_622), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_669), .B(n_547), .Y(n_756) );
BUFx2_ASAP7_75t_L g757 ( .A(n_644), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_695), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_654), .A2(n_605), .B1(n_576), .B2(n_579), .C(n_571), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_642), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_672), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_669), .B(n_547), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_639), .B(n_584), .Y(n_763) );
INVxp67_ASAP7_75t_L g764 ( .A(n_654), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_641), .B(n_622), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_648), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_697), .B(n_622), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_699), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_678), .B(n_622), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_663), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_663), .Y(n_771) );
OAI21x1_ASAP7_75t_L g772 ( .A1(n_704), .A2(n_580), .B(n_570), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_649), .B(n_567), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_647), .B(n_567), .Y(n_774) );
INVxp67_ASAP7_75t_L g775 ( .A(n_639), .Y(n_775) );
INVx2_ASAP7_75t_SL g776 ( .A(n_662), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g777 ( .A(n_685), .B(n_570), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_672), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_656), .B(n_652), .Y(n_779) );
AND2x4_ASAP7_75t_SL g780 ( .A(n_675), .B(n_571), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_668), .B(n_576), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_688), .B(n_589), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_688), .B(n_589), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_698), .B(n_589), .Y(n_784) );
INVx2_ASAP7_75t_SL g785 ( .A(n_675), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_702), .B(n_580), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_702), .B(n_580), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_666), .B(n_579), .Y(n_788) );
INVx2_ASAP7_75t_SL g789 ( .A(n_670), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_720), .B(n_608), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_720), .B(n_608), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_734), .B(n_612), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_650), .Y(n_793) );
NAND2x1p5_ASAP7_75t_L g794 ( .A(n_691), .B(n_612), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_667), .B(n_665), .Y(n_795) );
NAND2x1p5_ASAP7_75t_SL g796 ( .A(n_728), .B(n_709), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_734), .B(n_693), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_650), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_658), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_653), .B(n_657), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_671), .B(n_655), .Y(n_801) );
INVxp67_ASAP7_75t_L g802 ( .A(n_644), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_659), .B(n_671), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_722), .B(n_714), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_696), .Y(n_805) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_659), .Y(n_806) );
OR2x2_ASAP7_75t_L g807 ( .A(n_643), .B(n_717), .Y(n_807) );
NAND2xp5_ASAP7_75t_SL g808 ( .A(n_706), .B(n_689), .Y(n_808) );
INVx1_ASAP7_75t_SL g809 ( .A(n_681), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_687), .B(n_689), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_721), .A2(n_738), .B1(n_743), .B2(n_710), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_674), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_687), .B(n_731), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_731), .B(n_704), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_703), .B(n_714), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_701), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_713), .B(n_707), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_713), .B(n_643), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_721), .A2(n_738), .B1(n_743), .B2(n_711), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_661), .B(n_706), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_676), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_677), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_717), .B(n_684), .Y(n_823) );
BUFx2_ASAP7_75t_SL g824 ( .A(n_686), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_718), .B(n_682), .Y(n_825) );
INVx1_ASAP7_75t_SL g826 ( .A(n_712), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_718), .B(n_740), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_770), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_777), .A2(n_732), .B1(n_700), .B2(n_708), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_761), .Y(n_830) );
BUFx2_ASAP7_75t_L g831 ( .A(n_796), .Y(n_831) );
INVx2_ASAP7_75t_SL g832 ( .A(n_776), .Y(n_832) );
AOI22xp33_ASAP7_75t_SL g833 ( .A1(n_746), .A2(n_673), .B1(n_744), .B2(n_705), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_771), .Y(n_834) );
OR2x2_ASAP7_75t_L g835 ( .A(n_796), .B(n_679), .Y(n_835) );
OAI322xp33_ASAP7_75t_L g836 ( .A1(n_764), .A2(n_745), .A3(n_727), .B1(n_730), .B2(n_735), .C1(n_736), .C2(n_742), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_793), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_777), .A2(n_733), .B1(n_744), .B2(n_726), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_798), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_818), .B(n_660), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_801), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_748), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_810), .B(n_692), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_811), .B(n_692), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_750), .Y(n_845) );
OAI211xp5_ASAP7_75t_L g846 ( .A1(n_819), .A2(n_733), .B(n_739), .C(n_737), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_795), .Y(n_847) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_806), .Y(n_848) );
OR2x6_ASAP7_75t_L g849 ( .A(n_776), .B(n_715), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_810), .B(n_741), .Y(n_850) );
OAI33xp33_ASAP7_75t_L g851 ( .A1(n_775), .A2(n_664), .A3(n_680), .B1(n_690), .B2(n_724), .B3(n_723), .Y(n_851) );
AND2x4_ASAP7_75t_L g852 ( .A(n_747), .B(n_725), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_778), .Y(n_853) );
AND2x4_ASAP7_75t_L g854 ( .A(n_747), .B(n_725), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_815), .B(n_719), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_803), .Y(n_856) );
OR2x2_ASAP7_75t_L g857 ( .A(n_804), .B(n_726), .Y(n_857) );
OR2x2_ASAP7_75t_L g858 ( .A(n_817), .B(n_726), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_803), .Y(n_859) );
AND2x2_ASAP7_75t_L g860 ( .A(n_751), .B(n_726), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_751), .B(n_813), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_813), .B(n_797), .Y(n_862) );
INVxp67_ASAP7_75t_L g863 ( .A(n_757), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_754), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_760), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_815), .B(n_827), .Y(n_866) );
AND2x4_ASAP7_75t_L g867 ( .A(n_747), .B(n_785), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_766), .Y(n_868) );
INVxp67_ASAP7_75t_SL g869 ( .A(n_778), .Y(n_869) );
AND2x4_ASAP7_75t_L g870 ( .A(n_785), .B(n_752), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_799), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_759), .A2(n_780), .B1(n_763), .B2(n_784), .Y(n_872) );
NAND4xp75_ASAP7_75t_L g873 ( .A(n_820), .B(n_808), .C(n_784), .D(n_787), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_827), .B(n_814), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_800), .B(n_779), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g876 ( .A1(n_780), .A2(n_794), .B1(n_787), .B2(n_786), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_831), .A2(n_789), .B1(n_826), .B2(n_808), .Y(n_877) );
OAI21xp33_ASAP7_75t_SL g878 ( .A1(n_873), .A2(n_789), .B(n_797), .Y(n_878) );
A2O1A1Ixp33_ASAP7_75t_L g879 ( .A1(n_832), .A2(n_752), .B(n_814), .C(n_802), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_856), .Y(n_880) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_848), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_872), .A2(n_753), .B1(n_786), .B2(n_762), .Y(n_882) );
NAND4xp75_ASAP7_75t_L g883 ( .A(n_872), .B(n_783), .C(n_782), .D(n_762), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_846), .A2(n_753), .B1(n_756), .B2(n_769), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_859), .Y(n_885) );
INVx1_ASAP7_75t_SL g886 ( .A(n_849), .Y(n_886) );
OAI21xp5_ASAP7_75t_L g887 ( .A1(n_838), .A2(n_794), .B(n_772), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_837), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_839), .Y(n_889) );
OAI21xp5_ASAP7_75t_L g890 ( .A1(n_849), .A2(n_772), .B(n_752), .Y(n_890) );
OAI31xp33_ASAP7_75t_L g891 ( .A1(n_867), .A2(n_809), .A3(n_756), .B(n_782), .Y(n_891) );
OAI21xp33_ASAP7_75t_L g892 ( .A1(n_833), .A2(n_783), .B(n_825), .Y(n_892) );
XOR2x2_ASAP7_75t_L g893 ( .A(n_875), .B(n_825), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_842), .Y(n_894) );
INVx1_ASAP7_75t_SL g895 ( .A(n_867), .Y(n_895) );
AOI21xp33_ASAP7_75t_L g896 ( .A1(n_844), .A2(n_781), .B(n_755), .Y(n_896) );
OAI21xp33_ASAP7_75t_SL g897 ( .A1(n_876), .A2(n_790), .B(n_792), .Y(n_897) );
NAND3xp33_ASAP7_75t_L g898 ( .A(n_863), .B(n_812), .C(n_822), .Y(n_898) );
OAI21xp5_ASAP7_75t_L g899 ( .A1(n_835), .A2(n_807), .B(n_773), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_852), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_876), .A2(n_829), .B1(n_870), .B2(n_866), .Y(n_901) );
OAI221xp5_ASAP7_75t_L g902 ( .A1(n_829), .A2(n_824), .B1(n_823), .B2(n_755), .C(n_774), .Y(n_902) );
OR4x1_ASAP7_75t_L g903 ( .A(n_841), .B(n_821), .C(n_767), .D(n_769), .Y(n_903) );
OR2x2_ASAP7_75t_L g904 ( .A(n_881), .B(n_840), .Y(n_904) );
NAND2xp5_ASAP7_75t_SL g905 ( .A(n_878), .B(n_870), .Y(n_905) );
OAI221xp5_ASAP7_75t_L g906 ( .A1(n_887), .A2(n_847), .B1(n_858), .B2(n_857), .C(n_828), .Y(n_906) );
OAI31xp33_ASAP7_75t_L g907 ( .A1(n_901), .A2(n_854), .A3(n_852), .B(n_860), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_880), .B(n_834), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_888), .Y(n_909) );
OAI22xp33_ASAP7_75t_SL g910 ( .A1(n_877), .A2(n_854), .B1(n_871), .B2(n_865), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_903), .Y(n_911) );
OR2x2_ASAP7_75t_L g912 ( .A(n_885), .B(n_874), .Y(n_912) );
OR2x2_ASAP7_75t_L g913 ( .A(n_886), .B(n_830), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_889), .Y(n_914) );
AOI221xp5_ASAP7_75t_L g915 ( .A1(n_892), .A2(n_851), .B1(n_836), .B2(n_864), .C(n_868), .Y(n_915) );
AOI22xp5_ASAP7_75t_L g916 ( .A1(n_893), .A2(n_861), .B1(n_845), .B2(n_843), .Y(n_916) );
OAI21xp33_ASAP7_75t_SL g917 ( .A1(n_890), .A2(n_862), .B(n_869), .Y(n_917) );
A2O1A1Ixp33_ASAP7_75t_L g918 ( .A1(n_897), .A2(n_850), .B(n_855), .C(n_792), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_915), .B(n_894), .Y(n_919) );
NAND3xp33_ASAP7_75t_L g920 ( .A(n_907), .B(n_887), .C(n_890), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_911), .B(n_895), .Y(n_921) );
NAND3xp33_ASAP7_75t_SL g922 ( .A(n_905), .B(n_891), .C(n_879), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_916), .B(n_882), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_913), .B(n_900), .Y(n_924) );
NAND3xp33_ASAP7_75t_L g925 ( .A(n_917), .B(n_884), .C(n_898), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_904), .Y(n_926) );
AOI21xp5_ASAP7_75t_L g927 ( .A1(n_919), .A2(n_910), .B(n_906), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_926), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_924), .B(n_916), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g930 ( .A1(n_922), .A2(n_883), .B1(n_902), .B2(n_914), .Y(n_930) );
AOI222xp33_ASAP7_75t_L g931 ( .A1(n_928), .A2(n_920), .B1(n_925), .B2(n_923), .C1(n_909), .C2(n_899), .Y(n_931) );
AOI21xp5_ASAP7_75t_L g932 ( .A1(n_927), .A2(n_921), .B(n_918), .Y(n_932) );
OAI21xp5_ASAP7_75t_SL g933 ( .A1(n_930), .A2(n_899), .B(n_896), .Y(n_933) );
INVx1_ASAP7_75t_SL g934 ( .A(n_932), .Y(n_934) );
INVx2_ASAP7_75t_L g935 ( .A(n_933), .Y(n_935) );
NOR3xp33_ASAP7_75t_L g936 ( .A(n_934), .B(n_929), .C(n_931), .Y(n_936) );
INVx3_ASAP7_75t_SL g937 ( .A(n_935), .Y(n_937) );
BUFx2_ASAP7_75t_L g938 ( .A(n_937), .Y(n_938) );
OR2x2_ASAP7_75t_L g939 ( .A(n_936), .B(n_912), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_938), .A2(n_908), .B1(n_853), .B2(n_765), .Y(n_940) );
XOR2xp5_ASAP7_75t_L g941 ( .A(n_939), .B(n_765), .Y(n_941) );
HB1xp67_ASAP7_75t_L g942 ( .A(n_941), .Y(n_942) );
AO22x2_ASAP7_75t_L g943 ( .A1(n_942), .A2(n_940), .B1(n_791), .B2(n_790), .Y(n_943) );
XNOR2xp5_ASAP7_75t_L g944 ( .A(n_943), .B(n_791), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_944), .A2(n_836), .B1(n_788), .B2(n_805), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_945), .A2(n_788), .B1(n_805), .B2(n_816), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_946), .B(n_816), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_947), .A2(n_768), .B1(n_749), .B2(n_758), .Y(n_948) );
endmodule