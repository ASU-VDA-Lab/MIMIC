module fake_aes_5536_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
OA21x2_ASAP7_75t_L g12 ( .A1(n_3), .A2(n_2), .B(n_8), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
BUFx3_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_14), .B(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_14), .B(n_0), .Y(n_17) );
AND2x6_ASAP7_75t_SL g18 ( .A(n_11), .B(n_1), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_12), .B(n_13), .Y(n_20) );
BUFx3_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
BUFx2_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
AOI221xp5_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_19), .B1(n_13), .B2(n_11), .C(n_15), .Y(n_24) );
XNOR2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_12), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_23), .B(n_21), .Y(n_26) );
OAI22xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_21), .B1(n_12), .B2(n_18), .Y(n_27) );
OAI21xp5_ASAP7_75t_SL g28 ( .A1(n_25), .A2(n_11), .B(n_4), .Y(n_28) );
OR5x1_ASAP7_75t_L g29 ( .A(n_28), .B(n_2), .C(n_5), .D(n_11), .E(n_15), .Y(n_29) );
AOI21xp5_ASAP7_75t_SL g30 ( .A1(n_27), .A2(n_26), .B(n_21), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
AOI222xp33_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_11), .B1(n_5), .B2(n_21), .C1(n_10), .C2(n_6), .Y(n_33) );
OA21x2_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_31), .B(n_9), .Y(n_34) );
endmodule