module fake_jpeg_30810_n_28 (n_3, n_2, n_1, n_0, n_4, n_5, n_28);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_28;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx16f_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_2),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_3),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_7),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_9),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_0),
.B1(n_4),
.B2(n_2),
.Y(n_14)
);

AOI22x1_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_15),
.B1(n_6),
.B2(n_7),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g15 ( 
.A1(n_11),
.A2(n_1),
.B1(n_3),
.B2(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_17),
.B(n_8),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_18),
.A2(n_6),
.B1(n_12),
.B2(n_10),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_21),
.B1(n_10),
.B2(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_20),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_23),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_23),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_24),
.Y(n_28)
);


endmodule