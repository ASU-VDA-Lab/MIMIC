module fake_aes_9658_n_616 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_616);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_616;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_599;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g72 ( .A(n_62), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_59), .Y(n_73) );
INVx2_ASAP7_75t_L g74 ( .A(n_49), .Y(n_74) );
INVx2_ASAP7_75t_L g75 ( .A(n_50), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_25), .Y(n_76) );
CKINVDCx16_ASAP7_75t_R g77 ( .A(n_60), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_31), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_45), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_36), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_0), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_12), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_67), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_4), .Y(n_84) );
BUFx2_ASAP7_75t_L g85 ( .A(n_69), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_13), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_23), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_8), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_57), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_70), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_1), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_0), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_65), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_58), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_24), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_33), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_47), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_21), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_29), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_63), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_22), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_4), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_37), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_10), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_44), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_11), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_10), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_2), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_52), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_16), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_66), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_13), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_28), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_8), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_85), .B(n_1), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
INVx3_ASAP7_75t_L g118 ( .A(n_104), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_85), .B(n_2), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_73), .Y(n_120) );
AND2x4_ASAP7_75t_L g121 ( .A(n_109), .B(n_3), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_104), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_78), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_87), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_74), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_109), .B(n_3), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_91), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_77), .B(n_5), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_84), .B(n_5), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_79), .Y(n_133) );
INVx1_ASAP7_75t_SL g134 ( .A(n_91), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_87), .B(n_6), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_105), .B(n_6), .Y(n_137) );
INVx1_ASAP7_75t_SL g138 ( .A(n_107), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_80), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_92), .B(n_7), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_80), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_87), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_87), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_74), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_90), .Y(n_146) );
CKINVDCx16_ASAP7_75t_R g147 ( .A(n_72), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_94), .Y(n_148) );
NOR2x1_ASAP7_75t_L g149 ( .A(n_95), .B(n_7), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_75), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_86), .B(n_9), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_82), .B(n_9), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g153 ( .A1(n_108), .A2(n_11), .B1(n_12), .B2(n_14), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_86), .B(n_15), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_151), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_151), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_148), .B(n_75), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_121), .Y(n_158) );
INVx2_ASAP7_75t_SL g159 ( .A(n_130), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_117), .B(n_76), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_121), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_117), .B(n_96), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_120), .B(n_76), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_151), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_122), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_147), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_120), .B(n_96), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_154), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_124), .B(n_103), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_124), .B(n_103), .Y(n_172) );
OR2x2_ASAP7_75t_L g173 ( .A(n_136), .B(n_81), .Y(n_173) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_134), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_154), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_147), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_138), .B(n_102), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_131), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_122), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_122), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
NOR2xp33_ASAP7_75t_SL g182 ( .A(n_131), .B(n_98), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_122), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_148), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_137), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_126), .B(n_101), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_121), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_148), .Y(n_188) );
AND2x6_ASAP7_75t_L g189 ( .A(n_119), .B(n_113), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_122), .Y(n_190) );
OR2x6_ASAP7_75t_L g191 ( .A(n_153), .B(n_102), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_126), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_127), .Y(n_193) );
INVx6_ASAP7_75t_L g194 ( .A(n_119), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_127), .B(n_101), .Y(n_195) );
AO22x2_ASAP7_75t_L g196 ( .A1(n_137), .A2(n_106), .B1(n_112), .B2(n_88), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_133), .B(n_89), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_133), .B(n_89), .Y(n_198) );
INVx4_ASAP7_75t_SL g199 ( .A(n_139), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_139), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_128), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_125), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_164), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_174), .B(n_129), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g205 ( .A1(n_156), .A2(n_141), .B(n_146), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_192), .B(n_143), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_164), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_178), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_177), .B(n_152), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_194), .B(n_116), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_158), .B(n_132), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_158), .B(n_140), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_170), .A2(n_143), .B(n_146), .C(n_141), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_201), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_189), .A2(n_153), .B1(n_149), .B2(n_135), .Y(n_215) );
OR2x2_ASAP7_75t_L g216 ( .A(n_173), .B(n_118), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_162), .A2(n_150), .B(n_128), .C(n_145), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_178), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_189), .A2(n_149), .B1(n_112), .B2(n_106), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_201), .Y(n_220) );
INVx2_ASAP7_75t_SL g221 ( .A(n_194), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_158), .B(n_100), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_189), .A2(n_115), .B1(n_93), .B2(n_145), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_159), .B(n_118), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_194), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_185), .Y(n_227) );
INVx1_ASAP7_75t_SL g228 ( .A(n_189), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_163), .B(n_123), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_193), .B(n_150), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_184), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_169), .B(n_123), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_175), .B(n_118), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_188), .Y(n_234) );
NAND2xp33_ASAP7_75t_L g235 ( .A(n_189), .B(n_111), .Y(n_235) );
OR2x6_ASAP7_75t_L g236 ( .A(n_196), .B(n_123), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_187), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_161), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_171), .B(n_123), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_161), .B(n_97), .Y(n_240) );
BUFx12f_ASAP7_75t_L g241 ( .A(n_168), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_187), .B(n_99), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_185), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_161), .B(n_113), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_172), .B(n_111), .Y(n_245) );
INVx5_ASAP7_75t_L g246 ( .A(n_155), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_166), .B(n_110), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_199), .B(n_110), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_200), .B(n_94), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_155), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_182), .A2(n_114), .B1(n_83), .B2(n_125), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_168), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_195), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_198), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_176), .B(n_197), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_199), .B(n_114), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_250), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_206), .Y(n_258) );
NOR2xp33_ASAP7_75t_R g259 ( .A(n_241), .B(n_186), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_243), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_238), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_213), .A2(n_197), .B(n_165), .C(n_160), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_238), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_253), .B(n_199), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_204), .A2(n_196), .B1(n_191), .B2(n_165), .Y(n_265) );
AO22x1_ASAP7_75t_L g266 ( .A1(n_252), .A2(n_191), .B1(n_196), .B2(n_186), .Y(n_266) );
OAI22xp5_ASAP7_75t_SL g267 ( .A1(n_236), .A2(n_191), .B1(n_160), .B2(n_83), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_206), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_238), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_203), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_228), .B(n_157), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_236), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_203), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_205), .A2(n_157), .B(n_142), .C(n_144), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_236), .B(n_144), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_254), .B(n_144), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_205), .B(n_144), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_226), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_219), .A2(n_125), .B1(n_142), .B2(n_144), .Y(n_279) );
AOI22xp33_ASAP7_75t_SL g280 ( .A1(n_235), .A2(n_125), .B1(n_142), .B2(n_202), .Y(n_280) );
INVx5_ASAP7_75t_L g281 ( .A(n_203), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_231), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_207), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_228), .B(n_125), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_234), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_210), .B(n_17), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_207), .B(n_142), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_208), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_218), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_227), .Y(n_290) );
AO22x1_ASAP7_75t_L g291 ( .A1(n_255), .A2(n_142), .B1(n_19), .B2(n_20), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_245), .B(n_209), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_207), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_246), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_244), .A2(n_190), .B(n_183), .C(n_180), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g296 ( .A1(n_217), .A2(n_190), .B(n_183), .C(n_180), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_209), .B(n_18), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_246), .Y(n_298) );
OA21x2_ASAP7_75t_L g299 ( .A1(n_249), .A2(n_179), .B(n_167), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_215), .A2(n_179), .B1(n_167), .B2(n_202), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_223), .Y(n_301) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_296), .A2(n_256), .B(n_230), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_258), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_260), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_268), .B(n_232), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_292), .B(n_216), .Y(n_306) );
INVx6_ASAP7_75t_L g307 ( .A(n_281), .Y(n_307) );
OA21x2_ASAP7_75t_L g308 ( .A1(n_274), .A2(n_230), .B(n_229), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_278), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_301), .A2(n_225), .B1(n_221), .B2(n_224), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_281), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_289), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_292), .B(n_239), .Y(n_313) );
OA21x2_ASAP7_75t_L g314 ( .A1(n_277), .A2(n_295), .B(n_276), .Y(n_314) );
AOI22xp33_ASAP7_75t_SL g315 ( .A1(n_267), .A2(n_242), .B1(n_233), .B2(n_246), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_272), .B(n_246), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_296), .A2(n_248), .B(n_251), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_265), .A2(n_220), .B1(n_214), .B2(n_247), .Y(n_319) );
OA21x2_ASAP7_75t_L g320 ( .A1(n_277), .A2(n_240), .B(n_222), .Y(n_320) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_276), .A2(n_212), .B(n_211), .Y(n_321) );
INVxp67_ASAP7_75t_L g322 ( .A(n_290), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_263), .Y(n_323) );
OAI21x1_ASAP7_75t_L g324 ( .A1(n_299), .A2(n_26), .B(n_27), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_285), .B(n_237), .Y(n_325) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_281), .B(n_202), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_281), .Y(n_327) );
AOI22xp33_ASAP7_75t_SL g328 ( .A1(n_288), .A2(n_202), .B1(n_32), .B2(n_34), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_257), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_266), .A2(n_30), .B1(n_35), .B2(n_38), .C(n_39), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_315), .A2(n_286), .B1(n_297), .B2(n_259), .Y(n_331) );
OAI211xp5_ASAP7_75t_L g332 ( .A1(n_310), .A2(n_262), .B(n_300), .C(n_280), .Y(n_332) );
AOI222xp33_ASAP7_75t_L g333 ( .A1(n_306), .A2(n_286), .B1(n_279), .B2(n_275), .C1(n_271), .C2(n_298), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_312), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_309), .Y(n_336) );
AOI222xp33_ASAP7_75t_L g337 ( .A1(n_306), .A2(n_279), .B1(n_283), .B2(n_294), .C1(n_291), .C2(n_264), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_304), .B(n_294), .Y(n_338) );
OA21x2_ASAP7_75t_L g339 ( .A1(n_324), .A2(n_287), .B(n_284), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_303), .B(n_264), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_319), .A2(n_261), .B1(n_263), .B2(n_269), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_313), .B(n_262), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_313), .B(n_263), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_303), .B(n_269), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_309), .Y(n_345) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_304), .A2(n_319), .B1(n_317), .B2(n_305), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_307), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_317), .A2(n_283), .B1(n_280), .B2(n_269), .C(n_270), .Y(n_348) );
OAI321xp33_ASAP7_75t_L g349 ( .A1(n_330), .A2(n_293), .A3(n_273), .B1(n_42), .B2(n_43), .C(n_46), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_322), .A2(n_270), .B1(n_299), .B2(n_273), .C(n_293), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_329), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_305), .B(n_273), .Y(n_352) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_329), .A2(n_293), .B1(n_41), .B2(n_48), .C1(n_51), .C2(n_53), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_307), .A2(n_325), .B1(n_311), .B2(n_327), .Y(n_354) );
OAI22xp33_ASAP7_75t_L g355 ( .A1(n_330), .A2(n_40), .B1(n_54), .B2(n_55), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_335), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_345), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_345), .B(n_327), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_343), .B(n_311), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_343), .B(n_323), .Y(n_360) );
INVx2_ASAP7_75t_R g361 ( .A(n_336), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_352), .Y(n_362) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_352), .Y(n_363) );
OAI221xp5_ASAP7_75t_L g364 ( .A1(n_331), .A2(n_328), .B1(n_325), .B2(n_308), .C(n_314), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_340), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_351), .B(n_323), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_346), .A2(n_316), .B1(n_323), .B2(n_326), .C(n_308), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_340), .B(n_323), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_342), .B(n_314), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_334), .B(n_314), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_340), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_344), .Y(n_372) );
BUFx2_ASAP7_75t_L g373 ( .A(n_335), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_344), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_339), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_339), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_347), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_350), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_338), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_347), .B(n_314), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_347), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_341), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_348), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_354), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_333), .B(n_308), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_369), .B(n_308), .Y(n_387) );
BUFx12f_ASAP7_75t_L g388 ( .A(n_373), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_357), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_358), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_373), .Y(n_391) );
AOI21xp5_ASAP7_75t_SL g392 ( .A1(n_367), .A2(n_355), .B(n_349), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_357), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_376), .Y(n_394) );
AO21x2_ASAP7_75t_L g395 ( .A1(n_379), .A2(n_324), .B(n_332), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_369), .B(n_321), .Y(n_396) );
INVx4_ASAP7_75t_L g397 ( .A(n_365), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_381), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_381), .B(n_302), .Y(n_399) );
INVxp33_ASAP7_75t_L g400 ( .A(n_356), .Y(n_400) );
OR2x6_ASAP7_75t_L g401 ( .A(n_386), .B(n_307), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_358), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_386), .B(n_321), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_370), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_376), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_370), .B(n_302), .Y(n_406) );
INVx4_ASAP7_75t_L g407 ( .A(n_365), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_380), .B(n_321), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_361), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_380), .B(n_362), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_361), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_380), .B(n_337), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_385), .A2(n_307), .B1(n_316), .B2(n_320), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_361), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_376), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_362), .B(n_321), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_374), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_363), .B(n_320), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_374), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_372), .B(n_320), .Y(n_420) );
OAI33xp33_ASAP7_75t_L g421 ( .A1(n_372), .A2(n_353), .A3(n_61), .B1(n_64), .B2(n_68), .B3(n_56), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_360), .B(n_320), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_375), .B(n_326), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_359), .B(n_316), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_360), .B(n_318), .Y(n_425) );
OR2x2_ASAP7_75t_SL g426 ( .A(n_385), .B(n_326), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_377), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_359), .B(n_318), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_365), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_385), .B(n_316), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_403), .B(n_375), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_394), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_393), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_393), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_390), .B(n_402), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_398), .B(n_379), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_394), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_403), .B(n_377), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
OAI21xp5_ASAP7_75t_SL g440 ( .A1(n_391), .A2(n_384), .B(n_364), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_388), .Y(n_441) );
NOR2x1_ASAP7_75t_L g442 ( .A(n_397), .B(n_378), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_398), .B(n_383), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_387), .B(n_377), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_404), .B(n_383), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_389), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_417), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_402), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_387), .B(n_377), .Y(n_449) );
INVxp67_ASAP7_75t_SL g450 ( .A(n_418), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_388), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_396), .B(n_377), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_417), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_429), .B(n_384), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_396), .B(n_377), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_405), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_419), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_405), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_404), .B(n_371), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_415), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_415), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_422), .B(n_425), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_422), .B(n_366), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_429), .B(n_371), .Y(n_465) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_418), .Y(n_466) );
NAND2xp33_ASAP7_75t_L g467 ( .A(n_400), .B(n_366), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_424), .B(n_371), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_425), .B(n_382), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_420), .Y(n_470) );
AOI22x1_ASAP7_75t_L g471 ( .A1(n_397), .A2(n_368), .B1(n_382), .B2(n_378), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_428), .B(n_378), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_420), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_408), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_408), .Y(n_475) );
OAI222xp33_ASAP7_75t_L g476 ( .A1(n_401), .A2(n_368), .B1(n_397), .B2(n_407), .C1(n_412), .C2(n_423), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_409), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_399), .B(n_368), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_410), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_428), .B(n_368), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_409), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_416), .B(n_410), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_416), .B(n_401), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_436), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_479), .B(n_401), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_463), .B(n_406), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_463), .B(n_406), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_448), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_448), .Y(n_489) );
OAI21xp33_ASAP7_75t_L g490 ( .A1(n_440), .A2(n_392), .B(n_430), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_432), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_436), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_431), .B(n_406), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_438), .B(n_406), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_433), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_431), .B(n_407), .Y(n_496) );
XNOR2x2_ASAP7_75t_L g497 ( .A(n_435), .B(n_413), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_442), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_471), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_482), .B(n_401), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_433), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_482), .B(n_401), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_434), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_434), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_451), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_464), .B(n_407), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_467), .A2(n_392), .B(n_423), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_447), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_478), .B(n_414), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_447), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_464), .B(n_407), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_438), .B(n_399), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_477), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_444), .B(n_399), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_480), .B(n_399), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_443), .B(n_426), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_453), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_454), .B(n_421), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_453), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_432), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_444), .B(n_449), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_477), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_455), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_443), .B(n_426), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_470), .B(n_395), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_449), .B(n_411), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_455), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_458), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_441), .B(n_411), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_481), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_458), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_484), .B(n_470), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_492), .B(n_473), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_521), .B(n_478), .Y(n_534) );
BUFx2_ASAP7_75t_L g535 ( .A(n_488), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_499), .A2(n_476), .B(n_471), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_495), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_501), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_529), .B(n_473), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_490), .A2(n_478), .B1(n_480), .B2(n_483), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_518), .A2(n_468), .B1(n_469), .B2(n_478), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_518), .A2(n_451), .B(n_465), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_493), .B(n_450), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_503), .Y(n_544) );
NOR2xp67_ASAP7_75t_SL g545 ( .A(n_499), .B(n_483), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_498), .B(n_481), .Y(n_546) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_497), .A2(n_466), .B1(n_472), .B2(n_452), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_529), .B(n_469), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g549 ( .A1(n_507), .A2(n_475), .B1(n_474), .B2(n_445), .C(n_472), .Y(n_549) );
OAI221xp5_ASAP7_75t_L g550 ( .A1(n_505), .A2(n_445), .B1(n_460), .B2(n_481), .C(n_474), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_500), .A2(n_460), .B1(n_475), .B2(n_456), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_504), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_508), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_491), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_498), .B(n_439), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_510), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_488), .A2(n_414), .B(n_446), .C(n_439), .Y(n_557) );
INVxp33_ASAP7_75t_L g558 ( .A(n_506), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_517), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_496), .A2(n_456), .B1(n_452), .B2(n_446), .Y(n_560) );
NOR3xp33_ASAP7_75t_SL g561 ( .A(n_497), .B(n_395), .C(n_427), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_489), .B(n_437), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_521), .B(n_437), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_519), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_536), .A2(n_489), .B(n_511), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_563), .B(n_526), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_554), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_541), .B(n_526), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_532), .Y(n_569) );
XNOR2xp5_ASAP7_75t_L g570 ( .A(n_560), .B(n_487), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_542), .A2(n_516), .B(n_524), .C(n_525), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_533), .Y(n_572) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_547), .A2(n_485), .B1(n_502), .B2(n_530), .C(n_531), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_537), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_535), .Y(n_575) );
XNOR2xp5_ASAP7_75t_L g576 ( .A(n_558), .B(n_487), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_538), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_557), .A2(n_530), .B(n_520), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_534), .B(n_486), .Y(n_579) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_561), .B(n_530), .C(n_520), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_539), .B(n_549), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_548), .B(n_486), .Y(n_582) );
A2O1A1Ixp33_ASAP7_75t_L g583 ( .A1(n_545), .A2(n_509), .B(n_515), .C(n_494), .Y(n_583) );
NOR3xp33_ASAP7_75t_L g584 ( .A(n_547), .B(n_528), .C(n_527), .Y(n_584) );
AO21x1_ASAP7_75t_L g585 ( .A1(n_584), .A2(n_557), .B(n_555), .Y(n_585) );
CKINVDCx14_ASAP7_75t_R g586 ( .A(n_576), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_574), .Y(n_587) );
XNOR2x1_ASAP7_75t_L g588 ( .A(n_565), .B(n_543), .Y(n_588) );
AOI211xp5_ASAP7_75t_L g589 ( .A1(n_573), .A2(n_550), .B(n_551), .C(n_546), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_577), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_575), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_567), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_583), .A2(n_562), .B(n_540), .Y(n_593) );
NOR3xp33_ASAP7_75t_L g594 ( .A(n_571), .B(n_564), .C(n_553), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_SL g595 ( .A1(n_571), .A2(n_544), .B(n_552), .C(n_556), .Y(n_595) );
AOI21xp33_ASAP7_75t_L g596 ( .A1(n_581), .A2(n_580), .B(n_568), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_586), .A2(n_570), .B1(n_569), .B2(n_572), .Y(n_597) );
OAI211xp5_ASAP7_75t_L g598 ( .A1(n_596), .A2(n_561), .B(n_578), .C(n_582), .Y(n_598) );
AOI222xp33_ASAP7_75t_L g599 ( .A1(n_595), .A2(n_559), .B1(n_523), .B2(n_579), .C1(n_509), .C2(n_494), .Y(n_599) );
NOR2xp67_ASAP7_75t_L g600 ( .A(n_593), .B(n_578), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_596), .A2(n_566), .B1(n_509), .B2(n_514), .C(n_512), .Y(n_601) );
CKINVDCx16_ASAP7_75t_R g602 ( .A(n_591), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_585), .A2(n_514), .B1(n_512), .B2(n_513), .Y(n_603) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_603), .B(n_594), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_600), .Y(n_605) );
NAND4xp75_ASAP7_75t_L g606 ( .A(n_597), .B(n_592), .C(n_590), .D(n_587), .Y(n_606) );
AND3x4_ASAP7_75t_L g607 ( .A(n_602), .B(n_599), .C(n_598), .Y(n_607) );
NOR3xp33_ASAP7_75t_L g608 ( .A(n_606), .B(n_601), .C(n_589), .Y(n_608) );
OR4x2_ASAP7_75t_L g609 ( .A(n_607), .B(n_588), .C(n_491), .D(n_513), .Y(n_609) );
OAI22xp5_ASAP7_75t_SL g610 ( .A1(n_609), .A2(n_604), .B1(n_605), .B2(n_522), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_608), .Y(n_611) );
AND3x4_ASAP7_75t_L g612 ( .A(n_611), .B(n_605), .C(n_522), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_612), .Y(n_613) );
AOI22xp5_ASAP7_75t_SL g614 ( .A1(n_613), .A2(n_610), .B1(n_457), .B2(n_459), .Y(n_614) );
OAI221xp5_ASAP7_75t_R g615 ( .A1(n_614), .A2(n_395), .B1(n_427), .B2(n_457), .C(n_459), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_615), .A2(n_461), .B1(n_462), .B2(n_611), .C(n_608), .Y(n_616) );
endmodule