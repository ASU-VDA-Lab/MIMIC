module fake_jpeg_29085_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_62),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_19),
.B(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_63),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_29),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_14),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_7),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_28),
.Y(n_86)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_68),
.B(n_82),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_35),
.B1(n_38),
.B2(n_37),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_72),
.A2(n_79),
.B1(n_85),
.B2(n_93),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_35),
.B1(n_38),
.B2(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_18),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_35),
.B1(n_26),
.B2(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_90),
.B(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_17),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_108),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_42),
.A2(n_35),
.B1(n_17),
.B2(n_27),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_27),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_16),
.B1(n_23),
.B2(n_22),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_100),
.B1(n_110),
.B2(n_15),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_39),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_29),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_20),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_58),
.B1(n_56),
.B2(n_51),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_20),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_45),
.B(n_16),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_23),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_109),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_49),
.B(n_22),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_43),
.B(n_21),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_18),
.B1(n_15),
.B2(n_24),
.Y(n_110)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_125),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_117),
.B(n_123),
.Y(n_193)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_29),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_121),
.B(n_124),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_50),
.C(n_48),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_136),
.C(n_148),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_29),
.B1(n_26),
.B2(n_2),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_139),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_26),
.B1(n_9),
.B2(n_11),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_68),
.B(n_0),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_0),
.B(n_1),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_149),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_9),
.C(n_12),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_74),
.A2(n_9),
.B(n_12),
.C(n_11),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_87),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_92),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_77),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_107),
.A2(n_5),
.B1(n_12),
.B2(n_13),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_145),
.A2(n_154),
.B1(n_89),
.B2(n_76),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_91),
.A2(n_13),
.B1(n_2),
.B2(n_4),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_147),
.A2(n_70),
.B1(n_111),
.B2(n_83),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_80),
.B(n_0),
.C(n_4),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_73),
.B(n_0),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_73),
.B(n_4),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_155),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_105),
.A2(n_91),
.B1(n_106),
.B2(n_78),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_151),
.A2(n_127),
.B1(n_146),
.B2(n_113),
.Y(n_189)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_105),
.A2(n_88),
.B1(n_89),
.B2(n_70),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_89),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_159),
.B(n_161),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_193),
.B1(n_165),
.B2(n_190),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_87),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_83),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_81),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_183),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_95),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_179),
.C(n_185),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_122),
.C(n_129),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_101),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_121),
.B(n_95),
.C(n_111),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_116),
.B(n_136),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_187),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_189),
.A2(n_160),
.B1(n_180),
.B2(n_166),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_133),
.B(n_134),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_114),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_150),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_121),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_200),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_190),
.A2(n_124),
.B(n_140),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_195),
.A2(n_203),
.B(n_207),
.Y(n_236)
);

AND2x4_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_124),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_196),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_124),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_132),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_211),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_178),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_202),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_SL g203 ( 
.A(n_161),
.B(n_142),
.C(n_151),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_173),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_204),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_127),
.B1(n_137),
.B2(n_120),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_225),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_193),
.A2(n_114),
.B1(n_126),
.B2(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_156),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_177),
.C(n_167),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_182),
.C(n_184),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_173),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_220),
.C(n_168),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_156),
.B(n_167),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_174),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_158),
.B(n_191),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_224),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_163),
.A2(n_165),
.B(n_170),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_169),
.B(n_182),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_178),
.B(n_166),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_189),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_198),
.B1(n_213),
.B2(n_204),
.Y(n_248)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_163),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_164),
.B(n_162),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_162),
.B1(n_164),
.B2(n_184),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_235),
.C(n_236),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_228),
.A2(n_245),
.B(n_240),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_210),
.A2(n_176),
.B1(n_174),
.B2(n_169),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_232),
.A2(n_238),
.B1(n_241),
.B2(n_248),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_234),
.B(n_205),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_237),
.B(n_208),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_168),
.B1(n_176),
.B2(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_200),
.A2(n_168),
.B1(n_217),
.B2(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

AOI221xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_195),
.B1(n_197),
.B2(n_218),
.C(n_196),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_207),
.A2(n_199),
.B(n_216),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_223),
.B1(n_198),
.B2(n_199),
.Y(n_250)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_254),
.Y(n_285)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_256),
.B(n_263),
.Y(n_283)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_261),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_214),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_259),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_246),
.Y(n_259)
);

AOI221xp5_ASAP7_75t_L g260 ( 
.A1(n_245),
.A2(n_194),
.B1(n_196),
.B2(n_223),
.C(n_212),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_250),
.Y(n_281)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_196),
.C(n_205),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_221),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_230),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_249),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_226),
.C(n_235),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_281),
.C(n_256),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_241),
.B1(n_237),
.B2(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_279),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_253),
.B(n_231),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_231),
.Y(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_262),
.A2(n_249),
.B1(n_236),
.B2(n_238),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_271),
.B(n_227),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_247),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_281),
.C(n_277),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_285),
.B(n_266),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_288),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_233),
.C(n_264),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_273),
.A2(n_263),
.B(n_271),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_290),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_285),
.B(n_243),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_296),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_297),
.B(n_276),
.Y(n_304)
);

AOI31xp67_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_233),
.A3(n_251),
.B(n_243),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_283),
.B(n_288),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_227),
.A3(n_269),
.B1(n_257),
.B2(n_255),
.C1(n_267),
.C2(n_270),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_242),
.B(n_232),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_286),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_272),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_300),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_294),
.A2(n_278),
.B1(n_276),
.B2(n_283),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_305),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_301),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_307),
.B(n_295),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_310),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_289),
.B(n_303),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_298),
.C(n_304),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_311),
.Y(n_315)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_309),
.B(n_307),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_315),
.C(n_300),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_305),
.Y(n_317)
);


endmodule