module fake_aes_8237_n_322 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_322, n_660);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_322;
output n_660;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_575;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_64), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_36), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_69), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_45), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_10), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_67), .Y(n_81) );
INVx1_ASAP7_75t_SL g82 ( .A(n_35), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_51), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_54), .Y(n_84) );
INVxp67_ASAP7_75t_L g85 ( .A(n_37), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_72), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_15), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_27), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_8), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_43), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_13), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_10), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_11), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_75), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_55), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_73), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_24), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_15), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_61), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_17), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_5), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_9), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_70), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_59), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_6), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_11), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_33), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_14), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_17), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_65), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_21), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_19), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_9), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_18), .Y(n_114) );
INVxp33_ASAP7_75t_SL g115 ( .A(n_23), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_34), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_21), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_0), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_71), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_16), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_28), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_47), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_89), .Y(n_123) );
INVx4_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_76), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_94), .B(n_1), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_76), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_77), .Y(n_128) );
BUFx8_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_119), .B(n_1), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_97), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_97), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_78), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_83), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_120), .B(n_2), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_78), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_80), .B(n_2), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_89), .Y(n_141) );
OAI22xp5_ASAP7_75t_SL g142 ( .A1(n_93), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
INVxp67_ASAP7_75t_L g144 ( .A(n_120), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_84), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_80), .B(n_3), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_87), .B(n_4), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_88), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_87), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_88), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_122), .B(n_6), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_90), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g155 ( .A1(n_114), .A2(n_7), .B1(n_8), .B2(n_12), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_98), .B(n_7), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_95), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_96), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_96), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_98), .B(n_12), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_89), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_99), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_107), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_125), .A2(n_106), .B1(n_118), .B2(n_101), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_137), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_137), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_144), .B(n_85), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_144), .B(n_107), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_124), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_125), .B(n_100), .Y(n_172) );
INVx1_ASAP7_75t_SL g173 ( .A(n_131), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_147), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
OAI21xp33_ASAP7_75t_L g177 ( .A1(n_127), .A2(n_111), .B(n_118), .Y(n_177) );
NAND3x1_ASAP7_75t_L g178 ( .A(n_131), .B(n_111), .C(n_101), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_147), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_134), .Y(n_180) );
INVxp67_ASAP7_75t_L g181 ( .A(n_126), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_129), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_127), .B(n_92), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_149), .B(n_108), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_160), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_149), .B(n_164), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_128), .B(n_106), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_134), .Y(n_189) );
BUFx2_ASAP7_75t_L g190 ( .A(n_126), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_164), .B(n_105), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_128), .B(n_116), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_134), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_134), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_130), .B(n_91), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_124), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_130), .B(n_109), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_134), .Y(n_198) );
OR2x2_ASAP7_75t_L g199 ( .A(n_140), .B(n_117), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_135), .B(n_105), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_139), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_139), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_135), .B(n_116), .Y(n_203) );
INVxp67_ASAP7_75t_L g204 ( .A(n_138), .Y(n_204) );
INVxp67_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
INVxp67_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_161), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_145), .B(n_113), .Y(n_208) );
OR2x2_ASAP7_75t_L g209 ( .A(n_140), .B(n_112), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_139), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_150), .Y(n_211) );
AND2x6_ASAP7_75t_L g212 ( .A(n_148), .B(n_110), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_163), .B(n_113), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_148), .B(n_110), .Y(n_214) );
OR2x6_ASAP7_75t_L g215 ( .A(n_142), .B(n_102), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_150), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_129), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_150), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_151), .B(n_115), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_161), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_136), .Y(n_221) );
AND3x4_ASAP7_75t_L g222 ( .A(n_142), .B(n_86), .C(n_112), .Y(n_222) );
OR2x2_ASAP7_75t_L g223 ( .A(n_146), .B(n_102), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_186), .B(n_151), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_186), .B(n_163), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_201), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_186), .A2(n_155), .B1(n_159), .B2(n_153), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_217), .B(n_129), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_217), .B(n_129), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_189), .Y(n_230) );
INVx5_ASAP7_75t_L g231 ( .A(n_170), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_181), .B(n_153), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_174), .B(n_162), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_189), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_212), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_176), .A2(n_162), .B1(n_154), .B2(n_159), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_212), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_221), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_204), .B(n_154), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_212), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_221), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_182), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_179), .B(n_157), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_173), .B(n_146), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_212), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_185), .B(n_157), .Y(n_246) );
BUFx12f_ASAP7_75t_L g247 ( .A(n_215), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_202), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_212), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_184), .B(n_156), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_190), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_187), .Y(n_253) );
INVx1_ASAP7_75t_SL g254 ( .A(n_199), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_209), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_171), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_211), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_216), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_205), .B(n_124), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_215), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_218), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_187), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_187), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_191), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_188), .B(n_156), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_191), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_191), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_200), .Y(n_268) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_165), .B(n_152), .C(n_158), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_206), .B(n_124), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_178), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_219), .B(n_158), .Y(n_272) );
BUFx12f_ASAP7_75t_L g273 ( .A(n_215), .Y(n_273) );
INVx4_ASAP7_75t_L g274 ( .A(n_170), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_200), .B(n_103), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_223), .B(n_121), .Y(n_276) );
INVx2_ASAP7_75t_SL g277 ( .A(n_200), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_168), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_166), .B(n_132), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_171), .Y(n_280) );
INVx5_ASAP7_75t_L g281 ( .A(n_170), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_208), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_208), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_208), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_196), .A2(n_133), .B(n_132), .Y(n_285) );
CKINVDCx11_ASAP7_75t_R g286 ( .A(n_247), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_262), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_261), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_255), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_262), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_225), .B(n_167), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_247), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_231), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g294 ( .A1(n_254), .A2(n_214), .B(n_195), .C(n_183), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_225), .B(n_213), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_245), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_225), .B(n_213), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_278), .A2(n_178), .B1(n_168), .B2(n_213), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_225), .B(n_155), .Y(n_299) );
OAI221xp5_ASAP7_75t_L g300 ( .A1(n_227), .A2(n_165), .B1(n_172), .B2(n_169), .C(n_203), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_262), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_261), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_262), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_274), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_252), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_273), .Y(n_306) );
NOR2xp67_ASAP7_75t_L g307 ( .A(n_227), .B(n_169), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_224), .B(n_265), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_245), .Y(n_309) );
NOR2xp33_ASAP7_75t_R g310 ( .A(n_249), .B(n_197), .Y(n_310) );
OAI33xp33_ASAP7_75t_L g311 ( .A1(n_269), .A2(n_272), .A3(n_244), .B1(n_214), .B2(n_276), .B3(n_177), .Y(n_311) );
NOR2xp67_ASAP7_75t_R g312 ( .A(n_273), .B(n_222), .Y(n_312) );
NOR2xp67_ASAP7_75t_L g313 ( .A(n_260), .B(n_192), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_244), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_250), .B(n_196), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_274), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_284), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_261), .Y(n_318) );
BUFx12f_ASAP7_75t_L g319 ( .A(n_271), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_284), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_245), .Y(n_321) );
UNKNOWN g322 ( );
BUFx3_ASAP7_75t_L g323 ( .A(n_231), .Y(n_323) );
BUFx12f_ASAP7_75t_L g324 ( .A(n_271), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_282), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_253), .A2(n_222), .B1(n_196), .B2(n_82), .Y(n_326) );
INVx4_ASAP7_75t_L g327 ( .A(n_245), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_224), .B(n_133), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_245), .Y(n_329) );
CKINVDCx16_ASAP7_75t_R g330 ( .A(n_282), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_284), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_249), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_261), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_314), .A2(n_268), .B1(n_277), .B2(n_253), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_308), .A2(n_268), .B1(n_277), .B2(n_282), .Y(n_335) );
O2A1O1Ixp33_ASAP7_75t_SL g336 ( .A1(n_288), .A2(n_228), .B(n_229), .C(n_251), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_289), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_308), .A2(n_265), .B1(n_283), .B2(n_264), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_308), .B(n_265), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_286), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_295), .A2(n_283), .B1(n_263), .B2(n_264), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_297), .A2(n_263), .B1(n_266), .B2(n_267), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_291), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_307), .A2(n_266), .B1(n_267), .B2(n_265), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_328), .Y(n_345) );
AO21x2_ASAP7_75t_L g346 ( .A1(n_288), .A2(n_269), .B(n_285), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_299), .A2(n_233), .B1(n_232), .B2(n_279), .Y(n_347) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_319), .A2(n_242), .B1(n_233), .B2(n_235), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_328), .Y(n_349) );
INVxp67_ASAP7_75t_L g350 ( .A(n_305), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_300), .A2(n_246), .B1(n_243), .B2(n_233), .C(n_279), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_315), .A2(n_239), .B1(n_258), .B2(n_226), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_299), .A2(n_249), .B1(n_235), .B2(n_242), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_315), .A2(n_248), .B1(n_226), .B2(n_251), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_328), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_299), .A2(n_279), .B1(n_275), .B2(n_242), .Y(n_356) );
AOI22xp5_ASAP7_75t_SL g357 ( .A1(n_292), .A2(n_248), .B1(n_258), .B2(n_274), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_298), .B(n_257), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_287), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_290), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_301), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_322), .B(n_257), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g363 ( .A(n_293), .B(n_274), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_312), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_337), .A2(n_299), .B1(n_326), .B2(n_330), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_363), .Y(n_366) );
INVx4_ASAP7_75t_SL g367 ( .A(n_339), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_346), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_362), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_352), .A2(n_319), .B1(n_324), .B2(n_325), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_339), .B(n_303), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_363), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_346), .Y(n_373) );
OAI211xp5_ASAP7_75t_L g374 ( .A1(n_347), .A2(n_313), .B(n_286), .C(n_294), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_359), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_358), .B(n_325), .Y(n_376) );
OAI21x1_ASAP7_75t_L g377 ( .A1(n_354), .A2(n_333), .B(n_302), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_359), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_343), .B(n_293), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_351), .A2(n_311), .B1(n_324), .B2(n_331), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_350), .B(n_292), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_344), .A2(n_317), .B(n_320), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_336), .A2(n_333), .B(n_302), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_345), .B(n_306), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_356), .A2(n_310), .B1(n_304), .B2(n_316), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_357), .B(n_323), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_338), .B(n_306), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_349), .B(n_323), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_335), .A2(n_304), .B1(n_316), .B2(n_261), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_355), .A2(n_133), .B1(n_270), .B2(n_259), .C(n_89), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_360), .Y(n_391) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_372), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_375), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_369), .B(n_364), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_365), .A2(n_353), .B1(n_341), .B2(n_342), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_372), .B(n_361), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_369), .B(n_346), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_375), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g399 ( .A(n_380), .B(n_336), .C(n_161), .Y(n_399) );
AOI322xp5_ASAP7_75t_L g400 ( .A1(n_391), .A2(n_340), .A3(n_89), .B1(n_348), .B2(n_104), .C1(n_19), .C2(n_20), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_378), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_379), .Y(n_403) );
AOI222xp33_ASAP7_75t_L g404 ( .A1(n_370), .A2(n_340), .B1(n_304), .B2(n_141), .C1(n_123), .C2(n_143), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_378), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_380), .A2(n_334), .B(n_363), .Y(n_406) );
AO21x2_ASAP7_75t_L g407 ( .A1(n_377), .A2(n_318), .B(n_194), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_391), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_374), .A2(n_318), .B1(n_327), .B2(n_332), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_366), .B(n_13), .Y(n_410) );
AOI211xp5_ASAP7_75t_L g411 ( .A1(n_381), .A2(n_136), .B(n_143), .C(n_141), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_372), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_387), .A2(n_327), .B1(n_332), .B2(n_329), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_368), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_371), .B(n_14), .Y(n_415) );
INVx2_ASAP7_75t_SL g416 ( .A(n_366), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_366), .B(n_327), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_384), .A2(n_136), .B1(n_143), .B2(n_141), .C(n_123), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_371), .B(n_16), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_368), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_386), .B(n_332), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_366), .B(n_18), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
AOI222xp33_ASAP7_75t_L g424 ( .A1(n_367), .A2(n_123), .B1(n_141), .B2(n_136), .C1(n_143), .C2(n_161), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_388), .A2(n_136), .B1(n_143), .B2(n_123), .C(n_161), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_394), .Y(n_426) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_410), .A2(n_386), .B1(n_376), .B2(n_377), .Y(n_427) );
NAND4xp25_ASAP7_75t_L g428 ( .A(n_400), .B(n_385), .C(n_386), .D(n_389), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_397), .B(n_373), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_397), .B(n_373), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_398), .B(n_373), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
OAI33xp33_ASAP7_75t_L g433 ( .A1(n_408), .A2(n_376), .A3(n_368), .B1(n_20), .B2(n_198), .B3(n_194), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_414), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_412), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_402), .B(n_386), .Y(n_436) );
AND2x4_ASAP7_75t_SL g437 ( .A(n_396), .B(n_367), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_400), .B(n_390), .C(n_382), .D(n_383), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_401), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_402), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_403), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_408), .B(n_367), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_414), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_405), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_393), .B(n_367), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_404), .A2(n_136), .B1(n_143), .B2(n_161), .C(n_175), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_423), .B(n_367), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_410), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_405), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_422), .Y(n_450) );
NOR3xp33_ASAP7_75t_SL g451 ( .A(n_419), .B(n_22), .C(n_25), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_420), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_420), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_422), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_393), .B(n_161), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
AOI211xp5_ASAP7_75t_L g457 ( .A1(n_415), .A2(n_136), .B(n_143), .C(n_175), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_407), .Y(n_458) );
AOI22xp33_ASAP7_75t_SL g459 ( .A1(n_392), .A2(n_329), .B1(n_321), .B2(n_309), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_395), .B(n_180), .Y(n_461) );
AOI222xp33_ASAP7_75t_L g462 ( .A1(n_406), .A2(n_180), .B1(n_193), .B2(n_198), .C1(n_231), .C2(n_281), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_421), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_412), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_396), .B(n_193), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_396), .B(n_26), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_396), .Y(n_467) );
INVx5_ASAP7_75t_L g468 ( .A(n_417), .Y(n_468) );
INVx5_ASAP7_75t_SL g469 ( .A(n_417), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_416), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_416), .B(n_256), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_399), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_417), .Y(n_473) );
AND2x2_ASAP7_75t_SL g474 ( .A(n_417), .B(n_329), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_429), .B(n_399), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_467), .B(n_436), .Y(n_476) );
NAND2x2_ASAP7_75t_L g477 ( .A(n_447), .B(n_411), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_439), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_468), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_429), .B(n_409), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_441), .B(n_409), .Y(n_481) );
NAND3xp33_ASAP7_75t_L g482 ( .A(n_457), .B(n_411), .C(n_424), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g483 ( .A(n_433), .B(n_418), .C(n_425), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_431), .B(n_29), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_426), .B(n_413), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_432), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_431), .B(n_30), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_452), .B(n_31), .Y(n_488) );
INVxp67_ASAP7_75t_L g489 ( .A(n_448), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_432), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_440), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_440), .B(n_32), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_430), .B(n_38), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_428), .B(n_438), .C(n_446), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_444), .B(n_39), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_444), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_450), .B(n_40), .Y(n_497) );
NAND2x1p5_ASAP7_75t_L g498 ( .A(n_468), .B(n_321), .Y(n_498) );
NAND3xp33_ASAP7_75t_SL g499 ( .A(n_451), .B(n_41), .C(n_42), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_449), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_452), .B(n_44), .Y(n_501) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_454), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_436), .B(n_46), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_449), .B(n_48), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_434), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_453), .B(n_49), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_453), .B(n_435), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_467), .B(n_50), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_469), .B(n_52), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_434), .Y(n_510) );
NOR2x1_ASAP7_75t_SL g511 ( .A(n_468), .B(n_466), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_443), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_473), .B(n_53), .Y(n_513) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_466), .B(n_321), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_443), .B(n_56), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_442), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_470), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
OAI31xp33_ASAP7_75t_L g519 ( .A1(n_437), .A2(n_237), .A3(n_240), .B(n_256), .Y(n_519) );
OAI31xp33_ASAP7_75t_L g520 ( .A1(n_437), .A2(n_237), .A3(n_240), .B(n_256), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_469), .B(n_57), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_469), .B(n_58), .Y(n_522) );
BUFx2_ASAP7_75t_L g523 ( .A(n_468), .Y(n_523) );
AOI211xp5_ASAP7_75t_L g524 ( .A1(n_445), .A2(n_220), .B(n_207), .C(n_309), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_468), .B(n_60), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_456), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_445), .B(n_62), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_445), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_458), .B(n_63), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_478), .B(n_464), .Y(n_530) );
AOI21xp33_ASAP7_75t_SL g531 ( .A1(n_494), .A2(n_474), .B(n_427), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_507), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_486), .Y(n_533) );
OAI22xp33_ASAP7_75t_R g534 ( .A1(n_502), .A2(n_472), .B1(n_464), .B2(n_463), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_476), .B(n_489), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_516), .B(n_472), .Y(n_536) );
NOR2x1p5_ASAP7_75t_L g537 ( .A(n_479), .B(n_458), .Y(n_537) );
NOR2x1_ASAP7_75t_L g538 ( .A(n_479), .B(n_471), .Y(n_538) );
OAI21xp33_ASAP7_75t_L g539 ( .A1(n_481), .A2(n_461), .B(n_462), .Y(n_539) );
OAI21xp33_ASAP7_75t_L g540 ( .A1(n_485), .A2(n_455), .B(n_465), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_490), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_491), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_496), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_500), .B(n_455), .Y(n_544) );
XOR2xp5_ASAP7_75t_L g545 ( .A(n_511), .B(n_474), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_517), .B(n_460), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_518), .B(n_456), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_505), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_526), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_505), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_510), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_510), .B(n_471), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_512), .Y(n_553) );
AO21x1_ASAP7_75t_SL g554 ( .A1(n_528), .A2(n_459), .B(n_68), .Y(n_554) );
CKINVDCx8_ASAP7_75t_R g555 ( .A(n_523), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_480), .B(n_66), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_480), .B(n_74), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_484), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_475), .B(n_207), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_475), .B(n_220), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_483), .B(n_231), .C(n_281), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_524), .A2(n_309), .B(n_296), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_526), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_482), .B(n_231), .C(n_281), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_512), .B(n_231), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_514), .B(n_309), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_477), .A2(n_296), .B1(n_281), .B2(n_230), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_484), .B(n_281), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_527), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_529), .B(n_230), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_504), .Y(n_571) );
OAI21xp5_ASAP7_75t_L g572 ( .A1(n_499), .A2(n_281), .B(n_237), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_487), .B(n_234), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_493), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_493), .Y(n_575) );
OAI21xp33_ASAP7_75t_L g576 ( .A1(n_535), .A2(n_503), .B(n_497), .Y(n_576) );
INVxp67_ASAP7_75t_SL g577 ( .A(n_538), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_532), .B(n_529), .Y(n_578) );
XOR2xp5_ASAP7_75t_L g579 ( .A(n_545), .B(n_521), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_552), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_536), .B(n_487), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_533), .Y(n_582) );
INVxp67_ASAP7_75t_L g583 ( .A(n_530), .Y(n_583) );
AND2x4_ASAP7_75t_L g584 ( .A(n_537), .B(n_527), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_SL g585 ( .A1(n_531), .A2(n_522), .B(n_509), .C(n_525), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_569), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_541), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_548), .B(n_551), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_550), .B(n_508), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_542), .B(n_501), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_543), .B(n_488), .Y(n_591) );
OR2x6_ASAP7_75t_L g592 ( .A(n_569), .B(n_527), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_544), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_574), .B(n_488), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_558), .B(n_513), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_575), .B(n_515), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_546), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_547), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_553), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_549), .Y(n_600) );
OAI31xp33_ASAP7_75t_L g601 ( .A1(n_561), .A2(n_520), .A3(n_519), .B(n_498), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_571), .B(n_539), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_558), .B(n_495), .Y(n_603) );
AND3x2_ASAP7_75t_L g604 ( .A(n_534), .B(n_477), .C(n_506), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_563), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_565), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_559), .B(n_492), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_555), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_555), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_540), .A2(n_498), .B1(n_280), .B2(n_238), .C(n_234), .Y(n_610) );
A2O1A1Ixp33_ASAP7_75t_L g611 ( .A1(n_562), .A2(n_237), .B(n_240), .C(n_296), .Y(n_611) );
OAI21xp5_ASAP7_75t_L g612 ( .A1(n_567), .A2(n_240), .B(n_238), .Y(n_612) );
OA22x2_ASAP7_75t_L g613 ( .A1(n_556), .A2(n_566), .B1(n_557), .B2(n_568), .Y(n_613) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_560), .A2(n_241), .B(n_280), .Y(n_614) );
NAND4xp25_ASAP7_75t_L g615 ( .A(n_567), .B(n_241), .C(n_280), .D(n_572), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_573), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_570), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_566), .Y(n_618) );
XOR2xp5_ASAP7_75t_L g619 ( .A(n_554), .B(n_280), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_539), .A2(n_280), .B1(n_494), .B2(n_477), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_533), .Y(n_621) );
A2O1A1Ixp33_ASAP7_75t_L g622 ( .A1(n_531), .A2(n_537), .B(n_400), .C(n_538), .Y(n_622) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_538), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_534), .A2(n_494), .B1(n_539), .B2(n_569), .Y(n_624) );
NOR3xp33_ASAP7_75t_L g625 ( .A(n_531), .B(n_561), .C(n_564), .Y(n_625) );
OAI211xp5_ASAP7_75t_L g626 ( .A1(n_624), .A2(n_620), .B(n_601), .C(n_622), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_625), .A2(n_602), .B1(n_613), .B2(n_616), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_609), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_608), .B(n_580), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g630 ( .A1(n_583), .A2(n_593), .B1(n_623), .B2(n_577), .C1(n_597), .C2(n_598), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_588), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_584), .A2(n_577), .B(n_576), .C(n_615), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_604), .B(n_617), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_579), .B(n_604), .Y(n_634) );
AOI211x1_ASAP7_75t_SL g635 ( .A1(n_603), .A2(n_578), .B(n_589), .C(n_581), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_600), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_585), .B(n_618), .C(n_610), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_613), .A2(n_585), .B1(n_584), .B2(n_586), .Y(n_638) );
AOI211xp5_ASAP7_75t_SL g639 ( .A1(n_584), .A2(n_610), .B(n_595), .C(n_611), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_628), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g641 ( .A1(n_626), .A2(n_592), .B1(n_587), .B2(n_582), .C(n_621), .Y(n_641) );
OAI211xp5_ASAP7_75t_SL g642 ( .A1(n_627), .A2(n_612), .B(n_591), .C(n_590), .Y(n_642) );
NOR2x1_ASAP7_75t_L g643 ( .A(n_634), .B(n_592), .Y(n_643) );
NOR4xp75_ASAP7_75t_L g644 ( .A(n_633), .B(n_594), .C(n_596), .D(n_612), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_631), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_629), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g647 ( .A(n_637), .B(n_614), .C(n_606), .Y(n_647) );
OAI211xp5_ASAP7_75t_L g648 ( .A1(n_643), .A2(n_627), .B(n_634), .C(n_638), .Y(n_648) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_642), .B(n_632), .C(n_639), .Y(n_649) );
OAI22x1_ASAP7_75t_L g650 ( .A1(n_640), .A2(n_630), .B1(n_635), .B2(n_619), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_640), .Y(n_651) );
NOR3xp33_ASAP7_75t_L g652 ( .A(n_648), .B(n_641), .C(n_647), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_651), .B(n_646), .Y(n_653) );
NOR3xp33_ASAP7_75t_L g654 ( .A(n_649), .B(n_645), .C(n_644), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_653), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_654), .Y(n_656) );
AO21x2_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_652), .B(n_655), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_657), .Y(n_658) );
OR3x2_ASAP7_75t_L g659 ( .A(n_658), .B(n_657), .C(n_650), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_659), .A2(n_636), .B1(n_607), .B2(n_599), .C(n_605), .Y(n_660) );
endmodule