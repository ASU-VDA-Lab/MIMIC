module real_jpeg_24072_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_2),
.A2(n_19),
.B1(n_20),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_2),
.A2(n_41),
.B1(n_43),
.B2(n_48),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_5),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_5),
.A2(n_19),
.B1(n_20),
.B2(n_26),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_5),
.A2(n_26),
.B1(n_41),
.B2(n_43),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_8),
.A2(n_24),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_8),
.A2(n_33),
.B1(n_41),
.B2(n_43),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_8),
.A2(n_18),
.B(n_27),
.C(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_8),
.B(n_16),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_8),
.A2(n_19),
.B1(n_20),
.B2(n_33),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_8),
.B(n_39),
.C(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_8),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_8),
.B(n_37),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_77),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_75),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_59),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_12),
.B(n_59),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_49),
.Y(n_12)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_34),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_28),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_23),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_17)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_18),
.A2(n_22),
.B1(n_24),
.B2(n_27),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_19),
.A2(n_20),
.B1(n_38),
.B2(n_39),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_19),
.A2(n_22),
.B(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_85),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_44),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_47),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_41),
.B(n_103),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_45),
.B(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_56),
.B2(n_58),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B(n_55),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_73),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_52),
.B(n_55),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_94),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_56),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.C(n_65),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_65),
.A2(n_66),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_90),
.B(n_114),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_86),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_79),
.B(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_83),
.B1(n_84),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_100),
.B(n_113),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_108),
.B(n_112),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_109),
.B(n_110),
.Y(n_112)
);


endmodule