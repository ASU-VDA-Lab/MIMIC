module fake_jpeg_732_n_101 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_49),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_35),
.B1(n_27),
.B2(n_29),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_38),
.B(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_30),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_37),
.B1(n_40),
.B2(n_35),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_55),
.B1(n_48),
.B2(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_56),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_37),
.B1(n_47),
.B2(n_43),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_47),
.B1(n_49),
.B2(n_42),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_42),
.B1(n_34),
.B2(n_38),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_67),
.B(n_3),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_65),
.B(n_68),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_15),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_1),
.C(n_2),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_38),
.B1(n_2),
.B2(n_3),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_74),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_77),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_56),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_75),
.C(n_16),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_57),
.C(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

AOI32xp33_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_80),
.B(n_86),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_19),
.B1(n_25),
.B2(n_24),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_26),
.B(n_23),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_91),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_83),
.C(n_85),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_90),
.C(n_80),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_88),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_94),
.C(n_20),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_22),
.C(n_10),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_10),
.C(n_11),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_11),
.Y(n_101)
);


endmodule