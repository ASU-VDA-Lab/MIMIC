module fake_jpeg_26823_n_113 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_113);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_113;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_SL g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_1),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_14),
.A2(n_1),
.B(n_2),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_3),
.B(n_4),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_1),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_33),
.Y(n_39)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_18),
.Y(n_40)
);

CKINVDCx9p33_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_29),
.B1(n_31),
.B2(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_24),
.B1(n_16),
.B2(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_44),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_24),
.B1(n_16),
.B2(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_44),
.Y(n_59)
);

NOR2x1_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_21),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_60),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_54),
.B(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_34),
.B(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_15),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_39),
.B(n_36),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_74),
.B(n_43),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_41),
.B1(n_35),
.B2(n_39),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_67),
.B1(n_54),
.B2(n_57),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_38),
.B1(n_24),
.B2(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_70),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_R g70 ( 
.A(n_50),
.B(n_21),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_42),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_27),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_38),
.C(n_27),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_38),
.C(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_78),
.C(n_79),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_52),
.B(n_58),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_52),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_42),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_45),
.B1(n_28),
.B2(n_43),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_72),
.C(n_61),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_73),
.B(n_62),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_85),
.B(n_22),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_68),
.A3(n_63),
.B1(n_62),
.B2(n_66),
.C1(n_11),
.C2(n_12),
.Y(n_87)
);

OA21x2_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_89),
.B(n_93),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_79),
.C(n_78),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_11),
.C(n_81),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_61),
.B1(n_74),
.B2(n_45),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_27),
.C(n_26),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_76),
.C(n_82),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_30),
.B1(n_28),
.B2(n_22),
.Y(n_92)
);

INVxp33_ASAP7_75t_SL g94 ( 
.A(n_90),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_96),
.C(n_97),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_27),
.C(n_26),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_98),
.A2(n_95),
.B1(n_99),
.B2(n_20),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_26),
.C(n_21),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_26),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_26),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_3),
.B(n_4),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_6),
.B(n_7),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_104),
.B(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_6),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_107),
.B(n_103),
.CI(n_101),
.CON(n_109),
.SN(n_109)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_108),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_110),
.B1(n_109),
.B2(n_10),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_10),
.Y(n_113)
);


endmodule