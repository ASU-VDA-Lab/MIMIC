module fake_netlist_6_476_n_1719 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1719);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1719;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_108),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_32),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_10),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_139),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_14),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_27),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_34),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_21),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_24),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_72),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_97),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_98),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_67),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_119),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_109),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_118),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_48),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_40),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_40),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_29),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_13),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_29),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_70),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_18),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_64),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_88),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_39),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_60),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_124),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_94),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_135),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_23),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_36),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_133),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_7),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_46),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_16),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_103),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_87),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_106),
.Y(n_215)
);

INVx2_ASAP7_75t_R g216 ( 
.A(n_49),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_75),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_91),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_102),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_48),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_25),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_57),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_13),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_128),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_46),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_68),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_110),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_36),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_62),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_16),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_45),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_47),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_65),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_113),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_144),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_58),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_89),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_126),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_10),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_54),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_7),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_42),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_61),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_38),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_21),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_66),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_1),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_82),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_37),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_31),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_92),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_105),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_130),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_34),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_101),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_43),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_8),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_42),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_23),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_31),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_47),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_30),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_150),
.Y(n_265)
);

BUFx8_ASAP7_75t_SL g266 ( 
.A(n_83),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_81),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_41),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_51),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_39),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_95),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_84),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_149),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_116),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_32),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_30),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_63),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_96),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g279 ( 
.A(n_156),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_129),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_107),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_45),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_8),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_120),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_15),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_148),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_69),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_137),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_132),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_4),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_143),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_93),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_111),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_77),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_14),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_35),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_18),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_17),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_125),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_99),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_5),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_43),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_15),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_22),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_85),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_38),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_24),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_2),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_4),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_54),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_78),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_76),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_210),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_210),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_209),
.B(n_0),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_221),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_221),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_258),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_194),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_258),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_200),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_182),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_159),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_209),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_205),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_260),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_266),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_285),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_158),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_163),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_267),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_287),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_265),
.B(n_0),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_164),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_290),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_207),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_265),
.B(n_1),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_280),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_168),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_178),
.B(n_236),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_208),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_177),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_180),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_290),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_298),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_298),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_162),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_207),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_204),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_184),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_185),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_186),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_162),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_199),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_196),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_201),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_199),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_213),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_223),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_223),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_224),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_224),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_214),
.Y(n_367)
);

BUFx2_ASAP7_75t_SL g368 ( 
.A(n_187),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_215),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_226),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_226),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_229),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_229),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_218),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_219),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_220),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_227),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_160),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_230),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_233),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_233),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_240),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_237),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_240),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_242),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_166),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_244),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_242),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_322),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_340),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_386),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_315),
.B(n_204),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_378),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_322),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_336),
.B(n_204),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_216),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_316),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

BUFx8_ASAP7_75t_L g400 ( 
.A(n_353),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_322),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_368),
.B(n_187),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_322),
.B(n_178),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_313),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_341),
.B(n_204),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_351),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_313),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_357),
.A2(n_253),
.B(n_236),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_353),
.B(n_235),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_314),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_314),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_352),
.B(n_235),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_368),
.B(n_252),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_352),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_317),
.Y(n_416)
);

AND3x2_ASAP7_75t_L g417 ( 
.A(n_324),
.B(n_255),
.C(n_253),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_357),
.B(n_271),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_358),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_317),
.B(n_216),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_318),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_318),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_320),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_320),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_332),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_358),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_361),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_361),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_326),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_363),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_326),
.B(n_216),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_342),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_364),
.B(n_273),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_L g435 ( 
.A(n_364),
.B(n_275),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_365),
.B(n_274),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_327),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_365),
.B(n_281),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_327),
.B(n_192),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_323),
.B(n_197),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_366),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_366),
.Y(n_442)
);

NAND2xp33_ASAP7_75t_SL g443 ( 
.A(n_360),
.B(n_275),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_321),
.A2(n_232),
.B1(n_174),
.B2(n_170),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_329),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_329),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_330),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_370),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_370),
.B(n_257),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_330),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_331),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_371),
.B(n_288),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_331),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_372),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_338),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_369),
.A2(n_246),
.B1(n_222),
.B2(n_212),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_338),
.B(n_192),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_372),
.B(n_373),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_403),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_403),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_408),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_393),
.A2(n_276),
.B1(n_193),
.B2(n_310),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_440),
.B(n_333),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_403),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_408),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_403),
.Y(n_468)
);

AO22x2_ASAP7_75t_L g469 ( 
.A1(n_393),
.A2(n_276),
.B1(n_264),
.B2(n_262),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_396),
.B(n_375),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_403),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_403),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_414),
.B(n_337),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_395),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_426),
.B(n_339),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_408),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_394),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_395),
.Y(n_478)
);

BUFx10_ASAP7_75t_L g479 ( 
.A(n_440),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_397),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_433),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_395),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_397),
.B(n_420),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_397),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_420),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

AO22x2_ASAP7_75t_L g488 ( 
.A1(n_396),
.A2(n_406),
.B1(n_413),
.B2(n_410),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_SL g490 ( 
.A(n_406),
.B(n_376),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_411),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_433),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_420),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_414),
.B(n_343),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_395),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_444),
.A2(n_173),
.B1(n_270),
.B2(n_297),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_411),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_395),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_394),
.B(n_346),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_426),
.B(n_339),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_426),
.B(n_348),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_415),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_425),
.B(n_347),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_432),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_432),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_418),
.B(n_354),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_401),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_411),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_391),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_432),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_405),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_402),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_418),
.B(n_355),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_405),
.Y(n_515)
);

BUFx8_ASAP7_75t_SL g516 ( 
.A(n_391),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_410),
.B(n_356),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

OAI22xp33_ASAP7_75t_L g519 ( 
.A1(n_457),
.A2(n_283),
.B1(n_172),
.B2(n_188),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_411),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_407),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_419),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_402),
.B(n_359),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_439),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_401),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_434),
.B(n_362),
.Y(n_526)
);

INVxp33_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_425),
.B(n_367),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_422),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_434),
.B(n_374),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_409),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_436),
.B(n_377),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_419),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_422),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_449),
.A2(n_193),
.B1(n_262),
.B2(n_301),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_449),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_425),
.B(n_279),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_427),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_436),
.B(n_379),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_422),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_444),
.A2(n_413),
.B1(n_457),
.B2(n_443),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_427),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_409),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_421),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_425),
.B(n_383),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_428),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_428),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_423),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_423),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_438),
.B(n_387),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_425),
.B(n_345),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_400),
.B(n_328),
.Y(n_553)
);

BUFx8_ASAP7_75t_SL g554 ( 
.A(n_391),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_423),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_438),
.B(n_453),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_429),
.Y(n_557)
);

BUFx8_ASAP7_75t_SL g558 ( 
.A(n_453),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_402),
.A2(n_261),
.B1(n_248),
.B2(n_245),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_429),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_439),
.B(n_458),
.Y(n_561)
);

BUFx4f_ASAP7_75t_L g562 ( 
.A(n_449),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_392),
.B(n_325),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_431),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_449),
.A2(n_301),
.B1(n_264),
.B2(n_282),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_401),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_423),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_439),
.B(n_458),
.Y(n_568)
);

INVx4_ASAP7_75t_SL g569 ( 
.A(n_449),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_421),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_390),
.B(n_228),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_449),
.B(n_257),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_400),
.B(n_235),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_431),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_400),
.B(n_235),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_401),
.Y(n_576)
);

OAI21xp33_ASAP7_75t_SL g577 ( 
.A1(n_409),
.A2(n_310),
.B(n_309),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_458),
.B(n_381),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_400),
.B(n_289),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_459),
.B(n_279),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_400),
.B(n_292),
.Y(n_581)
);

NOR3xp33_ASAP7_75t_L g582 ( 
.A(n_443),
.B(n_382),
.C(n_385),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_417),
.B(n_334),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_441),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_389),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_421),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_441),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_435),
.A2(n_442),
.B1(n_455),
.B2(n_452),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_389),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_437),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_437),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_442),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_390),
.B(n_293),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_459),
.B(n_384),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_437),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_448),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_437),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_448),
.B(n_373),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_445),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_445),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_417),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_445),
.Y(n_602)
);

BUFx4f_ASAP7_75t_L g603 ( 
.A(n_421),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_390),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_412),
.B(n_348),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_400),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_445),
.Y(n_607)
);

BUFx4f_ASAP7_75t_L g608 ( 
.A(n_421),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_452),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_481),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_477),
.B(n_404),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_556),
.B(n_404),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_499),
.B(n_404),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_463),
.B(n_435),
.C(n_251),
.Y(n_614)
);

NOR2x1_ASAP7_75t_L g615 ( 
.A(n_538),
.B(n_335),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_486),
.B(n_182),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_510),
.B(n_455),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_481),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_513),
.B(n_243),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_486),
.B(n_182),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_462),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_511),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_485),
.B(n_404),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_513),
.B(n_189),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_485),
.B(n_404),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_493),
.B(n_182),
.Y(n_626)
);

OAI22xp33_ASAP7_75t_L g627 ( 
.A1(n_542),
.A2(n_594),
.B1(n_568),
.B2(n_580),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_511),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_484),
.B(n_424),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_531),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_493),
.B(n_182),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_488),
.A2(n_294),
.B1(n_299),
.B2(n_305),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_512),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_601),
.B(n_282),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_601),
.B(n_307),
.Y(n_635)
);

BUFx6f_ASAP7_75t_SL g636 ( 
.A(n_479),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_482),
.B(n_243),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_523),
.B(n_190),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_505),
.A2(n_506),
.B1(n_484),
.B2(n_469),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_484),
.B(n_424),
.Y(n_640)
);

BUFx4f_ASAP7_75t_L g641 ( 
.A(n_523),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_531),
.B(n_160),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_505),
.B(n_225),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_512),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_515),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_506),
.B(n_225),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_510),
.B(n_380),
.Y(n_647)
);

BUFx8_ASAP7_75t_L g648 ( 
.A(n_578),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_484),
.B(n_424),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_515),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_518),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_484),
.B(n_424),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_484),
.B(n_424),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_462),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_484),
.B(n_430),
.Y(n_655)
);

INVxp67_ASAP7_75t_SL g656 ( 
.A(n_531),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_507),
.B(n_430),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_514),
.B(n_430),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_518),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_526),
.B(n_195),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_572),
.B(n_225),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_530),
.B(n_206),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_537),
.B(n_562),
.Y(n_663)
);

OAI221xp5_ASAP7_75t_L g664 ( 
.A1(n_565),
.A2(n_307),
.B1(n_309),
.B2(n_239),
.C(n_234),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_467),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_521),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_537),
.B(n_225),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_562),
.A2(n_389),
.B(n_454),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_578),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_562),
.A2(n_389),
.B(n_454),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_532),
.B(n_430),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_540),
.B(n_430),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_561),
.B(n_524),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_537),
.B(n_225),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_521),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_551),
.B(n_211),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_475),
.Y(n_677)
);

OR2x6_ASAP7_75t_SL g678 ( 
.A(n_473),
.B(n_231),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_524),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_594),
.B(n_241),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_460),
.B(n_286),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_561),
.B(n_380),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_503),
.B(n_161),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_460),
.B(n_286),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_461),
.B(n_286),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_542),
.A2(n_179),
.B(n_161),
.C(n_312),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_522),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_582),
.B(n_256),
.C(n_250),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_494),
.B(n_446),
.Y(n_689)
);

AO221x1_ASAP7_75t_L g690 ( 
.A1(n_488),
.A2(n_286),
.B1(n_165),
.B2(n_239),
.C(n_167),
.Y(n_690)
);

OAI221xp5_ASAP7_75t_L g691 ( 
.A1(n_536),
.A2(n_176),
.B1(n_312),
.B2(n_300),
.C(n_291),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_522),
.B(n_446),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_461),
.B(n_286),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_534),
.B(n_446),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_L g695 ( 
.A1(n_577),
.A2(n_175),
.B(n_165),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_534),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_539),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_539),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_464),
.B(n_259),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_543),
.B(n_547),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_604),
.Y(n_701)
);

AOI22x1_ASAP7_75t_L g702 ( 
.A1(n_488),
.A2(n_311),
.B1(n_238),
.B2(n_234),
.Y(n_702)
);

AO221x1_ASAP7_75t_L g703 ( 
.A1(n_488),
.A2(n_171),
.B1(n_167),
.B2(n_169),
.C(n_175),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_543),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_479),
.B(n_243),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_476),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_466),
.B(n_311),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_598),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_466),
.B(n_421),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_475),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_547),
.Y(n_711)
);

NOR3xp33_ASAP7_75t_L g712 ( 
.A(n_563),
.B(n_269),
.C(n_263),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_572),
.B(n_169),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_548),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_548),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_476),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_468),
.B(n_421),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_568),
.A2(n_171),
.B(n_176),
.C(n_179),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_557),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_557),
.B(n_446),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_468),
.B(n_421),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_560),
.Y(n_722)
);

AND2x6_ASAP7_75t_SL g723 ( 
.A(n_583),
.B(n_388),
.Y(n_723)
);

NOR2x1p5_ASAP7_75t_L g724 ( 
.A(n_598),
.B(n_295),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_479),
.B(n_296),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_560),
.B(n_446),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_604),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_492),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_564),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_479),
.B(n_243),
.Y(n_730)
);

INVxp33_ASAP7_75t_SL g731 ( 
.A(n_504),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_564),
.B(n_181),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_469),
.A2(n_300),
.B1(n_183),
.B2(n_191),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_574),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_574),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_527),
.B(n_559),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_584),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_584),
.B(n_198),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_500),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_587),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_587),
.B(n_198),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_517),
.B(n_302),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_592),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_487),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_471),
.A2(n_202),
.B1(n_203),
.B2(n_217),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_471),
.B(n_202),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_491),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_592),
.B(n_203),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_491),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_497),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_497),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_472),
.B(n_217),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_596),
.B(n_238),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_496),
.B(n_388),
.Y(n_754)
);

NOR2x1p5_ASAP7_75t_L g755 ( 
.A(n_596),
.B(n_303),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_609),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_472),
.B(n_247),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_609),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_528),
.B(n_247),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_500),
.Y(n_760)
);

BUFx5_ASAP7_75t_L g761 ( 
.A(n_572),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_546),
.B(n_304),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_502),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_502),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_577),
.A2(n_249),
.B(n_254),
.C(n_272),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_538),
.A2(n_249),
.B1(n_254),
.B2(n_272),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_519),
.B(n_308),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_571),
.B(n_277),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_580),
.B(n_277),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_572),
.B(n_278),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_580),
.B(n_278),
.Y(n_771)
);

NAND3xp33_ASAP7_75t_SL g772 ( 
.A(n_496),
.B(n_306),
.C(n_291),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_580),
.B(n_284),
.Y(n_773)
);

O2A1O1Ixp5_ASAP7_75t_L g774 ( 
.A1(n_593),
.A2(n_284),
.B(n_454),
.C(n_451),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_605),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_531),
.B(n_447),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_509),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_531),
.B(n_544),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_509),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_673),
.B(n_469),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_L g781 ( 
.A(n_630),
.B(n_606),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_762),
.A2(n_470),
.B(n_490),
.C(n_552),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_680),
.B(n_669),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_627),
.A2(n_662),
.B1(n_676),
.B2(n_660),
.Y(n_784)
);

OAI21xp33_ASAP7_75t_L g785 ( 
.A1(n_680),
.A2(n_588),
.B(n_580),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_762),
.B(n_544),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_618),
.B(n_544),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_679),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_679),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_778),
.A2(n_544),
.B(n_608),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_630),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_731),
.B(n_728),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_778),
.A2(n_544),
.B(n_608),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_622),
.B(n_606),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_617),
.B(n_605),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_628),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_708),
.B(n_647),
.Y(n_797)
);

AO21x1_ASAP7_75t_L g798 ( 
.A1(n_695),
.A2(n_573),
.B(n_575),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_639),
.A2(n_538),
.B1(n_581),
.B2(n_579),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_610),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_686),
.A2(n_538),
.B(n_553),
.C(n_602),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_622),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_660),
.B(n_558),
.Y(n_803)
);

BUFx2_ASAP7_75t_SL g804 ( 
.A(n_636),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_754),
.B(n_538),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_622),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_677),
.B(n_349),
.Y(n_807)
);

O2A1O1Ixp5_ASAP7_75t_L g808 ( 
.A1(n_667),
.A2(n_608),
.B(n_603),
.C(n_501),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_676),
.B(n_516),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_656),
.A2(n_603),
.B(n_498),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_633),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_619),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_663),
.A2(n_611),
.B(n_629),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_686),
.A2(n_607),
.B(n_602),
.C(n_600),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_725),
.B(n_554),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_618),
.B(n_501),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_622),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_644),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_612),
.B(n_501),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_630),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_710),
.B(n_349),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_776),
.A2(n_674),
.B(n_667),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_776),
.A2(n_603),
.B(n_480),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_701),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_634),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_739),
.B(n_508),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_648),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_699),
.A2(n_767),
.B(n_742),
.C(n_759),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_613),
.A2(n_658),
.B(n_657),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_701),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_671),
.A2(n_672),
.B(n_663),
.Y(n_831)
);

AOI22x1_ASAP7_75t_L g832 ( 
.A1(n_645),
.A2(n_525),
.B1(n_566),
.B2(n_508),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_725),
.B(n_525),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_760),
.B(n_566),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_763),
.B(n_576),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_764),
.B(n_576),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_650),
.B(n_651),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_659),
.B(n_576),
.Y(n_838)
);

AO21x1_ASAP7_75t_L g839 ( 
.A1(n_766),
.A2(n_586),
.B(n_600),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_666),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_675),
.B(n_465),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_638),
.B(n_767),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_727),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_687),
.B(n_696),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_630),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_627),
.A2(n_699),
.B1(n_632),
.B2(n_638),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_697),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_698),
.B(n_465),
.Y(n_848)
);

NAND2x1p5_ASAP7_75t_L g849 ( 
.A(n_727),
.B(n_480),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_705),
.B(n_350),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_682),
.A2(n_572),
.B1(n_569),
.B2(n_465),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_730),
.B(n_624),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_704),
.B(n_474),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_641),
.B(n_569),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_682),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_SL g856 ( 
.A(n_641),
.B(n_572),
.Y(n_856)
);

NOR3xp33_ASAP7_75t_L g857 ( 
.A(n_772),
.B(n_450),
.C(n_456),
.Y(n_857)
);

OR2x6_ASAP7_75t_SL g858 ( 
.A(n_736),
.B(n_350),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_642),
.Y(n_859)
);

AO21x2_ASAP7_75t_L g860 ( 
.A1(n_690),
.A2(n_607),
.B(n_599),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_624),
.B(n_480),
.Y(n_861)
);

O2A1O1Ixp5_ASAP7_75t_L g862 ( 
.A1(n_674),
.A2(n_474),
.B(n_478),
.C(n_495),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_775),
.B(n_412),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_640),
.A2(n_474),
.B(n_478),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_711),
.B(n_478),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_742),
.A2(n_649),
.B1(n_652),
.B2(n_653),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_655),
.A2(n_495),
.B(n_597),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_689),
.A2(n_498),
.B(n_489),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_714),
.B(n_495),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_639),
.A2(n_599),
.B1(n_597),
.B2(n_595),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_715),
.B(n_572),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_623),
.A2(n_498),
.B(n_489),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_769),
.A2(n_595),
.B(n_591),
.C(n_590),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_771),
.A2(n_591),
.B(n_590),
.C(n_533),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_615),
.B(n_700),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_625),
.A2(n_489),
.B(n_483),
.Y(n_876)
);

BUFx8_ASAP7_75t_L g877 ( 
.A(n_636),
.Y(n_877)
);

NOR3xp33_ASAP7_75t_L g878 ( 
.A(n_688),
.B(n_456),
.C(n_416),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_719),
.B(n_483),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_722),
.B(n_483),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_761),
.B(n_569),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_661),
.A2(n_717),
.B(n_709),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_773),
.A2(n_765),
.B(n_752),
.C(n_757),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_709),
.A2(n_586),
.B(n_533),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_729),
.A2(n_569),
.B1(n_586),
.B2(n_585),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_734),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_634),
.B(n_412),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_735),
.B(n_529),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_SL g889 ( 
.A(n_637),
.B(n_450),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_717),
.A2(n_529),
.B(n_520),
.Y(n_890)
);

O2A1O1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_765),
.A2(n_567),
.B(n_555),
.C(n_550),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_621),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_683),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_737),
.Y(n_894)
);

INVx11_ASAP7_75t_L g895 ( 
.A(n_648),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_721),
.A2(n_535),
.B(n_520),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_654),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_755),
.B(n_456),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_721),
.A2(n_541),
.B(n_535),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_702),
.A2(n_541),
.B1(n_549),
.B2(n_567),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_692),
.A2(n_555),
.B(n_550),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_740),
.B(n_549),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_694),
.A2(n_589),
.B(n_585),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_743),
.B(n_589),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_720),
.A2(n_726),
.B(n_707),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_707),
.A2(n_589),
.B(n_585),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_634),
.B(n_589),
.Y(n_907)
);

INVx4_ASAP7_75t_L g908 ( 
.A(n_761),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_756),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_758),
.B(n_589),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_665),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_768),
.B(n_585),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_635),
.B(n_416),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_642),
.B(n_585),
.Y(n_914)
);

AO21x1_ASAP7_75t_L g915 ( 
.A1(n_616),
.A2(n_450),
.B(n_416),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_616),
.A2(n_570),
.B(n_545),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_718),
.A2(n_399),
.B(n_398),
.C(n_454),
.Y(n_917)
);

BUFx4f_ASAP7_75t_L g918 ( 
.A(n_635),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_620),
.A2(n_570),
.B(n_545),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_774),
.A2(n_620),
.B(n_626),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_724),
.B(n_398),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_631),
.A2(n_570),
.B(n_545),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_635),
.B(n_2),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_761),
.B(n_399),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_643),
.A2(n_570),
.B(n_545),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_683),
.B(n_451),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_642),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_642),
.B(n_451),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_646),
.A2(n_447),
.B(n_152),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_761),
.B(n_447),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_683),
.B(n_3),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_712),
.B(n_3),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_646),
.A2(n_145),
.B(n_140),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_642),
.B(n_5),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_706),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_668),
.A2(n_134),
.B(n_123),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_732),
.B(n_6),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_738),
.B(n_9),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_670),
.A2(n_121),
.B(n_117),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_713),
.A2(n_770),
.B(n_752),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_746),
.A2(n_115),
.B(n_114),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_746),
.A2(n_112),
.B(n_86),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_757),
.A2(n_80),
.B(n_79),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_681),
.A2(n_74),
.B(n_59),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_681),
.A2(n_685),
.B(n_693),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_684),
.A2(n_11),
.B(n_12),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_741),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_723),
.B(n_11),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_716),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_748),
.B(n_753),
.Y(n_950)
);

AOI21xp33_ASAP7_75t_L g951 ( 
.A1(n_733),
.A2(n_12),
.B(n_17),
.Y(n_951)
);

AO21x1_ASAP7_75t_L g952 ( 
.A1(n_684),
.A2(n_19),
.B(n_20),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_685),
.A2(n_19),
.B(n_20),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_691),
.A2(n_22),
.B(n_25),
.C(n_26),
.Y(n_954)
);

INVx11_ASAP7_75t_L g955 ( 
.A(n_678),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_744),
.B(n_26),
.Y(n_956)
);

OAI321xp33_ASAP7_75t_L g957 ( 
.A1(n_664),
.A2(n_27),
.A3(n_28),
.B1(n_33),
.B2(n_37),
.C(n_41),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_747),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_614),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_693),
.B(n_28),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_749),
.B(n_33),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_R g962 ( 
.A(n_750),
.B(n_44),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_751),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_825),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_820),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_820),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_877),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_842),
.A2(n_745),
.B(n_777),
.C(n_779),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_901),
.A2(n_703),
.B(n_49),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_858),
.Y(n_970)
);

OAI21x1_ASAP7_75t_L g971 ( 
.A1(n_901),
.A2(n_44),
.B(n_50),
.Y(n_971)
);

NAND2x1_ASAP7_75t_L g972 ( 
.A(n_820),
.B(n_50),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_949),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_852),
.B(n_51),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_792),
.B(n_52),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_784),
.A2(n_52),
.B(n_53),
.C(n_55),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_963),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_963),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_828),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_979)
);

BUFx8_ASAP7_75t_L g980 ( 
.A(n_959),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_908),
.A2(n_56),
.B(n_57),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_846),
.A2(n_785),
.B(n_782),
.C(n_883),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_845),
.Y(n_983)
);

INVx6_ASAP7_75t_L g984 ( 
.A(n_877),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_783),
.B(n_812),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_845),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_866),
.A2(n_932),
.B(n_813),
.C(n_801),
.Y(n_987)
);

BUFx6f_ASAP7_75t_SL g988 ( 
.A(n_921),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_795),
.B(n_950),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_951),
.A2(n_875),
.B(n_780),
.C(n_954),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_957),
.A2(n_937),
.B(n_938),
.C(n_960),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_908),
.A2(n_787),
.B(n_786),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_797),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_855),
.B(n_805),
.Y(n_994)
);

BUFx10_ASAP7_75t_L g995 ( 
.A(n_815),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_892),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_803),
.B(n_809),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_850),
.B(n_807),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_831),
.A2(n_829),
.B(n_810),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_811),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_897),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_893),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_947),
.B(n_833),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_818),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_855),
.B(n_898),
.Y(n_1005)
);

BUFx12f_ASAP7_75t_L g1006 ( 
.A(n_921),
.Y(n_1006)
);

AND2x6_ASAP7_75t_L g1007 ( 
.A(n_859),
.B(n_927),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_799),
.A2(n_837),
.B1(n_844),
.B2(n_909),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_845),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_855),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_831),
.A2(n_829),
.B(n_793),
.Y(n_1011)
);

O2A1O1Ixp5_ASAP7_75t_SL g1012 ( 
.A1(n_934),
.A2(n_943),
.B(n_920),
.C(n_794),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_887),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_840),
.A2(n_894),
.B1(n_886),
.B2(n_847),
.Y(n_1014)
);

CKINVDCx11_ASAP7_75t_R g1015 ( 
.A(n_827),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_947),
.B(n_863),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_889),
.B(n_800),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_911),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_918),
.B(n_947),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_790),
.A2(n_793),
.B(n_868),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_918),
.B(n_856),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_790),
.A2(n_868),
.B(n_864),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_859),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_SL g1024 ( 
.A(n_804),
.B(n_923),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_913),
.Y(n_1025)
);

BUFx8_ASAP7_75t_L g1026 ( 
.A(n_898),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_798),
.A2(n_857),
.B1(n_878),
.B2(n_796),
.Y(n_1027)
);

O2A1O1Ixp5_ASAP7_75t_L g1028 ( 
.A1(n_861),
.A2(n_839),
.B(n_808),
.C(n_940),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_788),
.B(n_789),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_821),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_888),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_902),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_958),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_940),
.A2(n_882),
.B(n_945),
.C(n_907),
.Y(n_1034)
);

AOI21x1_ASAP7_75t_L g1035 ( 
.A1(n_822),
.A2(n_823),
.B(n_905),
.Y(n_1035)
);

OAI21xp33_ASAP7_75t_SL g1036 ( 
.A1(n_867),
.A2(n_834),
.B(n_835),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_956),
.A2(n_931),
.B(n_917),
.C(n_926),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_824),
.B(n_830),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_819),
.A2(n_912),
.B(n_882),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_961),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_849),
.A2(n_823),
.B(n_781),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_SL g1042 ( 
.A(n_962),
.B(n_948),
.C(n_946),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_961),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_895),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_SL g1045 ( 
.A(n_946),
.B(n_953),
.C(n_944),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_851),
.A2(n_885),
.B1(n_791),
.B2(n_836),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_859),
.B(n_927),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_849),
.A2(n_872),
.B(n_876),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_935),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_802),
.A2(n_806),
.B1(n_817),
.B2(n_843),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_826),
.B(n_838),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_958),
.B(n_871),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_927),
.Y(n_1053)
);

BUFx10_ASAP7_75t_L g1054 ( 
.A(n_955),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_945),
.A2(n_905),
.B(n_873),
.C(n_814),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_816),
.B(n_879),
.Y(n_1056)
);

O2A1O1Ixp5_ASAP7_75t_L g1057 ( 
.A1(n_915),
.A2(n_862),
.B(n_854),
.C(n_914),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_880),
.B(n_910),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_870),
.A2(n_904),
.B1(n_900),
.B2(n_848),
.Y(n_1059)
);

OR2x6_ASAP7_75t_SL g1060 ( 
.A(n_928),
.B(n_841),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_853),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_865),
.A2(n_869),
.B1(n_953),
.B2(n_874),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_890),
.B(n_896),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_891),
.A2(n_936),
.B(n_939),
.C(n_884),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_872),
.A2(n_876),
.B(n_924),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_952),
.B(n_929),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_860),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_930),
.A2(n_881),
.B(n_903),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_903),
.A2(n_884),
.B(n_906),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_890),
.B(n_896),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_899),
.B(n_832),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_899),
.B(n_906),
.Y(n_1072)
);

NOR2x1_ASAP7_75t_L g1073 ( 
.A(n_939),
.B(n_933),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_916),
.A2(n_919),
.B(n_922),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_916),
.A2(n_919),
.B(n_922),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_933),
.A2(n_929),
.B1(n_944),
.B2(n_941),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_942),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_925),
.A2(n_656),
.B(n_630),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_925),
.B(n_784),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_842),
.A2(n_784),
.B1(n_846),
.B2(n_828),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_895),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_842),
.A2(n_828),
.B(n_396),
.C(n_406),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_858),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_784),
.B(n_842),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_842),
.A2(n_784),
.B(n_828),
.C(n_846),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_842),
.B(n_852),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_R g1087 ( 
.A(n_842),
.B(n_319),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_797),
.B(n_669),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_784),
.B(n_842),
.Y(n_1089)
);

AO32x2_ASAP7_75t_L g1090 ( 
.A1(n_799),
.A2(n_766),
.A3(n_870),
.B1(n_745),
.B2(n_690),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_877),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_855),
.B(n_673),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_811),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_811),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_842),
.A2(n_784),
.B(n_828),
.C(n_846),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_784),
.B(n_842),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_811),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_784),
.B(n_842),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_877),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_R g1100 ( 
.A(n_842),
.B(n_319),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_949),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_908),
.A2(n_656),
.B(n_630),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_812),
.B(n_728),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_784),
.B(n_842),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_842),
.A2(n_784),
.B1(n_846),
.B2(n_772),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_SL g1106 ( 
.A1(n_1085),
.A2(n_1095),
.B(n_1104),
.C(n_1089),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1048),
.A2(n_987),
.B(n_999),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_983),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_983),
.Y(n_1109)
);

AO31x2_ASAP7_75t_L g1110 ( 
.A1(n_1064),
.A2(n_982),
.A3(n_1055),
.B(n_1022),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_1020),
.A2(n_1011),
.A3(n_1034),
.B(n_1069),
.Y(n_1111)
);

AO21x1_ASAP7_75t_L g1112 ( 
.A1(n_1082),
.A2(n_1089),
.B(n_1084),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_964),
.Y(n_1113)
);

O2A1O1Ixp5_ASAP7_75t_L g1114 ( 
.A1(n_1084),
.A2(n_1104),
.B(n_1096),
.C(n_1098),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1000),
.Y(n_1115)
);

OAI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1096),
.A2(n_1098),
.B1(n_1080),
.B2(n_1024),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1004),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1105),
.A2(n_989),
.B1(n_1016),
.B2(n_998),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_975),
.B(n_1086),
.C(n_979),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1093),
.Y(n_1120)
);

AO21x2_ASAP7_75t_L g1121 ( 
.A1(n_1035),
.A2(n_1039),
.B(n_1065),
.Y(n_1121)
);

AO31x2_ASAP7_75t_L g1122 ( 
.A1(n_1062),
.A2(n_1076),
.A3(n_1071),
.B(n_1008),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_989),
.B(n_1031),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1094),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_1062),
.A2(n_1076),
.A3(n_1071),
.B(n_1008),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1041),
.A2(n_992),
.B(n_1102),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1023),
.Y(n_1127)
);

AOI221x1_ASAP7_75t_L g1128 ( 
.A1(n_979),
.A2(n_976),
.B1(n_1042),
.B2(n_1046),
.C(n_1079),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_1006),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_1010),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1012),
.A2(n_1028),
.B(n_1036),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1097),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_991),
.A2(n_990),
.B(n_1037),
.C(n_1017),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1014),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1032),
.B(n_1016),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_1007),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1074),
.A2(n_1075),
.B(n_1068),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_968),
.A2(n_1059),
.B(n_1072),
.Y(n_1138)
);

BUFx12f_ASAP7_75t_L g1139 ( 
.A(n_1015),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1003),
.B(n_1061),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1058),
.A2(n_1056),
.B(n_1078),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1003),
.A2(n_1073),
.B(n_1070),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_1081),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1063),
.A2(n_1057),
.B(n_1052),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1077),
.A2(n_1059),
.B(n_971),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_SL g1146 ( 
.A1(n_1021),
.A2(n_1019),
.B(n_974),
.C(n_1051),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1014),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1045),
.A2(n_969),
.B(n_1051),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1013),
.B(n_1025),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_SL g1150 ( 
.A1(n_972),
.A2(n_1038),
.B(n_1046),
.C(n_994),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1027),
.A2(n_1092),
.B(n_1029),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_L g1152 ( 
.A(n_997),
.B(n_985),
.C(n_1024),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_970),
.A2(n_1083),
.B1(n_1040),
.B2(n_1030),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1088),
.B(n_993),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_981),
.A2(n_1029),
.A3(n_1049),
.B(n_1067),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_L g1156 ( 
.A(n_980),
.B(n_1103),
.C(n_1043),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1050),
.A2(n_1033),
.B(n_1018),
.Y(n_1157)
);

AOI221x1_ASAP7_75t_L g1158 ( 
.A1(n_1060),
.A2(n_1090),
.B1(n_965),
.B2(n_966),
.C(n_1101),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1047),
.A2(n_1005),
.B(n_1001),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1026),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_996),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_973),
.B(n_978),
.Y(n_1162)
);

OA21x2_ASAP7_75t_L g1163 ( 
.A1(n_977),
.A2(n_1090),
.B(n_1002),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1087),
.B(n_1100),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_965),
.A2(n_966),
.B(n_1009),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_995),
.B(n_988),
.Y(n_1166)
);

AOI21xp33_ASAP7_75t_L g1167 ( 
.A1(n_1090),
.A2(n_980),
.B(n_1010),
.Y(n_1167)
);

AO21x2_ASAP7_75t_L g1168 ( 
.A1(n_1007),
.A2(n_1023),
.B(n_1053),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_988),
.A2(n_995),
.B1(n_1026),
.B2(n_1044),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1053),
.A2(n_986),
.B(n_1009),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1007),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_986),
.A2(n_1009),
.A3(n_1054),
.B(n_984),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_967),
.B(n_1091),
.Y(n_1173)
);

OA21x2_ASAP7_75t_L g1174 ( 
.A1(n_1099),
.A2(n_1028),
.B(n_1022),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1048),
.A2(n_908),
.B(n_656),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1020),
.A2(n_1048),
.B(n_1074),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1048),
.A2(n_908),
.B(n_656),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1048),
.A2(n_908),
.B(n_656),
.Y(n_1178)
);

NOR2xp67_ASAP7_75t_L g1179 ( 
.A(n_1044),
.B(n_728),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1084),
.A2(n_842),
.B1(n_1098),
.B2(n_1096),
.Y(n_1181)
);

AO22x1_ASAP7_75t_L g1182 ( 
.A1(n_975),
.A2(n_842),
.B1(n_731),
.B2(n_803),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1020),
.A2(n_1048),
.B(n_1074),
.Y(n_1183)
);

NOR4xp25_ASAP7_75t_L g1184 ( 
.A(n_1085),
.B(n_1095),
.C(n_828),
.D(n_979),
.Y(n_1184)
);

NOR2x1_ASAP7_75t_SL g1185 ( 
.A(n_1021),
.B(n_630),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1020),
.A2(n_1048),
.B(n_1074),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1020),
.A2(n_1048),
.B(n_1074),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1048),
.A2(n_908),
.B(n_656),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1048),
.A2(n_908),
.B(n_656),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_964),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1084),
.A2(n_842),
.B1(n_1098),
.B2(n_1096),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1085),
.A2(n_842),
.B(n_828),
.C(n_1095),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1020),
.A2(n_1048),
.B(n_1074),
.Y(n_1195)
);

NOR2x1_ASAP7_75t_R g1196 ( 
.A(n_1044),
.B(n_984),
.Y(n_1196)
);

AOI221x1_ASAP7_75t_L g1197 ( 
.A1(n_1085),
.A2(n_842),
.B1(n_1095),
.B2(n_828),
.C(n_979),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1048),
.A2(n_908),
.B(n_656),
.Y(n_1198)
);

INVx3_ASAP7_75t_SL g1199 ( 
.A(n_1081),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1085),
.A2(n_842),
.B(n_828),
.C(n_1095),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1023),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_998),
.B(n_842),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1105),
.A2(n_842),
.B1(n_1089),
.B2(n_1084),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1015),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1020),
.A2(n_1048),
.B(n_1074),
.Y(n_1205)
);

AOI221x1_ASAP7_75t_L g1206 ( 
.A1(n_1085),
.A2(n_842),
.B1(n_1095),
.B2(n_828),
.C(n_979),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1020),
.A2(n_1048),
.B(n_1074),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1048),
.A2(n_908),
.B(n_656),
.Y(n_1208)
);

AOI221x1_ASAP7_75t_L g1209 ( 
.A1(n_1085),
.A2(n_842),
.B1(n_1095),
.B2(n_828),
.C(n_979),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1000),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1006),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1085),
.A2(n_1095),
.A3(n_987),
.B(n_1064),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1015),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1085),
.A2(n_828),
.B(n_1095),
.C(n_842),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1006),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1048),
.A2(n_908),
.B(n_656),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1048),
.A2(n_908),
.B(n_656),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_983),
.Y(n_1220)
);

AOI31xp67_ASAP7_75t_L g1221 ( 
.A1(n_1080),
.A2(n_1066),
.A3(n_784),
.B(n_846),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1020),
.A2(n_1048),
.B(n_1074),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1020),
.A2(n_1048),
.B(n_1074),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1023),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1048),
.A2(n_908),
.B(n_656),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_993),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1000),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1013),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1085),
.A2(n_1095),
.B(n_784),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1084),
.B(n_842),
.Y(n_1232)
);

AO221x2_ASAP7_75t_L g1233 ( 
.A1(n_979),
.A2(n_1084),
.B1(n_1098),
.B2(n_1096),
.C(n_1089),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1000),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1084),
.A2(n_842),
.B1(n_1098),
.B2(n_1096),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1084),
.A2(n_842),
.B1(n_1098),
.B2(n_1096),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1085),
.A2(n_1095),
.B(n_784),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1048),
.A2(n_908),
.B(n_656),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1000),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1136),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1197),
.A2(n_1209),
.B1(n_1206),
.B2(n_1232),
.Y(n_1243)
);

CKINVDCx6p67_ASAP7_75t_R g1244 ( 
.A(n_1139),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1136),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1229),
.Y(n_1246)
);

CKINVDCx11_ASAP7_75t_R g1247 ( 
.A(n_1143),
.Y(n_1247)
);

CKINVDCx16_ASAP7_75t_R g1248 ( 
.A(n_1160),
.Y(n_1248)
);

BUFx2_ASAP7_75t_SL g1249 ( 
.A(n_1179),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1136),
.B(n_1171),
.Y(n_1250)
);

OAI21xp33_ASAP7_75t_L g1251 ( 
.A1(n_1203),
.A2(n_1119),
.B(n_1184),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1115),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1180),
.B(n_1188),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1231),
.A2(n_1237),
.B1(n_1181),
.B2(n_1192),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1231),
.A2(n_1237),
.B1(n_1181),
.B2(n_1192),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1117),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1233),
.A2(n_1152),
.B1(n_1235),
.B2(n_1236),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1108),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1124),
.Y(n_1259)
);

NAND2xp33_ASAP7_75t_SL g1260 ( 
.A(n_1199),
.B(n_1164),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1235),
.A2(n_1236),
.B1(n_1233),
.B2(n_1116),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1180),
.B(n_1188),
.Y(n_1262)
);

BUFx10_ASAP7_75t_L g1263 ( 
.A(n_1204),
.Y(n_1263)
);

CKINVDCx11_ASAP7_75t_R g1264 ( 
.A(n_1211),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1108),
.Y(n_1265)
);

BUFx12f_ASAP7_75t_L g1266 ( 
.A(n_1215),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1118),
.A2(n_1182),
.B1(n_1212),
.B2(n_1239),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1149),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1132),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_SL g1270 ( 
.A1(n_1153),
.A2(n_1194),
.B1(n_1238),
.B2(n_1226),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1210),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1112),
.A2(n_1226),
.B1(n_1238),
.B2(n_1230),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1228),
.Y(n_1273)
);

INVx6_ASAP7_75t_L g1274 ( 
.A(n_1130),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1227),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1234),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1241),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1172),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1214),
.A2(n_1230),
.B1(n_1202),
.B2(n_1138),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1214),
.A2(n_1123),
.B1(n_1200),
.B2(n_1193),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1128),
.A2(n_1123),
.B1(n_1135),
.B2(n_1140),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1138),
.A2(n_1167),
.B1(n_1134),
.B2(n_1147),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1156),
.A2(n_1166),
.B1(n_1184),
.B2(n_1174),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1167),
.A2(n_1135),
.B1(n_1140),
.B2(n_1151),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1161),
.A2(n_1141),
.B1(n_1154),
.B2(n_1216),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1172),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1169),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1162),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1148),
.A2(n_1174),
.B1(n_1131),
.B2(n_1142),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1111),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1133),
.A2(n_1191),
.B1(n_1113),
.B2(n_1159),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1129),
.A2(n_1217),
.B1(n_1173),
.B2(n_1130),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1148),
.A2(n_1131),
.B1(n_1106),
.B2(n_1163),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1221),
.A2(n_1114),
.B1(n_1144),
.B2(n_1145),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1121),
.A2(n_1213),
.B1(n_1157),
.B2(n_1126),
.Y(n_1295)
);

BUFx12f_ASAP7_75t_L g1296 ( 
.A(n_1109),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1127),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_SL g1298 ( 
.A(n_1109),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1168),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1168),
.Y(n_1300)
);

INVx6_ASAP7_75t_L g1301 ( 
.A(n_1109),
.Y(n_1301)
);

INVx3_ASAP7_75t_L g1302 ( 
.A(n_1127),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_1220),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1201),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1224),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1175),
.A2(n_1240),
.B1(n_1225),
.B2(n_1178),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1185),
.A2(n_1213),
.B1(n_1146),
.B2(n_1223),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1213),
.A2(n_1222),
.B1(n_1183),
.B2(n_1186),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1177),
.A2(n_1190),
.B1(n_1219),
.B2(n_1218),
.Y(n_1309)
);

BUFx8_ASAP7_75t_L g1310 ( 
.A(n_1196),
.Y(n_1310)
);

INVx6_ASAP7_75t_L g1311 ( 
.A(n_1170),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1111),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1155),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1176),
.A2(n_1207),
.B1(n_1195),
.B2(n_1205),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1187),
.A2(n_1158),
.B1(n_1110),
.B2(n_1137),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1121),
.A2(n_1165),
.B1(n_1110),
.B2(n_1208),
.Y(n_1316)
);

BUFx4f_ASAP7_75t_L g1317 ( 
.A(n_1150),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1155),
.Y(n_1318)
);

BUFx12f_ASAP7_75t_L g1319 ( 
.A(n_1122),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1122),
.Y(n_1320)
);

BUFx2_ASAP7_75t_SL g1321 ( 
.A(n_1189),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1125),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1198),
.A2(n_842),
.B1(n_1232),
.B2(n_1089),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1232),
.A2(n_842),
.B1(n_1089),
.B2(n_1084),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1229),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1232),
.A2(n_842),
.B1(n_1100),
.B2(n_1087),
.Y(n_1326)
);

INVx2_ASAP7_75t_R g1327 ( 
.A(n_1136),
.Y(n_1327)
);

CKINVDCx11_ASAP7_75t_R g1328 ( 
.A(n_1139),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1136),
.Y(n_1329)
);

CKINVDCx11_ASAP7_75t_R g1330 ( 
.A(n_1139),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1136),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1149),
.B(n_1013),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1232),
.A2(n_842),
.B1(n_1089),
.B2(n_1084),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1107),
.A2(n_1141),
.B(n_1216),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1232),
.A2(n_842),
.B1(n_1089),
.B2(n_1084),
.Y(n_1335)
);

CKINVDCx14_ASAP7_75t_R g1336 ( 
.A(n_1204),
.Y(n_1336)
);

OAI22xp33_ASAP7_75t_R g1337 ( 
.A1(n_1232),
.A2(n_948),
.B1(n_170),
.B2(n_336),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1203),
.B(n_784),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1232),
.A2(n_842),
.B1(n_1089),
.B2(n_1084),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1232),
.A2(n_842),
.B1(n_1089),
.B2(n_1084),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1120),
.Y(n_1341)
);

BUFx12f_ASAP7_75t_L g1342 ( 
.A(n_1139),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1136),
.Y(n_1343)
);

BUFx4f_ASAP7_75t_SL g1344 ( 
.A(n_1139),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1232),
.A2(n_842),
.B1(n_1105),
.B2(n_1080),
.Y(n_1345)
);

INVx6_ASAP7_75t_L g1346 ( 
.A(n_1136),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1120),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1232),
.B(n_1180),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1232),
.A2(n_842),
.B1(n_1089),
.B2(n_1084),
.Y(n_1349)
);

INVx6_ASAP7_75t_L g1350 ( 
.A(n_1136),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1120),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1232),
.A2(n_842),
.B1(n_1105),
.B2(n_1080),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1247),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1334),
.A2(n_1309),
.B(n_1306),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1290),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1252),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1313),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1257),
.B(n_1261),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1261),
.B(n_1254),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1254),
.B(n_1255),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1322),
.B(n_1312),
.Y(n_1361)
);

NAND2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1317),
.B(n_1278),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1317),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1319),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1318),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1278),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1286),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1337),
.A2(n_1345),
.B1(n_1352),
.B2(n_1338),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1328),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1255),
.B(n_1282),
.Y(n_1370)
);

AND2x2_ASAP7_75t_SL g1371 ( 
.A(n_1284),
.B(n_1320),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1275),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1322),
.B(n_1272),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1312),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1272),
.B(n_1276),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1320),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1299),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1291),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1300),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1338),
.A2(n_1251),
.B1(n_1326),
.B2(n_1349),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1256),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1259),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1269),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1271),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1324),
.A2(n_1340),
.B1(n_1333),
.B2(n_1339),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1273),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1348),
.A2(n_1243),
.B1(n_1287),
.B2(n_1280),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1279),
.B(n_1267),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1277),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1246),
.Y(n_1390)
);

INVx3_ASAP7_75t_SL g1391 ( 
.A(n_1298),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1323),
.A2(n_1335),
.B(n_1340),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1325),
.Y(n_1393)
);

CKINVDCx6p67_ASAP7_75t_R g1394 ( 
.A(n_1330),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1268),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1288),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1253),
.B(n_1262),
.Y(n_1397)
);

AO21x1_ASAP7_75t_L g1398 ( 
.A1(n_1243),
.A2(n_1281),
.B(n_1347),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1332),
.B(n_1324),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1279),
.B(n_1284),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1333),
.B(n_1349),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1293),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1341),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1293),
.B(n_1323),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1266),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1335),
.B(n_1339),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1315),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1351),
.B(n_1270),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1321),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1289),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1274),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1289),
.Y(n_1412)
);

NAND3xp33_ASAP7_75t_L g1413 ( 
.A(n_1285),
.B(n_1283),
.C(n_1307),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1295),
.A2(n_1294),
.B(n_1316),
.Y(n_1414)
);

OR2x6_ASAP7_75t_L g1415 ( 
.A(n_1311),
.B(n_1350),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1295),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1281),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1294),
.A2(n_1316),
.B(n_1285),
.Y(n_1418)
);

INVx5_ASAP7_75t_SL g1419 ( 
.A(n_1394),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1375),
.B(n_1308),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1368),
.A2(n_1260),
.B1(n_1292),
.B2(n_1249),
.Y(n_1421)
);

NAND4xp25_ASAP7_75t_L g1422 ( 
.A(n_1368),
.B(n_1380),
.C(n_1399),
.D(n_1392),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1387),
.A2(n_1311),
.B1(n_1344),
.B2(n_1248),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1413),
.A2(n_1242),
.B(n_1331),
.C(n_1329),
.Y(n_1424)
);

AO32x2_ASAP7_75t_L g1425 ( 
.A1(n_1356),
.A2(n_1314),
.A3(n_1327),
.B1(n_1305),
.B2(n_1301),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1381),
.Y(n_1426)
);

NOR2xp67_ASAP7_75t_SL g1427 ( 
.A(n_1378),
.B(n_1342),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1388),
.B(n_1311),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1385),
.A2(n_1297),
.B(n_1304),
.C(n_1250),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1401),
.A2(n_1250),
.B(n_1331),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1381),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1353),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1358),
.A2(n_1329),
.B(n_1245),
.C(n_1343),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1374),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1406),
.A2(n_1302),
.B(n_1303),
.Y(n_1435)
);

NOR2xp67_ASAP7_75t_L g1436 ( 
.A(n_1411),
.B(n_1296),
.Y(n_1436)
);

O2A1O1Ixp33_ASAP7_75t_SL g1437 ( 
.A1(n_1397),
.A2(n_1327),
.B(n_1344),
.C(n_1336),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1408),
.B(n_1258),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1391),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1415),
.B(n_1350),
.Y(n_1440)
);

OR2x6_ASAP7_75t_L g1441 ( 
.A(n_1415),
.B(n_1362),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1415),
.A2(n_1343),
.B(n_1346),
.Y(n_1442)
);

AO21x2_ASAP7_75t_L g1443 ( 
.A1(n_1398),
.A2(n_1343),
.B(n_1301),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1382),
.B(n_1244),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1375),
.B(n_1396),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_SL g1446 ( 
.A1(n_1398),
.A2(n_1336),
.B(n_1310),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1417),
.A2(n_1310),
.B(n_1264),
.C(n_1263),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1414),
.A2(n_1418),
.B(n_1417),
.Y(n_1448)
);

AO32x2_ASAP7_75t_L g1449 ( 
.A1(n_1411),
.A2(n_1265),
.A3(n_1274),
.B1(n_1402),
.B2(n_1412),
.Y(n_1449)
);

AOI211xp5_ASAP7_75t_L g1450 ( 
.A1(n_1388),
.A2(n_1265),
.B(n_1400),
.C(n_1370),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1359),
.A2(n_1360),
.B1(n_1370),
.B2(n_1371),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1390),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1393),
.Y(n_1453)
);

AO32x2_ASAP7_75t_L g1454 ( 
.A1(n_1402),
.A2(n_1410),
.A3(n_1412),
.B1(n_1373),
.B2(n_1361),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1354),
.A2(n_1371),
.B(n_1409),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_SL g1456 ( 
.A(n_1409),
.B(n_1364),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1403),
.B(n_1372),
.Y(n_1457)
);

OR2x6_ASAP7_75t_L g1458 ( 
.A(n_1362),
.B(n_1364),
.Y(n_1458)
);

NOR2x1_ASAP7_75t_SL g1459 ( 
.A(n_1364),
.B(n_1366),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1382),
.B(n_1383),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1360),
.B(n_1359),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1371),
.A2(n_1391),
.B1(n_1395),
.B2(n_1404),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_SL g1463 ( 
.A(n_1441),
.B(n_1367),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1448),
.B(n_1425),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1460),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_SL g1466 ( 
.A1(n_1451),
.A2(n_1404),
.B1(n_1410),
.B2(n_1407),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1426),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1434),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1431),
.Y(n_1469)
);

NOR2xp67_ASAP7_75t_L g1470 ( 
.A(n_1455),
.B(n_1384),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1441),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1434),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1445),
.B(n_1416),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1422),
.A2(n_1423),
.B1(n_1451),
.B2(n_1462),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1452),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1425),
.B(n_1449),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1428),
.B(n_1386),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1462),
.A2(n_1363),
.B1(n_1364),
.B2(n_1362),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1449),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1457),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1454),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1454),
.B(n_1376),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1454),
.B(n_1418),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1420),
.B(n_1355),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1441),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1461),
.B(n_1377),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1453),
.B(n_1361),
.Y(n_1487)
);

INVx4_ASAP7_75t_L g1488 ( 
.A(n_1471),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1471),
.A2(n_1423),
.B1(n_1421),
.B2(n_1440),
.Y(n_1489)
);

OAI33xp33_ASAP7_75t_L g1490 ( 
.A1(n_1486),
.A2(n_1389),
.A3(n_1444),
.B1(n_1447),
.B2(n_1365),
.B3(n_1357),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1474),
.B(n_1450),
.C(n_1427),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1480),
.B(n_1438),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1467),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1487),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1463),
.B(n_1458),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1463),
.B(n_1458),
.Y(n_1496)
);

OAI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1474),
.A2(n_1435),
.B1(n_1447),
.B2(n_1428),
.C(n_1424),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1467),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1487),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1482),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1465),
.B(n_1482),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1468),
.Y(n_1502)
);

OR2x6_ASAP7_75t_L g1503 ( 
.A(n_1471),
.B(n_1442),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1468),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1472),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1472),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1473),
.B(n_1374),
.Y(n_1507)
);

INVx4_ASAP7_75t_L g1508 ( 
.A(n_1471),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1463),
.B(n_1456),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1484),
.B(n_1367),
.Y(n_1510)
);

OR2x6_ASAP7_75t_L g1511 ( 
.A(n_1485),
.B(n_1440),
.Y(n_1511)
);

OAI211xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1475),
.A2(n_1435),
.B(n_1430),
.C(n_1429),
.Y(n_1512)
);

INVxp67_ASAP7_75t_L g1513 ( 
.A(n_1487),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1487),
.Y(n_1514)
);

OAI21xp33_ASAP7_75t_L g1515 ( 
.A1(n_1466),
.A2(n_1476),
.B(n_1483),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1484),
.B(n_1367),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1469),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1473),
.B(n_1379),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1509),
.B(n_1478),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1509),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1500),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1513),
.B(n_1505),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1491),
.B(n_1475),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1491),
.B(n_1439),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1498),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1493),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1497),
.A2(n_1466),
.B1(n_1446),
.B2(n_1478),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1501),
.B(n_1464),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1493),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1494),
.B(n_1479),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1495),
.B(n_1470),
.Y(n_1531)
);

NOR2x1_ASAP7_75t_L g1532 ( 
.A(n_1509),
.B(n_1443),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1494),
.B(n_1479),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1506),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1493),
.Y(n_1535)
);

OR2x6_ASAP7_75t_L g1536 ( 
.A(n_1511),
.B(n_1470),
.Y(n_1536)
);

INVxp67_ASAP7_75t_SL g1537 ( 
.A(n_1504),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1507),
.B(n_1481),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1506),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1510),
.B(n_1464),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1517),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1510),
.B(n_1464),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1516),
.B(n_1464),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1516),
.B(n_1479),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1517),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1545),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1522),
.B(n_1507),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1545),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1524),
.B(n_1394),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1520),
.B(n_1509),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1524),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1545),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1523),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_1523),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1520),
.B(n_1540),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1541),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1520),
.B(n_1495),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1526),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1534),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1527),
.A2(n_1515),
.B(n_1489),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1522),
.B(n_1518),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1541),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1520),
.B(n_1495),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1540),
.B(n_1542),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1541),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1537),
.B(n_1518),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1534),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1537),
.B(n_1499),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1541),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1540),
.B(n_1495),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1539),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1527),
.B(n_1515),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1526),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1539),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1538),
.B(n_1514),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1525),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1532),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1519),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1519),
.Y(n_1579)
);

NOR2x1_ASAP7_75t_L g1580 ( 
.A(n_1532),
.B(n_1488),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1526),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1538),
.B(n_1481),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1540),
.B(n_1477),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1544),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1542),
.B(n_1477),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1531),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1525),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1525),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1561),
.B(n_1538),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1564),
.B(n_1542),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1564),
.B(n_1542),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1546),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1553),
.B(n_1554),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1559),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1549),
.B(n_1369),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1546),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1551),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1555),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1579),
.B(n_1492),
.Y(n_1599)
);

OAI21xp33_ASAP7_75t_L g1600 ( 
.A1(n_1572),
.A2(n_1512),
.B(n_1532),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1548),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1578),
.B(n_1492),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1548),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1560),
.A2(n_1490),
.B1(n_1496),
.B2(n_1503),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1552),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1555),
.B(n_1543),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1583),
.B(n_1543),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1552),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1557),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1570),
.B(n_1543),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1557),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1571),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1561),
.B(n_1521),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1547),
.B(n_1521),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1576),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1563),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1570),
.B(n_1543),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1550),
.B(n_1544),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1574),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1547),
.B(n_1521),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1550),
.B(n_1544),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1585),
.B(n_1544),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1563),
.B(n_1528),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1576),
.Y(n_1624)
);

OA21x2_ASAP7_75t_L g1625 ( 
.A1(n_1600),
.A2(n_1577),
.B(n_1619),
.Y(n_1625)
);

AOI211xp5_ASAP7_75t_L g1626 ( 
.A1(n_1593),
.A2(n_1567),
.B(n_1577),
.C(n_1586),
.Y(n_1626)
);

OAI32xp33_ASAP7_75t_L g1627 ( 
.A1(n_1597),
.A2(n_1574),
.A3(n_1568),
.B1(n_1584),
.B2(n_1566),
.Y(n_1627)
);

AOI32xp33_ASAP7_75t_L g1628 ( 
.A1(n_1609),
.A2(n_1580),
.A3(n_1531),
.B1(n_1508),
.B2(n_1488),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1592),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1594),
.B(n_1566),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1592),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1595),
.A2(n_1568),
.B(n_1432),
.Y(n_1632)
);

OAI33xp33_ASAP7_75t_L g1633 ( 
.A1(n_1612),
.A2(n_1587),
.A3(n_1588),
.B1(n_1569),
.B2(n_1556),
.B3(n_1565),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1596),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1596),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1604),
.A2(n_1437),
.B(n_1405),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1616),
.B(n_1575),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1611),
.B(n_1531),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1611),
.B(n_1531),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1601),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1601),
.Y(n_1641)
);

NAND2x1_ASAP7_75t_L g1642 ( 
.A(n_1598),
.B(n_1531),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1599),
.B(n_1575),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1598),
.B(n_1531),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1623),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1603),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1602),
.A2(n_1536),
.B(n_1503),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1622),
.A2(n_1536),
.B(n_1587),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1603),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1627),
.A2(n_1625),
.B(n_1626),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1632),
.B(n_1630),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1637),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1645),
.B(n_1610),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1625),
.A2(n_1623),
.B1(n_1536),
.B2(n_1496),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1643),
.B(n_1607),
.Y(n_1655)
);

AOI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1627),
.A2(n_1624),
.B1(n_1605),
.B2(n_1615),
.C(n_1608),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1625),
.B(n_1608),
.C(n_1605),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1638),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1645),
.B(n_1610),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1629),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1631),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1628),
.B(n_1419),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1649),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1634),
.B(n_1589),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1636),
.A2(n_1648),
.B1(n_1647),
.B2(n_1642),
.C(n_1639),
.Y(n_1665)
);

AOI322xp5_ASAP7_75t_L g1666 ( 
.A1(n_1635),
.A2(n_1606),
.A3(n_1591),
.B1(n_1590),
.B2(n_1621),
.C1(n_1618),
.C2(n_1617),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1640),
.B(n_1617),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1641),
.Y(n_1668)
);

A2O1A1Ixp33_ASAP7_75t_L g1669 ( 
.A1(n_1650),
.A2(n_1642),
.B(n_1646),
.C(n_1639),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1663),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1663),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1652),
.B(n_1615),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1658),
.B(n_1638),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1651),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1659),
.B(n_1589),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1667),
.B(n_1590),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1664),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1665),
.B(n_1419),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1678),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1673),
.Y(n_1680)
);

OAI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1669),
.A2(n_1662),
.B1(n_1654),
.B2(n_1656),
.C(n_1655),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1670),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1671),
.B(n_1653),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1672),
.Y(n_1684)
);

NOR3xp33_ASAP7_75t_L g1685 ( 
.A(n_1674),
.B(n_1677),
.C(n_1672),
.Y(n_1685)
);

NAND4xp25_ASAP7_75t_L g1686 ( 
.A(n_1675),
.B(n_1676),
.C(n_1660),
.D(n_1661),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1670),
.Y(n_1687)
);

AOI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1681),
.A2(n_1685),
.B1(n_1682),
.B2(n_1684),
.C(n_1686),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1683),
.Y(n_1689)
);

OAI221xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1680),
.A2(n_1666),
.B1(n_1657),
.B2(n_1668),
.C(n_1644),
.Y(n_1690)
);

OAI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1679),
.A2(n_1687),
.B1(n_1668),
.B2(n_1624),
.C(n_1644),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1682),
.Y(n_1692)
);

O2A1O1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1690),
.A2(n_1633),
.B(n_1614),
.C(n_1620),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1688),
.A2(n_1606),
.B1(n_1621),
.B2(n_1618),
.C(n_1591),
.Y(n_1694)
);

AOI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1692),
.A2(n_1620),
.B1(n_1614),
.B2(n_1613),
.C(n_1556),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_L g1696 ( 
.A(n_1689),
.B(n_1419),
.Y(n_1696)
);

O2A1O1Ixp5_ASAP7_75t_SL g1697 ( 
.A1(n_1691),
.A2(n_1588),
.B(n_1562),
.C(n_1565),
.Y(n_1697)
);

A2O1A1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1688),
.A2(n_1613),
.B(n_1558),
.C(n_1581),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1698),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1696),
.Y(n_1700)
);

NOR2x1_ASAP7_75t_L g1701 ( 
.A(n_1693),
.B(n_1697),
.Y(n_1701)
);

XNOR2x1_ASAP7_75t_L g1702 ( 
.A(n_1694),
.B(n_1503),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_SL g1703 ( 
.A(n_1695),
.B(n_1391),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1703),
.A2(n_1581),
.B1(n_1573),
.B2(n_1558),
.Y(n_1704)
);

OR4x1_ASAP7_75t_L g1705 ( 
.A(n_1699),
.B(n_1562),
.C(n_1505),
.D(n_1502),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1700),
.B(n_1530),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1706),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_1707),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_SL g1709 ( 
.A(n_1708),
.B(n_1704),
.C(n_1701),
.Y(n_1709)
);

NAND4xp25_ASAP7_75t_L g1710 ( 
.A(n_1708),
.B(n_1705),
.C(n_1702),
.D(n_1436),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1709),
.A2(n_1573),
.B1(n_1582),
.B2(n_1521),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1710),
.A2(n_1582),
.B1(n_1529),
.B2(n_1526),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1711),
.A2(n_1712),
.B1(n_1488),
.B2(n_1508),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1711),
.A2(n_1535),
.B(n_1529),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_SL g1715 ( 
.A1(n_1714),
.A2(n_1433),
.B(n_1459),
.Y(n_1715)
);

OAI21xp33_ASAP7_75t_L g1716 ( 
.A1(n_1715),
.A2(n_1713),
.B(n_1533),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1716),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1717),
.A2(n_1535),
.B1(n_1529),
.B2(n_1530),
.C(n_1533),
.Y(n_1718)
);

AOI211xp5_ASAP7_75t_L g1719 ( 
.A1(n_1718),
.A2(n_1363),
.B(n_1530),
.C(n_1533),
.Y(n_1719)
);


endmodule