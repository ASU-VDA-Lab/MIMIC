module fake_aes_2402_n_47 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_47);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_47;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_SL g10 ( .A(n_3), .B(n_8), .Y(n_10) );
BUFx6f_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
INVx1_ASAP7_75t_SL g12 ( .A(n_4), .Y(n_12) );
AND3x2_ASAP7_75t_L g13 ( .A(n_0), .B(n_1), .C(n_7), .Y(n_13) );
NOR2xp33_ASAP7_75t_R g14 ( .A(n_1), .B(n_4), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_5), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_9), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_15), .B(n_2), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_17), .B(n_7), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_18), .B(n_5), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_11), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_16), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_11), .Y(n_24) );
BUFx6f_ASAP7_75t_L g25 ( .A(n_11), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_16), .Y(n_26) );
OAI221xp5_ASAP7_75t_L g27 ( .A1(n_19), .A2(n_12), .B1(n_10), .B2(n_11), .C(n_13), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_24), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_24), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_23), .Y(n_30) );
AOI221xp5_ASAP7_75t_SL g31 ( .A1(n_26), .A2(n_11), .B1(n_10), .B2(n_14), .C(n_6), .Y(n_31) );
AOI221xp5_ASAP7_75t_L g32 ( .A1(n_27), .A2(n_20), .B1(n_21), .B2(n_22), .C(n_25), .Y(n_32) );
INVx2_ASAP7_75t_SL g33 ( .A(n_30), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_28), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
NAND2xp5_ASAP7_75t_L g36 ( .A(n_33), .B(n_31), .Y(n_36) );
AND2x2_ASAP7_75t_L g37 ( .A(n_34), .B(n_6), .Y(n_37) );
INVx8_ASAP7_75t_L g38 ( .A(n_37), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
NOR4xp25_ASAP7_75t_SL g40 ( .A(n_35), .B(n_32), .C(n_28), .D(n_29), .Y(n_40) );
NOR2x1_ASAP7_75t_L g41 ( .A(n_39), .B(n_35), .Y(n_41) );
AOI22xp5_ASAP7_75t_L g42 ( .A1(n_38), .A2(n_36), .B1(n_29), .B2(n_25), .Y(n_42) );
O2A1O1Ixp33_ASAP7_75t_L g43 ( .A1(n_38), .A2(n_22), .B(n_25), .C(n_40), .Y(n_43) );
INVx1_ASAP7_75t_L g44 ( .A(n_41), .Y(n_44) );
INVx1_ASAP7_75t_L g45 ( .A(n_43), .Y(n_45) );
OAI221xp5_ASAP7_75t_L g46 ( .A1(n_44), .A2(n_42), .B1(n_25), .B2(n_22), .C(n_38), .Y(n_46) );
AOI22xp5_ASAP7_75t_L g47 ( .A1(n_46), .A2(n_45), .B1(n_44), .B2(n_22), .Y(n_47) );
endmodule