module fake_jpeg_6714_n_70 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_70);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_70;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_4),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_18),
.B(n_3),
.C(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_6),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_9),
.B(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_13),
.Y(n_30)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_20),
.Y(n_41)
);

CKINVDCx12_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_12),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_21),
.A2(n_15),
.B1(n_17),
.B2(n_11),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_17),
.B1(n_16),
.B2(n_19),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_44),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_47),
.B1(n_45),
.B2(n_41),
.Y(n_54)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_23),
.C(n_22),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_38),
.C(n_35),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_46),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_29),
.A2(n_19),
.B1(n_22),
.B2(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_31),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_33),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_52),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_53),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_54),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_48),
.B(n_49),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_56),
.B(n_60),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_51),
.B(n_33),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_53),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_64),
.A2(n_57),
.B1(n_43),
.B2(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_43),
.Y(n_68)
);

FAx1_ASAP7_75t_SL g67 ( 
.A(n_65),
.B(n_44),
.CI(n_57),
.CON(n_67),
.SN(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_67),
.B(n_68),
.Y(n_70)
);


endmodule