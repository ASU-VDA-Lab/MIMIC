module fake_ariane_652_n_2109 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2109);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2109;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_279;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_261;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_2075;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_180),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_13),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_56),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_64),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_61),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_63),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_115),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_111),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_198),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_151),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_201),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_152),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_45),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_103),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_173),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_118),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_19),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_23),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_86),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_184),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_124),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_187),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_142),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_123),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_26),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_98),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_20),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_85),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_33),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_29),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_106),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_15),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_164),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_83),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_42),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_143),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_147),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_57),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_100),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_60),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_7),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_88),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_75),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_73),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_4),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_203),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_89),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_52),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_91),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_53),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_126),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_70),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_19),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_25),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_40),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_114),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_53),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_13),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_80),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_165),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_0),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_153),
.Y(n_275)
);

BUFx8_ASAP7_75t_SL g276 ( 
.A(n_137),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_52),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_75),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_205),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_76),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_42),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_44),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_25),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_182),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_176),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_80),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_167),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_33),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_150),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_6),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_127),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_15),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_135),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_8),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_73),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_62),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_64),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_83),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_4),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_138),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_160),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_2),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_102),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_81),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_7),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_129),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_121),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_69),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_189),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_26),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_163),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_172),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_141),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_122),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_9),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_97),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_3),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_31),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_131),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_8),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_40),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_162),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_94),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_69),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_74),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_178),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_63),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_113),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_10),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_46),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_65),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_41),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_76),
.Y(n_333)
);

BUFx2_ASAP7_75t_SL g334 ( 
.A(n_130),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_3),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_31),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_38),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_125),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_62),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_66),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_55),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_6),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_21),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_57),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_72),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_23),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_104),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_14),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_132),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_37),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_192),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_27),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_183),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_144),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_95),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_54),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_36),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_56),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_108),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_177),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_48),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_28),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_202),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_190),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_84),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_204),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_82),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_107),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_134),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_199),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_90),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_28),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_5),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_87),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_24),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_197),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_179),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_38),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_9),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_55),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_168),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_140),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_1),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_16),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_50),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_21),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_48),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_105),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_154),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_193),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_1),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_81),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_18),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_34),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_27),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_169),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_51),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_35),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_11),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_0),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_2),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_59),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_18),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_51),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_72),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_357),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_237),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_209),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_224),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_258),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_319),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_208),
.B(n_5),
.Y(n_412)
);

NOR2x1_ASAP7_75t_L g413 ( 
.A(n_237),
.B(n_92),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_354),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_209),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_357),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_400),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_276),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_208),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_331),
.Y(n_420)
);

INVxp33_ASAP7_75t_SL g421 ( 
.A(n_400),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_274),
.B(n_10),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_223),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_223),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_331),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_211),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_263),
.B(n_11),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_227),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_227),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_212),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_281),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_229),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_237),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_222),
.Y(n_434)
);

INVxp33_ASAP7_75t_SL g435 ( 
.A(n_213),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_214),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_215),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_229),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_281),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_226),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_230),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_222),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_246),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_230),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_240),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_232),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_232),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_239),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_239),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_263),
.B(n_12),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_249),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_249),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_243),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_250),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_251),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_247),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_251),
.Y(n_457)
);

INVxp33_ASAP7_75t_SL g458 ( 
.A(n_253),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_274),
.B(n_12),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_228),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_371),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_247),
.Y(n_462)
);

BUFx6f_ASAP7_75t_SL g463 ( 
.A(n_269),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_271),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_273),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_260),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_281),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_273),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_300),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_262),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_300),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_307),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_307),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_277),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_375),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_296),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_265),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_267),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_228),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_299),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_313),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_238),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_356),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_268),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_313),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_322),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_270),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_238),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_322),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_323),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_365),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_272),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_278),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_323),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_280),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_359),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_282),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_326),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_359),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_283),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_326),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_351),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_341),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_351),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_286),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_355),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_288),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g508 ( 
.A(n_274),
.B(n_14),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_355),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_292),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_371),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_375),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_360),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_269),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_360),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_269),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_375),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_463),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_408),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_408),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_431),
.B(n_363),
.Y(n_522)
);

AND2x4_ASAP7_75t_SL g523 ( 
.A(n_514),
.B(n_341),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_418),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_407),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_423),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_433),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_433),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_420),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_421),
.A2(n_320),
.B1(n_329),
.B2(n_236),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_423),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_424),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_439),
.B(n_363),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_424),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_428),
.B(n_379),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_428),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_429),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_429),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_432),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_432),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_438),
.B(n_368),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_438),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_441),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_441),
.B(n_379),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_444),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_444),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_446),
.B(n_368),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_409),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_511),
.A2(n_320),
.B1(n_329),
.B2(n_236),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_446),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_456),
.B(n_207),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_447),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_447),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_448),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g557 ( 
.A(n_456),
.B(n_225),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_512),
.B(n_379),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_448),
.B(n_369),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_449),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_449),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_451),
.B(n_452),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_451),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_410),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_452),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_455),
.B(n_266),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_455),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_425),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_457),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_503),
.B(n_406),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_457),
.B(n_304),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_465),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_465),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_468),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_468),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_469),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_469),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_413),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_471),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_471),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_472),
.Y(n_581)
);

CKINVDCx11_ASAP7_75t_R g582 ( 
.A(n_445),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_472),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_473),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_412),
.B(n_207),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_473),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_481),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_481),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_485),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_485),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_486),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_486),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_489),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_489),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_490),
.Y(n_595)
);

AND3x2_ASAP7_75t_L g596 ( 
.A(n_416),
.B(n_302),
.C(n_266),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_490),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_494),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_494),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_498),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_498),
.B(n_369),
.Y(n_601)
);

OA21x2_ASAP7_75t_L g602 ( 
.A1(n_501),
.A2(n_390),
.B(n_370),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_501),
.Y(n_603)
);

OA21x2_ASAP7_75t_L g604 ( 
.A1(n_502),
.A2(n_390),
.B(n_370),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_539),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_539),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_539),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_539),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_520),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_557),
.B(n_426),
.Y(n_610)
);

AND3x2_ASAP7_75t_L g611 ( 
.A(n_557),
.B(n_427),
.C(n_417),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_539),
.B(n_347),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_518),
.Y(n_613)
);

CKINVDCx6p67_ASAP7_75t_R g614 ( 
.A(n_582),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_539),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_531),
.B(n_430),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_539),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_539),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_518),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_520),
.Y(n_620)
);

AND3x2_ASAP7_75t_L g621 ( 
.A(n_531),
.B(n_568),
.C(n_466),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_524),
.B(n_496),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_550),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_566),
.B(n_467),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_540),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_517),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_564),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_540),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_L g629 ( 
.A(n_540),
.B(n_347),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_540),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_540),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_541),
.B(n_462),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_540),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_585),
.A2(n_461),
.B1(n_419),
.B2(n_450),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_517),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_522),
.Y(n_636)
);

AND2x4_ASAP7_75t_SL g637 ( 
.A(n_518),
.B(n_499),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_520),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_526),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_531),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_541),
.B(n_475),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_526),
.Y(n_642)
);

INVxp33_ASAP7_75t_SL g643 ( 
.A(n_568),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_522),
.B(n_440),
.C(n_436),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_544),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_585),
.A2(n_461),
.B1(n_419),
.B2(n_508),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_541),
.B(n_503),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_544),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_544),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_568),
.B(n_443),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_535),
.Y(n_651)
);

OR2x6_ASAP7_75t_L g652 ( 
.A(n_553),
.B(n_508),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_553),
.A2(n_435),
.B1(n_458),
.B2(n_454),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_544),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_520),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_535),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_529),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_570),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_532),
.A2(n_459),
.B1(n_422),
.B2(n_434),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_519),
.Y(n_660)
);

INVxp33_ASAP7_75t_L g661 ( 
.A(n_570),
.Y(n_661)
);

NOR2x1p5_ASAP7_75t_L g662 ( 
.A(n_517),
.B(n_470),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_SL g663 ( 
.A(n_532),
.B(n_478),
.C(n_477),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_529),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_526),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_519),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_529),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_544),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_566),
.B(n_502),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_558),
.B(n_484),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_541),
.B(n_504),
.Y(n_671)
);

AND2x2_ASAP7_75t_SL g672 ( 
.A(n_518),
.B(n_266),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_558),
.B(n_487),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_544),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_566),
.B(n_562),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_558),
.B(n_492),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_529),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_541),
.B(n_552),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_544),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_526),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_544),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_547),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_SL g683 ( 
.A(n_518),
.B(n_493),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_547),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_571),
.B(n_495),
.Y(n_685)
);

CKINVDCx16_ASAP7_75t_R g686 ( 
.A(n_551),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_547),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_571),
.A2(n_500),
.B1(n_505),
.B2(n_497),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_551),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_552),
.B(n_504),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_547),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_562),
.B(n_506),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_547),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_547),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_552),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_547),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_552),
.B(n_506),
.Y(n_697)
);

BUFx10_ASAP7_75t_L g698 ( 
.A(n_571),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_571),
.A2(n_510),
.B1(n_507),
.B2(n_516),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_547),
.Y(n_700)
);

BUFx10_ASAP7_75t_L g701 ( 
.A(n_571),
.Y(n_701)
);

OR2x6_ASAP7_75t_L g702 ( 
.A(n_543),
.B(n_442),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_SL g703 ( 
.A(n_521),
.B(n_437),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_552),
.B(n_509),
.Y(n_704)
);

BUFx4f_ASAP7_75t_L g705 ( 
.A(n_602),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_548),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_548),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_548),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_548),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_548),
.Y(n_710)
);

BUFx4f_ASAP7_75t_L g711 ( 
.A(n_602),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_548),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_521),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_548),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_561),
.B(n_509),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_548),
.Y(n_716)
);

AND2x6_ASAP7_75t_L g717 ( 
.A(n_533),
.B(n_413),
.Y(n_717)
);

INVx6_ASAP7_75t_L g718 ( 
.A(n_578),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_523),
.B(n_460),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_561),
.B(n_513),
.Y(n_720)
);

INVx6_ASAP7_75t_L g721 ( 
.A(n_578),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_561),
.B(n_575),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_602),
.A2(n_513),
.B1(n_515),
.B2(n_463),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_555),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_555),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_555),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_555),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_555),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_555),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_555),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_561),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_602),
.A2(n_515),
.B1(n_463),
.B2(n_304),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_596),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_555),
.B(n_347),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_577),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_582),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_561),
.B(n_341),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_537),
.A2(n_405),
.B1(n_333),
.B2(n_479),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_577),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_602),
.A2(n_304),
.B1(n_394),
.B2(n_330),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_575),
.B(n_225),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_525),
.B(n_527),
.Y(n_742)
);

BUFx4f_ASAP7_75t_L g743 ( 
.A(n_602),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_575),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_577),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_525),
.B(n_527),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_575),
.B(n_235),
.Y(n_747)
);

NOR2x1p5_ASAP7_75t_L g748 ( 
.A(n_543),
.B(n_241),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_575),
.B(n_235),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_528),
.B(n_482),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_549),
.B(n_488),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_577),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_523),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_577),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_604),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_692),
.B(n_595),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_705),
.B(n_578),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_652),
.A2(n_578),
.B1(n_604),
.B2(n_523),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_660),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_705),
.B(n_578),
.Y(n_760)
);

OR2x6_ASAP7_75t_L g761 ( 
.A(n_652),
.B(n_537),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_609),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_692),
.B(n_595),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_666),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_609),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_675),
.B(n_595),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_705),
.B(n_578),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_675),
.B(n_595),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_669),
.B(n_595),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_669),
.B(n_528),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_750),
.B(n_542),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_620),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_698),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_647),
.B(n_542),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_711),
.B(n_578),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_713),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_698),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_640),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_624),
.B(n_545),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_620),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_695),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_626),
.A2(n_554),
.B(n_556),
.C(n_545),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_673),
.Y(n_783)
);

O2A1O1Ixp5_ASAP7_75t_L g784 ( 
.A1(n_704),
.A2(n_554),
.B(n_560),
.C(n_556),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_698),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_695),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_744),
.Y(n_787)
);

AND2x6_ASAP7_75t_L g788 ( 
.A(n_744),
.B(n_537),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_678),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_736),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_624),
.B(n_523),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_626),
.B(n_560),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_722),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_731),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_623),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_755),
.B(n_577),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_671),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_701),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_627),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_663),
.B(n_405),
.C(n_333),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_652),
.A2(n_689),
.B1(n_740),
.B2(n_659),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_635),
.B(n_563),
.Y(n_802)
);

NAND3xp33_ASAP7_75t_L g803 ( 
.A(n_676),
.B(n_565),
.C(n_563),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_635),
.B(n_565),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_702),
.B(n_537),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_690),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_652),
.A2(n_578),
.B1(n_604),
.B2(n_537),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_641),
.B(n_572),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_697),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_636),
.B(n_572),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_636),
.B(n_573),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_638),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_622),
.Y(n_813)
);

NAND2x1p5_ASAP7_75t_L g814 ( 
.A(n_672),
.B(n_604),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_638),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_719),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_711),
.B(n_577),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_689),
.A2(n_604),
.B1(n_546),
.B2(n_574),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_655),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_636),
.B(n_573),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_661),
.B(n_411),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_715),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_702),
.A2(n_751),
.B1(n_651),
.B2(n_656),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_702),
.A2(n_581),
.B1(n_583),
.B2(n_574),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_655),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_742),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_701),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_746),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_720),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_651),
.B(n_581),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_651),
.B(n_583),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_657),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_656),
.B(n_586),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_657),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_702),
.A2(n_546),
.B1(n_588),
.B2(n_586),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_643),
.B(n_414),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_658),
.B(n_546),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_632),
.A2(n_559),
.B(n_549),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_719),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_711),
.B(n_577),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_664),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_SL g842 ( 
.A(n_643),
.B(n_453),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_656),
.B(n_588),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_751),
.B(n_590),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_701),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_664),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_751),
.B(n_546),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_699),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_667),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_743),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_751),
.B(n_590),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_748),
.B(n_591),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_672),
.B(n_591),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_731),
.B(n_597),
.Y(n_854)
);

AND2x4_ASAP7_75t_SL g855 ( 
.A(n_614),
.B(n_464),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_731),
.B(n_597),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_703),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_741),
.B(n_599),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_743),
.B(n_587),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_743),
.B(n_587),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_733),
.B(n_599),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_639),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_667),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_677),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_639),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_677),
.Y(n_866)
);

NOR3xp33_ASAP7_75t_L g867 ( 
.A(n_616),
.B(n_245),
.C(n_241),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_747),
.B(n_749),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_646),
.B(n_600),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_717),
.A2(n_604),
.B1(n_600),
.B2(n_603),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_679),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_639),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_755),
.A2(n_533),
.B(n_536),
.C(n_534),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_706),
.B(n_587),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_644),
.B(n_474),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_706),
.B(n_587),
.Y(n_876)
);

INVx8_ASAP7_75t_L g877 ( 
.A(n_717),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_706),
.B(n_587),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_634),
.B(n_603),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_642),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_642),
.Y(n_881)
);

OAI22xp33_ASAP7_75t_L g882 ( 
.A1(n_653),
.A2(n_738),
.B1(n_688),
.B2(n_686),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_706),
.B(n_587),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_723),
.B(n_538),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_665),
.B(n_538),
.Y(n_885)
);

INVxp33_ASAP7_75t_L g886 ( 
.A(n_670),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_665),
.B(n_611),
.Y(n_887)
);

INVx8_ASAP7_75t_L g888 ( 
.A(n_717),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_732),
.B(n_538),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_650),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_754),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_639),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_639),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_737),
.B(n_685),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_610),
.A2(n_567),
.B1(n_576),
.B2(n_569),
.Y(n_895)
);

OAI22xp33_ASAP7_75t_L g896 ( 
.A1(n_733),
.A2(n_559),
.B1(n_601),
.B2(n_394),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_753),
.B(n_476),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_662),
.A2(n_601),
.B1(n_533),
.B2(n_536),
.Y(n_898)
);

OAI221xp5_ASAP7_75t_L g899 ( 
.A1(n_683),
.A2(n_394),
.B1(n_252),
.B2(n_255),
.C(n_256),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_637),
.B(n_480),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_754),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_717),
.B(n_567),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_680),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_717),
.B(n_567),
.Y(n_904)
);

NOR3xp33_ASAP7_75t_L g905 ( 
.A(n_736),
.B(n_252),
.C(n_245),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_752),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_752),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_717),
.B(n_569),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_706),
.B(n_587),
.Y(n_909)
);

NAND3xp33_ASAP7_75t_L g910 ( 
.A(n_621),
.B(n_589),
.C(n_587),
.Y(n_910)
);

INVx5_ASAP7_75t_L g911 ( 
.A(n_718),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_680),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_613),
.B(n_589),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_680),
.B(n_569),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_680),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_679),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_682),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_613),
.B(n_589),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_680),
.B(n_576),
.Y(n_919)
);

OAI221xp5_ASAP7_75t_L g920 ( 
.A1(n_612),
.A2(n_308),
.B1(n_297),
.B2(n_255),
.C(n_310),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_682),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_605),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_615),
.B(n_579),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_605),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_615),
.B(n_579),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_850),
.B(n_613),
.Y(n_926)
);

INVx4_ASAP7_75t_L g927 ( 
.A(n_877),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_861),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_759),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_826),
.A2(n_534),
.B(n_536),
.C(n_533),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_783),
.B(n_637),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_796),
.A2(n_619),
.B(n_607),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_873),
.A2(n_607),
.B(n_606),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_873),
.A2(n_608),
.B(n_606),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_828),
.B(n_579),
.Y(n_935)
);

OAI21xp33_ASAP7_75t_L g936 ( 
.A1(n_810),
.A2(n_295),
.B(n_294),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_796),
.A2(n_619),
.B(n_617),
.Y(n_937)
);

AOI21x1_ASAP7_75t_L g938 ( 
.A1(n_913),
.A2(n_617),
.B(n_608),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_771),
.B(n_779),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_756),
.A2(n_763),
.B(n_853),
.C(n_838),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_778),
.B(n_483),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_850),
.B(n_619),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_766),
.A2(n_536),
.B(n_594),
.C(n_534),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_853),
.A2(n_594),
.B(n_534),
.C(n_584),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_868),
.A2(n_625),
.B(n_618),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_811),
.B(n_580),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_764),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_794),
.B(n_630),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_839),
.B(n_491),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_776),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_795),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_820),
.B(n_580),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_877),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_791),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_817),
.A2(n_625),
.B(n_618),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_817),
.A2(n_631),
.B(n_628),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_877),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_794),
.B(n_630),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_770),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_813),
.B(n_530),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_830),
.B(n_580),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_769),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_848),
.B(n_630),
.Y(n_963)
);

AO21x1_ASAP7_75t_L g964 ( 
.A1(n_840),
.A2(n_629),
.B(n_612),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_842),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_762),
.Y(n_966)
);

AO21x1_ASAP7_75t_L g967 ( 
.A1(n_859),
.A2(n_734),
.B(n_629),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_791),
.B(n_816),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_792),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_877),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_860),
.A2(n_856),
.B(n_854),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_831),
.B(n_584),
.Y(n_972)
);

OAI321xp33_ASAP7_75t_L g973 ( 
.A1(n_882),
.A2(n_308),
.A3(n_344),
.B1(n_343),
.B2(n_342),
.C(n_391),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_768),
.A2(n_823),
.B1(n_843),
.B2(n_833),
.Y(n_974)
);

NOR2x1_ASAP7_75t_R g975 ( 
.A(n_790),
.B(n_298),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_861),
.B(n_584),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_791),
.B(n_596),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_794),
.B(n_649),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_L g979 ( 
.A(n_836),
.B(n_257),
.C(n_256),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_773),
.B(n_649),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_773),
.B(n_649),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_861),
.B(n_592),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_801),
.B(n_592),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_774),
.A2(n_594),
.B(n_592),
.C(n_257),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_852),
.B(n_594),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_852),
.B(n_589),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_799),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_821),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_777),
.B(n_654),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_923),
.A2(n_645),
.B(n_633),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_765),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_925),
.A2(n_918),
.B(n_913),
.Y(n_992)
);

NAND2x1p5_ASAP7_75t_L g993 ( 
.A(n_911),
.B(n_530),
.Y(n_993)
);

OAI22xp33_ASAP7_75t_L g994 ( 
.A1(n_835),
.A2(n_305),
.B1(n_317),
.B2(n_315),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_851),
.B(n_589),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_851),
.B(n_589),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_851),
.B(n_589),
.Y(n_997)
);

AOI21xp33_ASAP7_75t_L g998 ( 
.A1(n_886),
.A2(n_668),
.B(n_648),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_918),
.A2(n_668),
.B(n_648),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_897),
.B(n_530),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_858),
.A2(n_681),
.B(n_674),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_911),
.B(n_530),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_777),
.B(n_654),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_808),
.A2(n_681),
.B(n_674),
.Y(n_1004)
);

BUFx12f_ASAP7_75t_L g1005 ( 
.A(n_790),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_855),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_844),
.B(n_589),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_797),
.B(n_593),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_806),
.B(n_593),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_837),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_900),
.B(n_530),
.Y(n_1011)
);

AOI21xp33_ASAP7_75t_L g1012 ( 
.A1(n_886),
.A2(n_691),
.B(n_684),
.Y(n_1012)
);

BUFx4f_ASAP7_75t_L g1013 ( 
.A(n_855),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_785),
.B(n_654),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_824),
.A2(n_290),
.B(n_310),
.C(n_297),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_802),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_804),
.A2(n_290),
.B(n_321),
.C(n_318),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_834),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_875),
.B(n_341),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_814),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_809),
.B(n_593),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_890),
.B(n_593),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_765),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_782),
.A2(n_330),
.B(n_361),
.C(n_302),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_L g1025 ( 
.A(n_888),
.B(n_684),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_788),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_849),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_822),
.B(n_593),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_789),
.A2(n_321),
.B(n_325),
.C(n_318),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_772),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_793),
.B(n_593),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_785),
.A2(n_745),
.B1(n_714),
.B2(n_691),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_914),
.A2(n_694),
.B(n_693),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_879),
.B(n_593),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_798),
.A2(n_745),
.B1(n_714),
.B2(n_693),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_863),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_784),
.A2(n_700),
.B(n_694),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_896),
.B(n_805),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_805),
.B(n_593),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_847),
.B(n_598),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_902),
.A2(n_707),
.B(n_700),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_888),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_L g1043 ( 
.A(n_800),
.B(n_857),
.C(n_803),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_894),
.B(n_714),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_919),
.A2(n_876),
.B(n_874),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_874),
.A2(n_710),
.B(n_707),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_876),
.A2(n_724),
.B(n_710),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_772),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_888),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_798),
.B(n_745),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_847),
.B(n_598),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_758),
.B(n_598),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_870),
.A2(n_696),
.B(n_687),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_818),
.B(n_598),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_807),
.A2(n_761),
.B1(n_888),
.B2(n_869),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_827),
.A2(n_739),
.B1(n_735),
.B2(n_730),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_788),
.B(n_598),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_780),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_866),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_827),
.B(n_687),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_878),
.A2(n_725),
.B(n_724),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_780),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_788),
.B(n_598),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_878),
.A2(n_909),
.B(n_883),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_898),
.A2(n_373),
.B(n_325),
.C(n_327),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_867),
.B(n_598),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_883),
.A2(n_726),
.B(n_725),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_899),
.A2(n_373),
.B(n_327),
.C(n_332),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_L g1069 ( 
.A(n_905),
.B(n_342),
.C(n_332),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_845),
.A2(n_814),
.B1(n_781),
.B2(n_787),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_788),
.B(n_598),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_L g1072 ( 
.A1(n_904),
.A2(n_727),
.B(n_726),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_812),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_909),
.A2(n_728),
.B(n_727),
.Y(n_1074)
);

NOR2xp67_ASAP7_75t_L g1075 ( 
.A(n_910),
.B(n_696),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_895),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_812),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_815),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_908),
.A2(n_730),
.B(n_728),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_815),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_757),
.A2(n_739),
.B(n_735),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_757),
.A2(n_709),
.B(n_708),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_760),
.A2(n_709),
.B(n_708),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_760),
.A2(n_716),
.B(n_712),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_767),
.A2(n_716),
.B(n_712),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_L g1086 ( 
.A(n_887),
.B(n_729),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_788),
.B(n_845),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_767),
.A2(n_729),
.B(n_734),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_788),
.B(n_718),
.Y(n_1089)
);

CKINVDCx14_ASAP7_75t_R g1090 ( 
.A(n_761),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_761),
.A2(n_242),
.B1(n_718),
.B2(n_721),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_761),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_829),
.B(n_718),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_775),
.A2(n_242),
.B(n_217),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_922),
.A2(n_396),
.B(n_216),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_786),
.A2(n_343),
.B(n_393),
.C(n_391),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_880),
.B(n_721),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_911),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_920),
.A2(n_383),
.B(n_367),
.C(n_344),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_924),
.A2(n_330),
.B(n_361),
.C(n_403),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_881),
.B(n_721),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_775),
.A2(n_218),
.B(n_210),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_871),
.A2(n_396),
.B(n_216),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_885),
.A2(n_220),
.B(n_219),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_871),
.A2(n_231),
.B(n_221),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_872),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_872),
.B(n_207),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_819),
.B(n_721),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_892),
.B(n_324),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_893),
.A2(n_383),
.B(n_393),
.C(n_302),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_903),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_987),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_939),
.A2(n_865),
.B1(n_862),
.B2(n_912),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_959),
.A2(n_865),
.B1(n_862),
.B2(n_912),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_1005),
.Y(n_1115)
);

OR2x6_ASAP7_75t_L g1116 ( 
.A(n_928),
.B(n_872),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_979),
.A2(n_403),
.B(n_361),
.C(n_862),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_988),
.B(n_872),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1005),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1013),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_968),
.B(n_865),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_932),
.A2(n_915),
.B(n_901),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_928),
.B(n_911),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_R g1124 ( 
.A(n_1013),
.B(n_915),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1106),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_1026),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_954),
.B(n_911),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_1106),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1106),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_937),
.A2(n_915),
.B(n_921),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_969),
.B(n_825),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_949),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_SL g1133 ( 
.A1(n_931),
.A2(n_943),
.B(n_984),
.C(n_1109),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_951),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_931),
.B(n_915),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_SL g1136 ( 
.A1(n_965),
.A2(n_345),
.B1(n_404),
.B2(n_362),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1016),
.B(n_825),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_971),
.A2(n_940),
.B(n_1045),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_968),
.B(n_832),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_962),
.B(n_1019),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_974),
.A2(n_921),
.B1(n_917),
.B2(n_916),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_940),
.A2(n_917),
.B(n_901),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_929),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_947),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_963),
.B(n_1010),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_945),
.A2(n_992),
.B(n_1004),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_994),
.A2(n_403),
.B(n_907),
.C(n_906),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_941),
.B(n_891),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1043),
.B(n_891),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1069),
.A2(n_916),
.B(n_907),
.C(n_906),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_963),
.B(n_832),
.Y(n_1151)
);

AO32x1_ASAP7_75t_L g1152 ( 
.A1(n_1070),
.A2(n_864),
.A3(n_846),
.B1(n_841),
.B2(n_275),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_SL g1153 ( 
.A(n_1068),
.B(n_336),
.C(n_335),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1000),
.B(n_841),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1006),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1026),
.A2(n_889),
.B1(n_884),
.B2(n_864),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_955),
.A2(n_846),
.B(n_275),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_957),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_950),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_977),
.B(n_337),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1011),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_973),
.B(n_339),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1106),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_1092),
.B(n_334),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1065),
.A2(n_311),
.B(n_275),
.C(n_309),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_956),
.A2(n_309),
.B(n_216),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1038),
.B(n_340),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_976),
.B(n_346),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1015),
.A2(n_311),
.B(n_309),
.C(n_314),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_982),
.B(n_348),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1099),
.A2(n_314),
.B(n_311),
.C(n_334),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1018),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1055),
.A2(n_402),
.B1(n_401),
.B2(n_380),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_985),
.B(n_350),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1027),
.Y(n_1175)
);

AOI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1072),
.A2(n_314),
.B(n_311),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_936),
.A2(n_352),
.B(n_358),
.C(n_372),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_957),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_957),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_SL g1180 ( 
.A(n_975),
.B(n_233),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_983),
.B(n_378),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1055),
.A2(n_399),
.B1(n_398),
.B2(n_397),
.Y(n_1182)
);

INVxp67_ASAP7_75t_L g1183 ( 
.A(n_1109),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1036),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_935),
.B(n_384),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1087),
.B(n_385),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1022),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_946),
.B(n_952),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1091),
.B(n_386),
.Y(n_1189)
);

BUFx4_ASAP7_75t_SL g1190 ( 
.A(n_1111),
.Y(n_1190)
);

BUFx4f_ASAP7_75t_L g1191 ( 
.A(n_957),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1059),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_995),
.A2(n_395),
.B1(n_392),
.B2(n_387),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1044),
.A2(n_944),
.B(n_986),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1095),
.A2(n_1044),
.B(n_1029),
.C(n_1017),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_927),
.B(n_970),
.Y(n_1196)
);

AO32x1_ASAP7_75t_L g1197 ( 
.A1(n_1032),
.A2(n_16),
.A3(n_17),
.B1(n_20),
.B2(n_22),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_996),
.A2(n_389),
.B1(n_388),
.B2(n_382),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1090),
.B(n_234),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1024),
.A2(n_1096),
.B(n_930),
.C(n_944),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1090),
.A2(n_1020),
.B1(n_1078),
.B2(n_1077),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1024),
.A2(n_17),
.B(n_22),
.C(n_24),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1041),
.A2(n_381),
.B(n_377),
.C(n_376),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_927),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_961),
.B(n_29),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1081),
.A2(n_374),
.B(n_366),
.Y(n_1206)
);

NOR2xp67_ASAP7_75t_SL g1207 ( 
.A(n_1098),
.B(n_244),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1001),
.A2(n_364),
.B(n_353),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_997),
.Y(n_1209)
);

NOR3xp33_ASAP7_75t_SL g1210 ( 
.A(n_930),
.B(n_349),
.C(n_338),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1039),
.B(n_248),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1040),
.B(n_254),
.Y(n_1212)
);

NOR2xp67_ASAP7_75t_L g1213 ( 
.A(n_1098),
.B(n_93),
.Y(n_1213)
);

OAI21xp33_ASAP7_75t_SL g1214 ( 
.A1(n_1103),
.A2(n_30),
.B(n_32),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_966),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_927),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1053),
.A2(n_128),
.B(n_206),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1051),
.B(n_259),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_972),
.B(n_30),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1079),
.A2(n_328),
.B(n_316),
.C(n_312),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_993),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_991),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_960),
.B(n_32),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1008),
.A2(n_306),
.B1(n_303),
.B2(n_301),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_991),
.B(n_1023),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1064),
.A2(n_293),
.B(n_291),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_993),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1110),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1088),
.A2(n_289),
.B(n_287),
.Y(n_1229)
);

AND2x6_ASAP7_75t_L g1230 ( 
.A(n_1049),
.B(n_953),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1066),
.A2(n_285),
.B1(n_284),
.B2(n_279),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1023),
.B(n_37),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_970),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_998),
.A2(n_1012),
.B(n_1076),
.C(n_1063),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_990),
.A2(n_1085),
.B(n_1084),
.Y(n_1235)
);

O2A1O1Ixp5_ASAP7_75t_L g1236 ( 
.A1(n_964),
.A2(n_39),
.B(n_41),
.C(n_43),
.Y(n_1236)
);

BUFx4f_ASAP7_75t_L g1237 ( 
.A(n_1002),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1082),
.A2(n_264),
.B(n_261),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1030),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1002),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_970),
.B(n_39),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1048),
.B(n_43),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1048),
.B(n_44),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1058),
.B(n_45),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1053),
.A2(n_112),
.B(n_194),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1042),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1042),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1058),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1083),
.A2(n_110),
.B(n_188),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1042),
.B(n_46),
.Y(n_1250)
);

BUFx8_ASAP7_75t_L g1251 ( 
.A(n_1062),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1031),
.A2(n_109),
.B(n_186),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_953),
.B(n_47),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1062),
.B(n_47),
.Y(n_1254)
);

BUFx2_ASAP7_75t_SL g1255 ( 
.A(n_1086),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1009),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1073),
.B(n_58),
.Y(n_1257)
);

NAND2xp33_ASAP7_75t_SL g1258 ( 
.A(n_1049),
.B(n_58),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1057),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1025),
.A2(n_133),
.B(n_185),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1049),
.B(n_65),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1025),
.A2(n_136),
.B(n_181),
.Y(n_1262)
);

OAI21xp33_ASAP7_75t_SL g1263 ( 
.A1(n_933),
.A2(n_934),
.B(n_1021),
.Y(n_1263)
);

O2A1O1Ixp5_ASAP7_75t_L g1264 ( 
.A1(n_967),
.A2(n_67),
.B(n_68),
.C(n_70),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1073),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1089),
.B(n_67),
.Y(n_1266)
);

OAI222xp33_ASAP7_75t_L g1267 ( 
.A1(n_1052),
.A2(n_68),
.B1(n_71),
.B2(n_74),
.C1(n_77),
.C2(n_78),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1080),
.Y(n_1268)
);

AO32x2_ASAP7_75t_L g1269 ( 
.A1(n_1141),
.A2(n_1035),
.A3(n_1056),
.B1(n_1100),
.B2(n_938),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1156),
.A2(n_1100),
.A3(n_1034),
.B(n_1054),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1145),
.B(n_1080),
.Y(n_1271)
);

XOR2xp5_ASAP7_75t_L g1272 ( 
.A(n_1115),
.B(n_1094),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1138),
.A2(n_926),
.B(n_942),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1146),
.A2(n_926),
.B(n_942),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1183),
.B(n_1007),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1143),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1263),
.A2(n_1028),
.B(n_1071),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1263),
.A2(n_948),
.B(n_978),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1188),
.A2(n_948),
.B(n_978),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_1119),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1132),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1134),
.Y(n_1282)
);

CKINVDCx14_ASAP7_75t_R g1283 ( 
.A(n_1120),
.Y(n_1283)
);

NAND2xp33_ASAP7_75t_SL g1284 ( 
.A(n_1124),
.B(n_989),
.Y(n_1284)
);

NAND3xp33_ASAP7_75t_L g1285 ( 
.A(n_1195),
.B(n_981),
.C(n_1014),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1235),
.A2(n_958),
.B(n_1033),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1173),
.A2(n_1075),
.B1(n_980),
.B2(n_981),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1122),
.A2(n_958),
.B(n_1060),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1217),
.A2(n_1061),
.B(n_1074),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1191),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1148),
.B(n_1140),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1123),
.B(n_980),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1130),
.A2(n_1060),
.B(n_999),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1194),
.A2(n_1067),
.B(n_1046),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1142),
.A2(n_1037),
.B(n_1107),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1245),
.A2(n_1047),
.B(n_1107),
.Y(n_1296)
);

NAND3x1_ASAP7_75t_L g1297 ( 
.A(n_1173),
.B(n_1102),
.C(n_1101),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1123),
.B(n_989),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_SL g1299 ( 
.A1(n_1200),
.A2(n_1097),
.B(n_1105),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1161),
.B(n_1050),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1151),
.A2(n_1050),
.B(n_1014),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1211),
.A2(n_1104),
.B(n_1003),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1144),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1251),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1112),
.B(n_1003),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1133),
.A2(n_1108),
.B(n_1093),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1234),
.A2(n_145),
.A3(n_175),
.B(n_174),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1113),
.A2(n_139),
.B(n_171),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1160),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1121),
.B(n_78),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1176),
.A2(n_146),
.B(n_166),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1159),
.B(n_79),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1214),
.A2(n_82),
.B(n_84),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1155),
.Y(n_1314)
);

AO21x1_ASAP7_75t_L g1315 ( 
.A1(n_1149),
.A2(n_96),
.B(n_99),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1251),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1214),
.A2(n_101),
.B(n_116),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1260),
.A2(n_117),
.B(n_120),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1116),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1199),
.B(n_196),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1191),
.Y(n_1321)
);

AO32x2_ASAP7_75t_L g1322 ( 
.A1(n_1256),
.A2(n_149),
.A3(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1116),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1262),
.A2(n_159),
.B(n_161),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_SL g1325 ( 
.A1(n_1203),
.A2(n_1220),
.B(n_1250),
.C(n_1241),
.Y(n_1325)
);

AO32x2_ASAP7_75t_L g1326 ( 
.A1(n_1114),
.A2(n_1187),
.A3(n_1182),
.B1(n_1209),
.B2(n_1193),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1172),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1139),
.B(n_1175),
.Y(n_1328)
);

AO21x1_ASAP7_75t_L g1329 ( 
.A1(n_1226),
.A2(n_1258),
.B(n_1205),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1116),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1267),
.A2(n_1167),
.B(n_1153),
.C(n_1259),
.Y(n_1331)
);

BUFx12f_ASAP7_75t_L g1332 ( 
.A(n_1164),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1219),
.A2(n_1252),
.B(n_1237),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1157),
.A2(n_1249),
.B(n_1166),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1237),
.A2(n_1135),
.B(n_1196),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1184),
.B(n_1192),
.Y(n_1336)
);

OR2x6_ASAP7_75t_L g1337 ( 
.A(n_1126),
.B(n_1127),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1127),
.B(n_1126),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1239),
.A2(n_1268),
.A3(n_1265),
.B(n_1248),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1196),
.A2(n_1229),
.B(n_1154),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1150),
.A2(n_1225),
.B(n_1244),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1174),
.B(n_1162),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1168),
.B(n_1170),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1164),
.Y(n_1344)
);

NOR2xp67_ASAP7_75t_SL g1345 ( 
.A(n_1247),
.B(n_1216),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1232),
.A2(n_1242),
.B(n_1243),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1212),
.A2(n_1218),
.B(n_1171),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1215),
.A2(n_1222),
.A3(n_1257),
.B(n_1254),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1131),
.A2(n_1137),
.B(n_1186),
.Y(n_1349)
);

AO32x2_ASAP7_75t_L g1350 ( 
.A1(n_1231),
.A2(n_1136),
.A3(n_1197),
.B1(n_1152),
.B2(n_1224),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1236),
.A2(n_1264),
.B(n_1246),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1164),
.B(n_1180),
.Y(n_1352)
);

CKINVDCx6p67_ASAP7_75t_R g1353 ( 
.A(n_1247),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1204),
.A2(n_1233),
.B(n_1246),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1204),
.A2(n_1233),
.B(n_1216),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1147),
.A2(n_1152),
.B(n_1261),
.Y(n_1356)
);

NOR2xp67_ASAP7_75t_L g1357 ( 
.A(n_1247),
.B(n_1158),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1190),
.Y(n_1358)
);

AO21x1_ASAP7_75t_L g1359 ( 
.A1(n_1202),
.A2(n_1118),
.B(n_1223),
.Y(n_1359)
);

INVx5_ASAP7_75t_L g1360 ( 
.A(n_1125),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1253),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1253),
.B(n_1185),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1152),
.A2(n_1261),
.B(n_1266),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1181),
.B(n_1201),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1189),
.A2(n_1210),
.B1(n_1117),
.B2(n_1228),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1213),
.A2(n_1238),
.B(n_1165),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1125),
.Y(n_1367)
);

NAND3xp33_ASAP7_75t_SL g1368 ( 
.A(n_1177),
.B(n_1169),
.C(n_1208),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1125),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1221),
.A2(n_1227),
.B1(n_1240),
.B2(n_1178),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1255),
.B(n_1128),
.Y(n_1371)
);

NAND3xp33_ASAP7_75t_L g1372 ( 
.A(n_1207),
.B(n_1198),
.C(n_1206),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1213),
.A2(n_1230),
.B(n_1178),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1128),
.Y(n_1374)
);

AO32x2_ASAP7_75t_L g1375 ( 
.A1(n_1197),
.A2(n_1158),
.A3(n_1129),
.B1(n_1128),
.B2(n_1163),
.Y(n_1375)
);

NAND2x1p5_ASAP7_75t_L g1376 ( 
.A(n_1179),
.B(n_1221),
.Y(n_1376)
);

AO21x1_ASAP7_75t_L g1377 ( 
.A1(n_1197),
.A2(n_1221),
.B(n_1227),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1129),
.A2(n_1163),
.B(n_1227),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1179),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1179),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1240),
.A2(n_796),
.B(n_1138),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1230),
.A2(n_940),
.B(n_1263),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1230),
.B(n_1132),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1230),
.B(n_1132),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1138),
.A2(n_796),
.B(n_1146),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1138),
.A2(n_796),
.B(n_1146),
.Y(n_1386)
);

AND2x2_ASAP7_75t_SL g1387 ( 
.A(n_1173),
.B(n_1013),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1138),
.A2(n_796),
.B(n_1146),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1145),
.B(n_783),
.Y(n_1389)
);

INVx6_ASAP7_75t_L g1390 ( 
.A(n_1251),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1138),
.A2(n_1235),
.B(n_1146),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1263),
.A2(n_940),
.B(n_1194),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1138),
.A2(n_796),
.B(n_1146),
.Y(n_1393)
);

NAND2x1p5_ASAP7_75t_L g1394 ( 
.A(n_1134),
.B(n_1013),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1132),
.B(n_1112),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1138),
.A2(n_1235),
.B(n_1146),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1138),
.A2(n_1146),
.B(n_1235),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1138),
.A2(n_1235),
.B(n_1146),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1143),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1115),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1138),
.A2(n_796),
.B(n_1146),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1143),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1263),
.A2(n_940),
.B(n_1194),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1123),
.B(n_928),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_SL g1405 ( 
.A1(n_1133),
.A2(n_940),
.B(n_939),
.C(n_1195),
.Y(n_1405)
);

CKINVDCx11_ASAP7_75t_R g1406 ( 
.A(n_1134),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1183),
.A2(n_783),
.B(n_1195),
.C(n_1173),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1138),
.A2(n_1235),
.B(n_1146),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1263),
.A2(n_940),
.B(n_1194),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1183),
.B(n_823),
.Y(n_1410)
);

NOR2x1_ASAP7_75t_R g1411 ( 
.A(n_1120),
.B(n_736),
.Y(n_1411)
);

NOR2xp67_ASAP7_75t_L g1412 ( 
.A(n_1247),
.B(n_1158),
.Y(n_1412)
);

AO21x1_ASAP7_75t_L g1413 ( 
.A1(n_1149),
.A2(n_974),
.B(n_1070),
.Y(n_1413)
);

AO31x2_ASAP7_75t_L g1414 ( 
.A1(n_1156),
.A2(n_1141),
.A3(n_1142),
.B(n_1234),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1112),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1115),
.Y(n_1416)
);

AOI31xp67_ASAP7_75t_L g1417 ( 
.A1(n_1151),
.A2(n_1107),
.A3(n_1060),
.B(n_1135),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1112),
.Y(n_1418)
);

OAI22x1_ASAP7_75t_L g1419 ( 
.A1(n_1173),
.A2(n_551),
.B1(n_836),
.B2(n_1183),
.Y(n_1419)
);

OA21x2_ASAP7_75t_L g1420 ( 
.A1(n_1138),
.A2(n_1146),
.B(n_1235),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1115),
.Y(n_1421)
);

AO31x2_ASAP7_75t_L g1422 ( 
.A1(n_1156),
.A2(n_1141),
.A3(n_1142),
.B(n_1234),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1162),
.A2(n_689),
.B1(n_557),
.B2(n_897),
.Y(n_1423)
);

AOI21x1_ASAP7_75t_SL g1424 ( 
.A1(n_1205),
.A2(n_811),
.B(n_810),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1263),
.A2(n_940),
.B(n_1194),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1138),
.A2(n_796),
.B(n_1146),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1134),
.Y(n_1427)
);

OR2x6_ASAP7_75t_L g1428 ( 
.A(n_1123),
.B(n_928),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1138),
.A2(n_796),
.B(n_1146),
.Y(n_1429)
);

AO31x2_ASAP7_75t_L g1430 ( 
.A1(n_1156),
.A2(n_1141),
.A3(n_1142),
.B(n_1234),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1143),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1138),
.A2(n_796),
.B(n_1146),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1183),
.A2(n_783),
.B(n_1195),
.C(n_1173),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1138),
.A2(n_1235),
.B(n_1146),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1407),
.A2(n_1433),
.B1(n_1310),
.B2(n_1423),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_SL g1436 ( 
.A1(n_1387),
.A2(n_1313),
.B1(n_1317),
.B2(n_1342),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1419),
.A2(n_1362),
.B1(n_1410),
.B2(n_1389),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1313),
.A2(n_1317),
.B1(n_1364),
.B2(n_1309),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1336),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1321),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1397),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1406),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1352),
.A2(n_1347),
.B1(n_1332),
.B2(n_1309),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1291),
.A2(n_1343),
.B1(n_1425),
.B2(n_1392),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1395),
.B(n_1281),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1304),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1379),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1282),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1276),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1321),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1303),
.Y(n_1451)
);

CKINVDCx20_ASAP7_75t_R g1452 ( 
.A(n_1316),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1327),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1328),
.B(n_1275),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1340),
.A2(n_1331),
.B(n_1285),
.Y(n_1455)
);

OAI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1392),
.A2(n_1409),
.B1(n_1425),
.B2(n_1403),
.Y(n_1456)
);

CKINVDCx11_ASAP7_75t_R g1457 ( 
.A(n_1280),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1399),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1390),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1403),
.A2(n_1409),
.B1(n_1329),
.B2(n_1413),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1402),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1382),
.A2(n_1365),
.B1(n_1361),
.B2(n_1287),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1320),
.A2(n_1382),
.B1(n_1344),
.B2(n_1377),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1380),
.Y(n_1464)
);

CKINVDCx11_ASAP7_75t_R g1465 ( 
.A(n_1421),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1359),
.A2(n_1272),
.B1(n_1368),
.B2(n_1292),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1431),
.A2(n_1312),
.B1(n_1271),
.B2(n_1315),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1383),
.A2(n_1384),
.B1(n_1287),
.B2(n_1305),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1390),
.A2(n_1372),
.B1(n_1285),
.B2(n_1302),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1415),
.B(n_1418),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1292),
.A2(n_1427),
.B1(n_1404),
.B2(n_1428),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1339),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1404),
.A2(n_1428),
.B1(n_1284),
.B2(n_1300),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1339),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1385),
.A2(n_1401),
.B(n_1432),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1339),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1338),
.A2(n_1428),
.B1(n_1358),
.B2(n_1394),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1337),
.Y(n_1478)
);

BUFx12f_ASAP7_75t_L g1479 ( 
.A(n_1400),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1372),
.A2(n_1349),
.B1(n_1323),
.B2(n_1338),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1358),
.A2(n_1337),
.B1(n_1314),
.B2(n_1298),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1297),
.A2(n_1290),
.B1(n_1283),
.B2(n_1337),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1319),
.B(n_1369),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1322),
.A2(n_1363),
.B1(n_1330),
.B2(n_1356),
.Y(n_1484)
);

CKINVDCx11_ASAP7_75t_R g1485 ( 
.A(n_1353),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1416),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1367),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1330),
.A2(n_1279),
.B1(n_1278),
.B2(n_1299),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1295),
.A2(n_1301),
.B1(n_1346),
.B2(n_1277),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1290),
.A2(n_1306),
.B1(n_1370),
.B2(n_1374),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1348),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1333),
.A2(n_1335),
.B1(n_1294),
.B2(n_1388),
.Y(n_1492)
);

AOI21xp33_ASAP7_75t_L g1493 ( 
.A1(n_1371),
.A2(n_1373),
.B(n_1341),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1386),
.A2(n_1429),
.B(n_1426),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1325),
.A2(n_1405),
.B1(n_1357),
.B2(n_1412),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1322),
.A2(n_1324),
.B1(n_1318),
.B2(n_1366),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1393),
.A2(n_1273),
.B1(n_1355),
.B2(n_1381),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1295),
.A2(n_1322),
.B1(n_1308),
.B2(n_1326),
.Y(n_1498)
);

OR2x6_ASAP7_75t_L g1499 ( 
.A(n_1378),
.B(n_1376),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1326),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1354),
.A2(n_1274),
.B1(n_1357),
.B2(n_1412),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1360),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1360),
.Y(n_1503)
);

BUFx10_ASAP7_75t_L g1504 ( 
.A(n_1411),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1326),
.A2(n_1350),
.B1(n_1288),
.B2(n_1351),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1345),
.A2(n_1360),
.B1(n_1411),
.B2(n_1311),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1397),
.Y(n_1507)
);

INVx8_ASAP7_75t_L g1508 ( 
.A(n_1424),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1414),
.B(n_1422),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1350),
.A2(n_1420),
.B1(n_1286),
.B2(n_1375),
.Y(n_1510)
);

OAI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1375),
.A2(n_1350),
.B1(n_1293),
.B2(n_1420),
.Y(n_1511)
);

OAI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1375),
.A2(n_1307),
.B1(n_1269),
.B2(n_1417),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1270),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1269),
.A2(n_1307),
.B1(n_1430),
.B2(n_1422),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1414),
.B(n_1430),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1414),
.B(n_1430),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1270),
.Y(n_1517)
);

BUFx4f_ASAP7_75t_SL g1518 ( 
.A(n_1269),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1334),
.A2(n_1396),
.B1(n_1408),
.B2(n_1398),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1391),
.A2(n_1434),
.B1(n_1296),
.B2(n_1289),
.Y(n_1520)
);

INVx3_ASAP7_75t_SL g1521 ( 
.A(n_1270),
.Y(n_1521)
);

CKINVDCx11_ASAP7_75t_R g1522 ( 
.A(n_1422),
.Y(n_1522)
);

BUFx4f_ASAP7_75t_SL g1523 ( 
.A(n_1280),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1336),
.Y(n_1524)
);

INVx6_ASAP7_75t_L g1525 ( 
.A(n_1321),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1313),
.A2(n_1173),
.B1(n_973),
.B2(n_1419),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1313),
.A2(n_1173),
.B1(n_973),
.B2(n_1419),
.Y(n_1527)
);

BUFx8_ASAP7_75t_L g1528 ( 
.A(n_1280),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1321),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_689),
.B2(n_652),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1280),
.Y(n_1531)
);

BUFx12f_ASAP7_75t_L g1532 ( 
.A(n_1406),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_689),
.B2(n_652),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_SL g1534 ( 
.A1(n_1387),
.A2(n_557),
.B1(n_410),
.B2(n_411),
.Y(n_1534)
);

BUFx4f_ASAP7_75t_SL g1535 ( 
.A(n_1280),
.Y(n_1535)
);

INVx6_ASAP7_75t_L g1536 ( 
.A(n_1321),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1406),
.Y(n_1537)
);

BUFx12f_ASAP7_75t_L g1538 ( 
.A(n_1406),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1390),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1291),
.B(n_1389),
.Y(n_1540)
);

CKINVDCx6p67_ASAP7_75t_R g1541 ( 
.A(n_1406),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_689),
.B2(n_652),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1390),
.Y(n_1543)
);

OAI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1342),
.A2(n_557),
.B1(n_686),
.B2(n_1173),
.Y(n_1544)
);

BUFx4f_ASAP7_75t_SL g1545 ( 
.A(n_1280),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1336),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1336),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1280),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1406),
.Y(n_1549)
);

CKINVDCx20_ASAP7_75t_R g1550 ( 
.A(n_1406),
.Y(n_1550)
);

INVx6_ASAP7_75t_L g1551 ( 
.A(n_1321),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1336),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_689),
.B2(n_652),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_689),
.B2(n_652),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1428),
.B(n_1338),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1387),
.A2(n_557),
.B1(n_410),
.B2(n_411),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1406),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1406),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1347),
.A2(n_783),
.B(n_1407),
.Y(n_1559)
);

BUFx8_ASAP7_75t_L g1560 ( 
.A(n_1280),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1321),
.Y(n_1561)
);

BUFx2_ASAP7_75t_SL g1562 ( 
.A(n_1304),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1406),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1379),
.Y(n_1564)
);

CKINVDCx14_ASAP7_75t_R g1565 ( 
.A(n_1283),
.Y(n_1565)
);

BUFx8_ASAP7_75t_SL g1566 ( 
.A(n_1280),
.Y(n_1566)
);

BUFx12f_ASAP7_75t_L g1567 ( 
.A(n_1406),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1291),
.B(n_1389),
.Y(n_1568)
);

BUFx10_ASAP7_75t_L g1569 ( 
.A(n_1390),
.Y(n_1569)
);

AOI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1385),
.A2(n_1388),
.B(n_1386),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_SL g1571 ( 
.A1(n_1419),
.A2(n_736),
.B1(n_1316),
.B2(n_1304),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1406),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_689),
.B2(n_652),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_689),
.B2(n_652),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1407),
.A2(n_1433),
.B1(n_1183),
.B2(n_823),
.Y(n_1575)
);

BUFx8_ASAP7_75t_L g1576 ( 
.A(n_1280),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1336),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_689),
.B2(n_652),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1406),
.Y(n_1579)
);

OAI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1313),
.A2(n_1173),
.B1(n_973),
.B2(n_1419),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1336),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_1406),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1336),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1423),
.A2(n_1419),
.B1(n_689),
.B2(n_652),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1336),
.Y(n_1585)
);

INVx4_ASAP7_75t_L g1586 ( 
.A(n_1321),
.Y(n_1586)
);

BUFx4f_ASAP7_75t_L g1587 ( 
.A(n_1321),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1407),
.A2(n_1433),
.B1(n_1183),
.B2(n_823),
.Y(n_1588)
);

NAND2x1p5_ASAP7_75t_L g1589 ( 
.A(n_1478),
.B(n_1495),
.Y(n_1589)
);

CKINVDCx8_ASAP7_75t_R g1590 ( 
.A(n_1562),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1472),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1454),
.B(n_1444),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1518),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1445),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1559),
.A2(n_1435),
.B(n_1575),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1486),
.B(n_1540),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1448),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1474),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1476),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1491),
.Y(n_1600)
);

INVx6_ASAP7_75t_L g1601 ( 
.A(n_1569),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1500),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1449),
.B(n_1451),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1470),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1513),
.Y(n_1605)
);

OA21x2_ASAP7_75t_L g1606 ( 
.A1(n_1475),
.A2(n_1570),
.B(n_1494),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1517),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1453),
.B(n_1458),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1487),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1478),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1456),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1456),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1446),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1444),
.B(n_1568),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1519),
.A2(n_1492),
.B(n_1520),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1461),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1509),
.Y(n_1617)
);

INVx4_ASAP7_75t_L g1618 ( 
.A(n_1508),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1439),
.B(n_1524),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1515),
.B(n_1516),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1478),
.B(n_1555),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1518),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1522),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1441),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1507),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1507),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1521),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1526),
.A2(n_1527),
.B1(n_1580),
.B2(n_1436),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1512),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1455),
.Y(n_1630)
);

AOI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1497),
.A2(n_1501),
.B(n_1482),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1526),
.A2(n_1580),
.B1(n_1527),
.B2(n_1438),
.C(n_1544),
.Y(n_1632)
);

OR2x6_ASAP7_75t_L g1633 ( 
.A(n_1462),
.B(n_1499),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1460),
.B(n_1510),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1503),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1546),
.B(n_1547),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1460),
.B(n_1510),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1514),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1483),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1552),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1499),
.B(n_1503),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1577),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1581),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1583),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1585),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1463),
.B(n_1505),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1438),
.A2(n_1588),
.B1(n_1514),
.B2(n_1463),
.C(n_1574),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1511),
.Y(n_1648)
);

O2A1O1Ixp33_ASAP7_75t_SL g1649 ( 
.A1(n_1442),
.A2(n_1563),
.B(n_1558),
.C(n_1579),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1511),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1437),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1534),
.A2(n_1556),
.B1(n_1530),
.B2(n_1533),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1505),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1499),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1489),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1502),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1468),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1468),
.B(n_1466),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1489),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1488),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1488),
.Y(n_1661)
);

OAI21xp33_ASAP7_75t_SL g1662 ( 
.A1(n_1506),
.A2(n_1467),
.B(n_1542),
.Y(n_1662)
);

BUFx2_ASAP7_75t_L g1663 ( 
.A(n_1481),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1496),
.A2(n_1498),
.B(n_1469),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1484),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1519),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1498),
.B(n_1480),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1481),
.B(n_1443),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1520),
.A2(n_1467),
.B(n_1480),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1569),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1493),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1452),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1490),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1473),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1473),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1571),
.B(n_1471),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1447),
.B(n_1564),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1471),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1477),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1440),
.Y(n_1680)
);

OAI21x1_ASAP7_75t_L g1681 ( 
.A1(n_1530),
.A2(n_1533),
.B(n_1553),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1464),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1566),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1529),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1529),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1542),
.A2(n_1578),
.B(n_1554),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_SL g1687 ( 
.A1(n_1553),
.A2(n_1578),
.B1(n_1584),
.B2(n_1573),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1554),
.B(n_1573),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1584),
.B(n_1561),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1529),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1561),
.Y(n_1691)
);

INVx2_ASAP7_75t_SL g1692 ( 
.A(n_1525),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1525),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1525),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1459),
.B(n_1543),
.Y(n_1695)
);

BUFx2_ASAP7_75t_L g1696 ( 
.A(n_1450),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1536),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1551),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1551),
.Y(n_1699)
);

OAI21x1_ASAP7_75t_L g1700 ( 
.A1(n_1551),
.A2(n_1450),
.B(n_1586),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1587),
.A2(n_1539),
.B(n_1565),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1587),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1485),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1504),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1541),
.B(n_1504),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1532),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1582),
.A2(n_1549),
.B(n_1572),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1538),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1567),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1523),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1523),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1479),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1609),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1639),
.B(n_1557),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1654),
.B(n_1537),
.Y(n_1715)
);

A2O1A1Ixp33_ASAP7_75t_L g1716 ( 
.A1(n_1632),
.A2(n_1628),
.B(n_1662),
.C(n_1595),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1594),
.B(n_1531),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1597),
.B(n_1550),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1639),
.B(n_1548),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1611),
.B(n_1528),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1611),
.B(n_1528),
.Y(n_1721)
);

OR2x6_ASAP7_75t_L g1722 ( 
.A(n_1633),
.B(n_1560),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1630),
.A2(n_1535),
.B1(n_1545),
.B2(n_1560),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1616),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1593),
.B(n_1457),
.Y(n_1725)
);

AO32x2_ASAP7_75t_L g1726 ( 
.A1(n_1682),
.A2(n_1535),
.A3(n_1545),
.B1(n_1576),
.B2(n_1465),
.Y(n_1726)
);

A2O1A1Ixp33_ASAP7_75t_L g1727 ( 
.A1(n_1647),
.A2(n_1576),
.B(n_1664),
.C(n_1658),
.Y(n_1727)
);

A2O1A1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1658),
.A2(n_1676),
.B(n_1665),
.C(n_1668),
.Y(n_1728)
);

AO21x1_ASAP7_75t_L g1729 ( 
.A1(n_1614),
.A2(n_1592),
.B(n_1612),
.Y(n_1729)
);

NAND2xp33_ASAP7_75t_L g1730 ( 
.A(n_1683),
.B(n_1613),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1616),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1593),
.B(n_1622),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1612),
.B(n_1630),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1676),
.A2(n_1665),
.B(n_1668),
.C(n_1652),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1672),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1617),
.B(n_1648),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1660),
.A2(n_1661),
.B(n_1657),
.Y(n_1737)
);

O2A1O1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1651),
.A2(n_1673),
.B(n_1671),
.C(n_1660),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1604),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1687),
.A2(n_1688),
.B1(n_1673),
.B2(n_1661),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1617),
.B(n_1648),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1603),
.B(n_1608),
.Y(n_1742)
);

OR2x6_ASAP7_75t_L g1743 ( 
.A(n_1633),
.B(n_1663),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1677),
.B(n_1635),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1646),
.A2(n_1667),
.B(n_1686),
.C(n_1681),
.Y(n_1745)
);

AO32x2_ASAP7_75t_L g1746 ( 
.A1(n_1692),
.A2(n_1670),
.A3(n_1618),
.B1(n_1629),
.B2(n_1650),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_SL g1747 ( 
.A(n_1633),
.B(n_1663),
.Y(n_1747)
);

AOI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1629),
.A2(n_1650),
.B1(n_1637),
.B2(n_1634),
.C(n_1646),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1634),
.A2(n_1637),
.B(n_1667),
.Y(n_1749)
);

O2A1O1Ixp33_ASAP7_75t_SL g1750 ( 
.A1(n_1707),
.A2(n_1703),
.B(n_1708),
.C(n_1711),
.Y(n_1750)
);

AO21x2_ASAP7_75t_L g1751 ( 
.A1(n_1671),
.A2(n_1655),
.B(n_1659),
.Y(n_1751)
);

NOR2xp67_ASAP7_75t_L g1752 ( 
.A(n_1670),
.B(n_1711),
.Y(n_1752)
);

AND2x6_ASAP7_75t_L g1753 ( 
.A(n_1641),
.B(n_1623),
.Y(n_1753)
);

AOI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1653),
.A2(n_1638),
.B1(n_1688),
.B2(n_1659),
.C(n_1655),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1620),
.B(n_1653),
.Y(n_1755)
);

OAI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1596),
.A2(n_1638),
.B1(n_1666),
.B2(n_1674),
.C(n_1675),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1678),
.A2(n_1674),
.B1(n_1675),
.B2(n_1686),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1678),
.A2(n_1681),
.B1(n_1689),
.B2(n_1679),
.Y(n_1758)
);

BUFx2_ASAP7_75t_L g1759 ( 
.A(n_1696),
.Y(n_1759)
);

AO32x2_ASAP7_75t_L g1760 ( 
.A1(n_1692),
.A2(n_1618),
.A3(n_1602),
.B1(n_1642),
.B2(n_1643),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1640),
.B(n_1644),
.Y(n_1761)
);

OA21x2_ASAP7_75t_L g1762 ( 
.A1(n_1615),
.A2(n_1669),
.B(n_1666),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1645),
.B(n_1602),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1672),
.B(n_1590),
.Y(n_1764)
);

AOI21x1_ASAP7_75t_L g1765 ( 
.A1(n_1631),
.A2(n_1696),
.B(n_1704),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1695),
.B(n_1690),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1656),
.B(n_1619),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1636),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1591),
.Y(n_1769)
);

NAND2xp33_ASAP7_75t_L g1770 ( 
.A(n_1683),
.B(n_1613),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1679),
.A2(n_1607),
.B1(n_1605),
.B2(n_1624),
.C(n_1626),
.Y(n_1771)
);

AOI211xp5_ASAP7_75t_L g1772 ( 
.A1(n_1649),
.A2(n_1701),
.B(n_1704),
.C(n_1703),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1693),
.Y(n_1773)
);

AOI21x1_ASAP7_75t_L g1774 ( 
.A1(n_1631),
.A2(n_1625),
.B(n_1691),
.Y(n_1774)
);

OAI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1606),
.A2(n_1700),
.B(n_1589),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1702),
.A2(n_1621),
.B1(n_1706),
.B2(n_1705),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1709),
.Y(n_1777)
);

OA21x2_ASAP7_75t_L g1778 ( 
.A1(n_1627),
.A2(n_1605),
.B(n_1600),
.Y(n_1778)
);

OA21x2_ASAP7_75t_L g1779 ( 
.A1(n_1600),
.A2(n_1599),
.B(n_1591),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1779),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1779),
.Y(n_1781)
);

INVx3_ASAP7_75t_SL g1782 ( 
.A(n_1777),
.Y(n_1782)
);

INVx1_ASAP7_75t_SL g1783 ( 
.A(n_1744),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1742),
.B(n_1606),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_SL g1785 ( 
.A1(n_1740),
.A2(n_1589),
.B1(n_1709),
.B2(n_1706),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1760),
.B(n_1606),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1760),
.B(n_1606),
.Y(n_1787)
);

AND2x4_ASAP7_75t_SL g1788 ( 
.A(n_1722),
.B(n_1610),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1778),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1760),
.B(n_1599),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1739),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1753),
.Y(n_1792)
);

NOR2x1_ASAP7_75t_SL g1793 ( 
.A(n_1722),
.B(n_1684),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1769),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1753),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1724),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1759),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1778),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1762),
.B(n_1598),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1762),
.B(n_1685),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1733),
.B(n_1685),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1733),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1735),
.B(n_1710),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1731),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1732),
.B(n_1775),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1755),
.B(n_1713),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1746),
.B(n_1680),
.Y(n_1807)
);

AOI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1716),
.A2(n_1621),
.B1(n_1601),
.B2(n_1712),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1763),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1746),
.B(n_1766),
.Y(n_1810)
);

AOI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1740),
.A2(n_1697),
.B1(n_1694),
.B2(n_1699),
.C(n_1698),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1773),
.Y(n_1812)
);

INVxp67_ASAP7_75t_SL g1813 ( 
.A(n_1774),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1734),
.A2(n_1601),
.B1(n_1712),
.B2(n_1698),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1736),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1718),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1736),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1791),
.B(n_1750),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1781),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1802),
.B(n_1771),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1780),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1781),
.Y(n_1822)
);

NAND2xp33_ASAP7_75t_SL g1823 ( 
.A(n_1782),
.B(n_1725),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1780),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1781),
.Y(n_1825)
);

INVxp67_ASAP7_75t_L g1826 ( 
.A(n_1800),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1785),
.A2(n_1728),
.B1(n_1727),
.B2(n_1749),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1784),
.B(n_1810),
.Y(n_1828)
);

AO21x2_ASAP7_75t_L g1829 ( 
.A1(n_1813),
.A2(n_1729),
.B(n_1751),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1785),
.A2(n_1738),
.B(n_1745),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1794),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1811),
.A2(n_1737),
.B(n_1749),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1811),
.A2(n_1748),
.B1(n_1722),
.B2(n_1756),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1789),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1789),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1794),
.Y(n_1836)
);

AOI33xp33_ASAP7_75t_L g1837 ( 
.A1(n_1786),
.A2(n_1772),
.A3(n_1757),
.B1(n_1758),
.B2(n_1754),
.B3(n_1768),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1798),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1798),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1795),
.B(n_1765),
.Y(n_1840)
);

BUFx3_ASAP7_75t_L g1841 ( 
.A(n_1792),
.Y(n_1841)
);

NOR2x1_ASAP7_75t_L g1842 ( 
.A(n_1795),
.B(n_1752),
.Y(n_1842)
);

BUFx2_ASAP7_75t_L g1843 ( 
.A(n_1792),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1805),
.B(n_1743),
.Y(n_1844)
);

INVx1_ASAP7_75t_SL g1845 ( 
.A(n_1797),
.Y(n_1845)
);

OAI21xp5_ASAP7_75t_SL g1846 ( 
.A1(n_1808),
.A2(n_1723),
.B(n_1764),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1796),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1802),
.B(n_1761),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1798),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1796),
.Y(n_1850)
);

INVxp67_ASAP7_75t_SL g1851 ( 
.A(n_1812),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1806),
.B(n_1761),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1799),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1815),
.B(n_1751),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1804),
.Y(n_1855)
);

OAI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1814),
.A2(n_1747),
.B1(n_1737),
.B2(n_1776),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1805),
.B(n_1721),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1804),
.Y(n_1858)
);

INVxp67_ASAP7_75t_SL g1859 ( 
.A(n_1786),
.Y(n_1859)
);

BUFx3_ASAP7_75t_L g1860 ( 
.A(n_1788),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1786),
.B(n_1721),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1787),
.B(n_1720),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1787),
.B(n_1720),
.Y(n_1863)
);

AOI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1787),
.A2(n_1741),
.B1(n_1772),
.B2(n_1723),
.C(n_1767),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1820),
.B(n_1817),
.Y(n_1865)
);

INVx4_ASAP7_75t_L g1866 ( 
.A(n_1841),
.Y(n_1866)
);

INVx1_ASAP7_75t_SL g1867 ( 
.A(n_1845),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1841),
.B(n_1793),
.Y(n_1868)
);

INVx1_ASAP7_75t_SL g1869 ( 
.A(n_1845),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1853),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1828),
.B(n_1783),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1820),
.B(n_1817),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1853),
.Y(n_1873)
);

NOR3xp33_ASAP7_75t_L g1874 ( 
.A(n_1864),
.B(n_1830),
.C(n_1827),
.Y(n_1874)
);

INVx2_ASAP7_75t_SL g1875 ( 
.A(n_1842),
.Y(n_1875)
);

BUFx2_ASAP7_75t_L g1876 ( 
.A(n_1823),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1859),
.B(n_1806),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1828),
.B(n_1783),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1831),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1831),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1823),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1848),
.B(n_1809),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1836),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1843),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1821),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1836),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1828),
.B(n_1797),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1859),
.B(n_1807),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1847),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1841),
.B(n_1793),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1847),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1852),
.B(n_1801),
.Y(n_1892)
);

AND2x2_ASAP7_75t_SL g1893 ( 
.A(n_1837),
.B(n_1747),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1852),
.B(n_1801),
.Y(n_1894)
);

AND2x4_ASAP7_75t_L g1895 ( 
.A(n_1841),
.B(n_1790),
.Y(n_1895)
);

INVx2_ASAP7_75t_SL g1896 ( 
.A(n_1840),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1852),
.B(n_1824),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1850),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1876),
.B(n_1881),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1867),
.B(n_1782),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1879),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1876),
.B(n_1861),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1874),
.B(n_1850),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1879),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1880),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1874),
.B(n_1855),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1870),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1865),
.B(n_1855),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1881),
.B(n_1861),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1868),
.B(n_1861),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1870),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1883),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1867),
.B(n_1869),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1892),
.B(n_1851),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1870),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1865),
.B(n_1858),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1883),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1868),
.B(n_1844),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1868),
.B(n_1862),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1886),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1868),
.B(n_1862),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1872),
.B(n_1858),
.Y(n_1922)
);

BUFx2_ASAP7_75t_L g1923 ( 
.A(n_1866),
.Y(n_1923)
);

OAI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1893),
.A2(n_1832),
.B(n_1864),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1886),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1872),
.B(n_1862),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1889),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1868),
.B(n_1863),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1890),
.B(n_1863),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1872),
.B(n_1863),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1889),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1873),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1891),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1892),
.B(n_1851),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1891),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1898),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1890),
.B(n_1871),
.Y(n_1937)
);

BUFx3_ASAP7_75t_L g1938 ( 
.A(n_1869),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1873),
.Y(n_1939)
);

NAND2x1p5_ASAP7_75t_L g1940 ( 
.A(n_1866),
.B(n_1860),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1890),
.B(n_1844),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1890),
.B(n_1857),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1898),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1885),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1884),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1894),
.B(n_1857),
.Y(n_1946)
);

INVx2_ASAP7_75t_SL g1947 ( 
.A(n_1890),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1903),
.B(n_1897),
.Y(n_1948)
);

INVx1_ASAP7_75t_SL g1949 ( 
.A(n_1938),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1902),
.B(n_1866),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1903),
.B(n_1906),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1900),
.B(n_1782),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1901),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1901),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1906),
.B(n_1884),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1938),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1938),
.Y(n_1957)
);

AOI211xp5_ASAP7_75t_L g1958 ( 
.A1(n_1924),
.A2(n_1846),
.B(n_1827),
.C(n_1830),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1904),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1924),
.B(n_1887),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1902),
.B(n_1866),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1945),
.B(n_1887),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1913),
.B(n_1887),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1899),
.B(n_1893),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1909),
.B(n_1899),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1946),
.B(n_1926),
.Y(n_1966)
);

OAI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1909),
.A2(n_1893),
.B(n_1818),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_1923),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1904),
.Y(n_1969)
);

OR2x6_ASAP7_75t_L g1970 ( 
.A(n_1940),
.B(n_1832),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1918),
.B(n_1818),
.Y(n_1971)
);

OAI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1926),
.A2(n_1833),
.B1(n_1856),
.B2(n_1814),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1907),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1930),
.B(n_1894),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1942),
.B(n_1871),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1905),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1946),
.B(n_1816),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1942),
.B(n_1871),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1940),
.B(n_1878),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1940),
.B(n_1878),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1918),
.B(n_1941),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1918),
.B(n_1896),
.Y(n_1982)
);

INVx1_ASAP7_75t_SL g1983 ( 
.A(n_1923),
.Y(n_1983)
);

HB1xp67_ASAP7_75t_L g1984 ( 
.A(n_1944),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1918),
.B(n_1896),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1941),
.B(n_1878),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1905),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1930),
.B(n_1882),
.Y(n_1988)
);

AOI21xp33_ASAP7_75t_SL g1989 ( 
.A1(n_1951),
.A2(n_1947),
.B(n_1875),
.Y(n_1989)
);

NAND3xp33_ASAP7_75t_L g1990 ( 
.A(n_1958),
.B(n_1944),
.C(n_1837),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1957),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_SL g1992 ( 
.A1(n_1967),
.A2(n_1960),
.B1(n_1957),
.B2(n_1970),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1953),
.Y(n_1993)
);

AOI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1958),
.A2(n_1964),
.B1(n_1967),
.B2(n_1972),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1949),
.B(n_1922),
.Y(n_1995)
);

OAI211xp5_ASAP7_75t_SL g1996 ( 
.A1(n_1955),
.A2(n_1947),
.B(n_1934),
.C(n_1914),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1953),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1954),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1954),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1957),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1959),
.Y(n_2001)
);

AND2x4_ASAP7_75t_L g2002 ( 
.A(n_1949),
.B(n_1941),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1948),
.B(n_1914),
.Y(n_2003)
);

NOR3xp33_ASAP7_75t_L g2004 ( 
.A(n_1956),
.B(n_1833),
.C(n_1846),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1956),
.B(n_1922),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1970),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1977),
.B(n_1730),
.Y(n_2007)
);

AOI221xp5_ASAP7_75t_L g2008 ( 
.A1(n_1948),
.A2(n_1888),
.B1(n_1916),
.B2(n_1908),
.C(n_1826),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1959),
.Y(n_2009)
);

AND3x1_ASAP7_75t_L g2010 ( 
.A(n_1965),
.B(n_1937),
.C(n_1875),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1969),
.Y(n_2011)
);

AOI211xp5_ASAP7_75t_L g2012 ( 
.A1(n_1971),
.A2(n_1888),
.B(n_1896),
.C(n_1856),
.Y(n_2012)
);

AOI221xp5_ASAP7_75t_L g2013 ( 
.A1(n_1988),
.A2(n_1888),
.B1(n_1908),
.B2(n_1916),
.C(n_1826),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1952),
.B(n_1770),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1969),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1965),
.B(n_1968),
.Y(n_2016)
);

OAI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1970),
.A2(n_1961),
.B(n_1950),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1981),
.B(n_1937),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1976),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1993),
.Y(n_2020)
);

INVx1_ASAP7_75t_SL g2021 ( 
.A(n_2002),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1997),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1998),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_2002),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1991),
.B(n_1968),
.Y(n_2025)
);

INVxp67_ASAP7_75t_L g2026 ( 
.A(n_2016),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1991),
.B(n_1981),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_2000),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1999),
.Y(n_2029)
);

OR2x2_ASAP7_75t_L g2030 ( 
.A(n_1990),
.B(n_1966),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2001),
.Y(n_2031)
);

AOI31xp33_ASAP7_75t_L g2032 ( 
.A1(n_1992),
.A2(n_1983),
.A3(n_1950),
.B(n_1961),
.Y(n_2032)
);

OAI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_1994),
.A2(n_1970),
.B1(n_1877),
.B2(n_1875),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2009),
.Y(n_2034)
);

XNOR2xp5_ASAP7_75t_L g2035 ( 
.A(n_1992),
.B(n_1970),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_2000),
.B(n_1983),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_2010),
.A2(n_1962),
.B1(n_1941),
.B2(n_1986),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_2003),
.B(n_1966),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_2004),
.B(n_1984),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_2018),
.B(n_1986),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_2006),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_2004),
.B(n_1975),
.Y(n_2042)
);

AOI221x1_ASAP7_75t_SL g2043 ( 
.A1(n_2012),
.A2(n_1982),
.B1(n_1985),
.B2(n_1963),
.C(n_1987),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2028),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2038),
.Y(n_2045)
);

INVxp67_ASAP7_75t_L g2046 ( 
.A(n_2036),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2038),
.Y(n_2047)
);

AOI222xp33_ASAP7_75t_L g2048 ( 
.A1(n_2035),
.A2(n_2006),
.B1(n_1996),
.B2(n_2008),
.C1(n_1995),
.C2(n_2005),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2024),
.Y(n_2049)
);

OAI21xp5_ASAP7_75t_L g2050 ( 
.A1(n_2035),
.A2(n_2017),
.B(n_1989),
.Y(n_2050)
);

XNOR2x2_ASAP7_75t_L g2051 ( 
.A(n_2030),
.B(n_2014),
.Y(n_2051)
);

OAI222xp33_ASAP7_75t_L g2052 ( 
.A1(n_2030),
.A2(n_2019),
.B1(n_2015),
.B2(n_2011),
.C1(n_1973),
.C2(n_1985),
.Y(n_2052)
);

AOI222xp33_ASAP7_75t_L g2053 ( 
.A1(n_2039),
.A2(n_2013),
.B1(n_1973),
.B2(n_1976),
.C1(n_1987),
.C2(n_1988),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2043),
.B(n_1974),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_2021),
.B(n_2007),
.Y(n_2055)
);

OAI21xp5_ASAP7_75t_SL g2056 ( 
.A1(n_2032),
.A2(n_2014),
.B(n_1980),
.Y(n_2056)
);

OAI322xp33_ASAP7_75t_L g2057 ( 
.A1(n_2033),
.A2(n_1934),
.A3(n_1973),
.B1(n_1877),
.B2(n_1917),
.C1(n_1925),
.C2(n_1912),
.Y(n_2057)
);

OAI221xp5_ASAP7_75t_L g2058 ( 
.A1(n_2042),
.A2(n_1911),
.B1(n_1939),
.B2(n_1915),
.C(n_1907),
.Y(n_2058)
);

NAND4xp25_ASAP7_75t_L g2059 ( 
.A(n_2055),
.B(n_2036),
.C(n_2026),
.D(n_2024),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2045),
.Y(n_2060)
);

INVx1_ASAP7_75t_SL g2061 ( 
.A(n_2051),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_2047),
.B(n_2025),
.Y(n_2062)
);

OAI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_2046),
.A2(n_2027),
.B(n_2037),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2044),
.B(n_2027),
.Y(n_2064)
);

NOR3xp33_ASAP7_75t_SL g2065 ( 
.A(n_2052),
.B(n_2022),
.C(n_2020),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2053),
.B(n_2027),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2049),
.Y(n_2067)
);

OAI21xp5_ASAP7_75t_SL g2068 ( 
.A1(n_2048),
.A2(n_2040),
.B(n_1980),
.Y(n_2068)
);

INVxp67_ASAP7_75t_L g2069 ( 
.A(n_2050),
.Y(n_2069)
);

NOR4xp25_ASAP7_75t_L g2070 ( 
.A(n_2054),
.B(n_2034),
.C(n_2031),
.D(n_2029),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_2056),
.B(n_2007),
.Y(n_2071)
);

AOI221xp5_ASAP7_75t_L g2072 ( 
.A1(n_2061),
.A2(n_2057),
.B1(n_2054),
.B2(n_2058),
.C(n_2023),
.Y(n_2072)
);

AOI211xp5_ASAP7_75t_L g2073 ( 
.A1(n_2068),
.A2(n_2041),
.B(n_2040),
.C(n_1985),
.Y(n_2073)
);

NOR4xp25_ASAP7_75t_L g2074 ( 
.A(n_2069),
.B(n_2066),
.C(n_2059),
.D(n_2067),
.Y(n_2074)
);

AOI221xp5_ASAP7_75t_L g2075 ( 
.A1(n_2069),
.A2(n_1911),
.B1(n_1907),
.B2(n_1915),
.C(n_1932),
.Y(n_2075)
);

AOI221xp5_ASAP7_75t_L g2076 ( 
.A1(n_2065),
.A2(n_1932),
.B1(n_1939),
.B2(n_1915),
.C(n_1911),
.Y(n_2076)
);

OAI221xp5_ASAP7_75t_L g2077 ( 
.A1(n_2070),
.A2(n_1932),
.B1(n_1939),
.B2(n_1979),
.C(n_1590),
.Y(n_2077)
);

AOI221xp5_ASAP7_75t_L g2078 ( 
.A1(n_2060),
.A2(n_1985),
.B1(n_1982),
.B2(n_1813),
.C(n_1979),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_L g2079 ( 
.A(n_2077),
.B(n_2071),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_2073),
.B(n_2063),
.Y(n_2080)
);

OAI211xp5_ASAP7_75t_L g2081 ( 
.A1(n_2074),
.A2(n_2064),
.B(n_2062),
.C(n_1712),
.Y(n_2081)
);

AOI211xp5_ASAP7_75t_SL g2082 ( 
.A1(n_2072),
.A2(n_1982),
.B(n_1978),
.C(n_1975),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_2076),
.A2(n_1829),
.B1(n_1982),
.B2(n_1834),
.Y(n_2083)
);

BUFx12f_ASAP7_75t_L g2084 ( 
.A(n_2078),
.Y(n_2084)
);

AOI221xp5_ASAP7_75t_L g2085 ( 
.A1(n_2075),
.A2(n_1895),
.B1(n_1943),
.B2(n_1936),
.C(n_1935),
.Y(n_2085)
);

AOI222xp33_ASAP7_75t_L g2086 ( 
.A1(n_2072),
.A2(n_1819),
.B1(n_1849),
.B2(n_1839),
.C1(n_1838),
.C2(n_1835),
.Y(n_2086)
);

AOI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_2086),
.A2(n_1978),
.B1(n_1895),
.B2(n_1921),
.Y(n_2087)
);

NAND4xp75_ASAP7_75t_L g2088 ( 
.A(n_2079),
.B(n_1910),
.C(n_1919),
.D(n_1921),
.Y(n_2088)
);

NAND4xp75_ASAP7_75t_L g2089 ( 
.A(n_2081),
.B(n_1910),
.C(n_1928),
.D(n_1929),
.Y(n_2089)
);

AO22x2_ASAP7_75t_L g2090 ( 
.A1(n_2080),
.A2(n_1717),
.B1(n_1936),
.B2(n_1935),
.Y(n_2090)
);

NOR3xp33_ASAP7_75t_L g2091 ( 
.A(n_2085),
.B(n_1726),
.C(n_1854),
.Y(n_2091)
);

AND2x2_ASAP7_75t_SL g2092 ( 
.A(n_2082),
.B(n_1712),
.Y(n_2092)
);

AOI211xp5_ASAP7_75t_L g2093 ( 
.A1(n_2091),
.A2(n_2084),
.B(n_2092),
.C(n_2087),
.Y(n_2093)
);

OAI221xp5_ASAP7_75t_L g2094 ( 
.A1(n_2090),
.A2(n_2083),
.B1(n_1943),
.B2(n_1933),
.C(n_1931),
.Y(n_2094)
);

AOI211xp5_ASAP7_75t_L g2095 ( 
.A1(n_2089),
.A2(n_1726),
.B(n_1929),
.C(n_1928),
.Y(n_2095)
);

INVxp67_ASAP7_75t_L g2096 ( 
.A(n_2088),
.Y(n_2096)
);

HB1xp67_ASAP7_75t_L g2097 ( 
.A(n_2096),
.Y(n_2097)
);

AO22x2_ASAP7_75t_L g2098 ( 
.A1(n_2093),
.A2(n_1933),
.B1(n_1931),
.B2(n_1927),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2097),
.Y(n_2099)
);

AO22x2_ASAP7_75t_L g2100 ( 
.A1(n_2099),
.A2(n_2098),
.B1(n_2095),
.B2(n_2094),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2099),
.Y(n_2101)
);

HB1xp67_ASAP7_75t_L g2102 ( 
.A(n_2101),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2100),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2102),
.A2(n_1819),
.B1(n_1822),
.B2(n_1825),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2104),
.B(n_2103),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2105),
.B(n_1714),
.Y(n_2106)
);

AOI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_2106),
.A2(n_1927),
.B1(n_1925),
.B2(n_1920),
.Y(n_2107)
);

AOI221xp5_ASAP7_75t_L g2108 ( 
.A1(n_2107),
.A2(n_1803),
.B1(n_1920),
.B2(n_1917),
.C(n_1912),
.Y(n_2108)
);

AOI211xp5_ASAP7_75t_L g2109 ( 
.A1(n_2108),
.A2(n_1726),
.B(n_1715),
.C(n_1719),
.Y(n_2109)
);


endmodule