module fake_netlist_6_3217_n_409 (n_41, n_52, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_54, n_27, n_3, n_14, n_38, n_0, n_61, n_39, n_63, n_60, n_59, n_32, n_4, n_66, n_36, n_22, n_26, n_55, n_13, n_35, n_11, n_28, n_17, n_23, n_58, n_12, n_20, n_50, n_49, n_7, n_30, n_64, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_62, n_31, n_65, n_25, n_40, n_57, n_53, n_51, n_44, n_56, n_409);

input n_41;
input n_52;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_54;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_61;
input n_39;
input n_63;
input n_60;
input n_59;
input n_32;
input n_4;
input n_66;
input n_36;
input n_22;
input n_26;
input n_55;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_58;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_64;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_62;
input n_31;
input n_65;
input n_25;
input n_40;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_409;

wire n_91;
wire n_326;
wire n_256;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_68;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_77;
wire n_106;
wire n_358;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_78;
wire n_84;
wire n_392;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_67;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_230;
wire n_141;
wire n_383;
wire n_200;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_71;
wire n_74;
wire n_229;
wire n_305;
wire n_72;
wire n_173;
wire n_250;
wire n_372;
wire n_111;
wire n_314;
wire n_378;
wire n_377;
wire n_183;
wire n_79;
wire n_375;
wire n_338;
wire n_360;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_344;
wire n_73;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_96;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_397;
wire n_155;
wire n_109;
wire n_122;
wire n_218;
wire n_70;
wire n_234;
wire n_381;
wire n_82;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_97;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_93;
wire n_80;
wire n_196;
wire n_402;
wire n_352;
wire n_107;
wire n_89;
wire n_374;
wire n_366;
wire n_407;
wire n_103;
wire n_272;
wire n_185;
wire n_348;
wire n_69;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_83;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_152;
wire n_92;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_406;
wire n_102;
wire n_204;
wire n_261;
wire n_312;
wire n_394;
wire n_130;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_76;
wire n_243;
wire n_124;
wire n_94;
wire n_282;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_95;
wire n_311;
wire n_403;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_88;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_317;
wire n_149;
wire n_90;
wire n_347;
wire n_328;
wire n_373;
wire n_87;
wire n_195;
wire n_285;
wire n_85;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_75;
wire n_401;
wire n_324;
wire n_335;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_81;
wire n_267;
wire n_339;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_351;
wire n_259;
wire n_177;
wire n_391;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_39),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_8),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_22),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_33),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_17),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_31),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_9),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_11),
.Y(n_99)
);

INVxp33_ASAP7_75t_SL g100 ( 
.A(n_21),
.Y(n_100)
);

INVxp33_ASAP7_75t_SL g101 ( 
.A(n_7),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_48),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_17),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_0),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_1),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_52),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_15),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_18),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_12),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_1),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_5),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_18),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_10),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_0),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_8),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_44),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_5),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_14),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_67),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_67),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_69),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_3),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_69),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_80),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_80),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_88),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_85),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_88),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_87),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_R g146 ( 
.A(n_102),
.B(n_37),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_87),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_R g149 ( 
.A(n_102),
.B(n_75),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_R g150 ( 
.A(n_75),
.B(n_40),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_4),
.Y(n_152)
);

NOR2x1p5_ASAP7_75t_L g153 ( 
.A(n_96),
.B(n_78),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_105),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_91),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_105),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_91),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_93),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

OR2x6_ASAP7_75t_L g164 ( 
.A(n_96),
.B(n_6),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

AND2x4_ASAP7_75t_L g167 ( 
.A(n_78),
.B(n_42),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_98),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_108),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_118),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_99),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_70),
.B(n_6),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_115),
.Y(n_178)
);

OAI21x1_ASAP7_75t_L g179 ( 
.A1(n_123),
.A2(n_7),
.B(n_10),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_83),
.Y(n_181)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_116),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_13),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_100),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_126),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_100),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_101),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_167),
.B(n_101),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_155),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_123),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_81),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_126),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_133),
.A2(n_125),
.B1(n_109),
.B2(n_90),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_76),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_73),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

NOR2x1p5_ASAP7_75t_L g209 ( 
.A(n_152),
.B(n_161),
.Y(n_209)
);

AND2x4_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_77),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

AO22x2_ASAP7_75t_L g212 ( 
.A1(n_164),
.A2(n_113),
.B1(n_111),
.B2(n_110),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_148),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_146),
.B(n_106),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_97),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_142),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_86),
.Y(n_220)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_170),
.B(n_92),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_128),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_82),
.B1(n_79),
.B2(n_15),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_163),
.Y(n_225)
);

BUFx8_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

NAND2x1p5_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_49),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_175),
.B(n_53),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_177),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_140),
.B(n_16),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_55),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_179),
.A2(n_16),
.B(n_20),
.C(n_25),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_171),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_131),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_173),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_194),
.A2(n_186),
.B(n_184),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_209),
.Y(n_242)
);

BUFx8_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_191),
.B(n_172),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_194),
.A2(n_178),
.B(n_185),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_136),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_205),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_192),
.B(n_150),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_134),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_213),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_SL g254 ( 
.A1(n_189),
.A2(n_187),
.B(n_174),
.Y(n_254)
);

OAI22x1_ASAP7_75t_L g255 ( 
.A1(n_195),
.A2(n_141),
.B1(n_145),
.B2(n_143),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_192),
.B(n_220),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_216),
.A2(n_138),
.B(n_139),
.Y(n_257)
);

AND3x4_ASAP7_75t_L g258 ( 
.A(n_210),
.B(n_132),
.C(n_158),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

BUFx4f_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_196),
.B(n_32),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_216),
.A2(n_59),
.B(n_60),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_224),
.A2(n_142),
.B1(n_147),
.B2(n_154),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_220),
.A2(n_61),
.B(n_197),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_196),
.B(n_193),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_198),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_SL g268 ( 
.A1(n_200),
.A2(n_199),
.B(n_202),
.C(n_230),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_218),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_196),
.B(n_232),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_210),
.B(n_206),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_210),
.A2(n_215),
.B(n_212),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_215),
.A2(n_212),
.B(n_207),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_214),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_212),
.A2(n_206),
.B(n_207),
.Y(n_276)
);

NAND2x1p5_ASAP7_75t_L g277 ( 
.A(n_219),
.B(n_222),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_234),
.A2(n_221),
.B1(n_235),
.B2(n_233),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_228),
.A2(n_237),
.B(n_221),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_223),
.B(n_226),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_225),
.B(n_231),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_231),
.B(n_227),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_208),
.Y(n_283)
);

CKINVDCx8_ASAP7_75t_R g284 ( 
.A(n_223),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_228),
.A2(n_227),
.B1(n_211),
.B2(n_217),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_237),
.A2(n_208),
.B(n_211),
.C(n_217),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_221),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_226),
.B(n_218),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_221),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_279),
.A2(n_289),
.B(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_270),
.Y(n_293)
);

INVx8_ASAP7_75t_L g294 ( 
.A(n_260),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_270),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_269),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_249),
.B(n_275),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_253),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_260),
.A2(n_271),
.B1(n_256),
.B2(n_240),
.Y(n_302)
);

BUFx4f_ASAP7_75t_SL g303 ( 
.A(n_243),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_271),
.A2(n_278),
.B1(n_240),
.B2(n_244),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_251),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_274),
.B(n_265),
.Y(n_307)
);

BUFx4_ASAP7_75t_SL g308 ( 
.A(n_258),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_259),
.Y(n_310)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_287),
.A2(n_262),
.B(n_263),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_266),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_242),
.B(n_241),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_262),
.A2(n_285),
.B1(n_261),
.B2(n_246),
.Y(n_315)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_277),
.A2(n_257),
.B(n_286),
.Y(n_316)
);

AO32x2_ASAP7_75t_L g317 ( 
.A1(n_264),
.A2(n_268),
.A3(n_255),
.B1(n_288),
.B2(n_280),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_192),
.Y(n_318)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

OA21x2_ASAP7_75t_L g320 ( 
.A1(n_286),
.A2(n_279),
.B(n_276),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_272),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g323 ( 
.A1(n_279),
.A2(n_289),
.B(n_276),
.Y(n_323)
);

OR2x6_ASAP7_75t_L g324 ( 
.A(n_273),
.B(n_276),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_279),
.A2(n_272),
.B(n_271),
.Y(n_325)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_279),
.A2(n_289),
.B(n_276),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_260),
.Y(n_327)
);

CKINVDCx11_ASAP7_75t_R g328 ( 
.A(n_284),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_245),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_245),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_248),
.A2(n_252),
.B1(n_234),
.B2(n_131),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_328),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_R g334 ( 
.A(n_328),
.B(n_298),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_308),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_322),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_303),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_318),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_295),
.Y(n_340)
);

CKINVDCx11_ASAP7_75t_R g341 ( 
.A(n_297),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_293),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_306),
.A2(n_321),
.B1(n_302),
.B2(n_304),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_310),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_332),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_325),
.Y(n_347)
);

NOR3xp33_ASAP7_75t_SL g348 ( 
.A(n_313),
.B(n_301),
.C(n_299),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

AOI221xp5_ASAP7_75t_L g350 ( 
.A1(n_291),
.A2(n_296),
.B1(n_315),
.B2(n_313),
.C(n_300),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_305),
.B(n_309),
.Y(n_351)
);

NAND4xp25_ASAP7_75t_L g352 ( 
.A(n_300),
.B(n_314),
.C(n_317),
.D(n_330),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_327),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_331),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_294),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_324),
.A2(n_320),
.B1(n_331),
.B2(n_329),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_R g357 ( 
.A(n_320),
.B(n_324),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_294),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_316),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_290),
.B(n_326),
.Y(n_360)
);

CKINVDCx11_ASAP7_75t_R g361 ( 
.A(n_317),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_329),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_361),
.A2(n_329),
.B1(n_327),
.B2(n_319),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_346),
.A2(n_347),
.B1(n_352),
.B2(n_350),
.Y(n_365)
);

INVx4_ASAP7_75t_R g366 ( 
.A(n_359),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_323),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_307),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_346),
.A2(n_311),
.B1(n_336),
.B2(n_359),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_342),
.Y(n_371)
);

OAI221xp5_ASAP7_75t_L g372 ( 
.A1(n_351),
.A2(n_344),
.B1(n_348),
.B2(n_356),
.C(n_357),
.Y(n_372)
);

OA21x2_ASAP7_75t_L g373 ( 
.A1(n_360),
.A2(n_345),
.B(n_354),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_334),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_354),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_355),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_363),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_353),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_362),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_373),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_345),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_343),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_343),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_358),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_374),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_378),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_381),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_368),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_371),
.Y(n_390)
);

NOR2x1_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_374),
.Y(n_391)
);

OAI322xp33_ASAP7_75t_L g392 ( 
.A1(n_390),
.A2(n_386),
.A3(n_371),
.B1(n_375),
.B2(n_379),
.C1(n_385),
.C2(n_380),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_383),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_391),
.A2(n_341),
.B1(n_384),
.B2(n_377),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_388),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_388),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_389),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_395),
.B(n_396),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_394),
.A2(n_377),
.B1(n_370),
.B2(n_358),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_399),
.A2(n_392),
.B1(n_333),
.B2(n_383),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_398),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_401),
.B(n_397),
.Y(n_402)
);

NAND3x1_ASAP7_75t_SL g403 ( 
.A(n_400),
.B(n_366),
.C(n_337),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_402),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_404),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_405),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_406),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_407),
.A2(n_401),
.B1(n_403),
.B2(n_335),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_408),
.A2(n_337),
.B(n_335),
.Y(n_409)
);


endmodule