module fake_jpeg_4186_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_33),
.Y(n_71)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_30),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_30),
.B1(n_21),
.B2(n_20),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_38),
.A2(n_30),
.B1(n_21),
.B2(n_20),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_40),
.Y(n_99)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_57),
.B1(n_18),
.B2(n_60),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_76),
.A2(n_100),
.B1(n_59),
.B2(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_88),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_21),
.B1(n_59),
.B2(n_73),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_85),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_97),
.Y(n_114)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_72),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_33),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_56),
.A2(n_30),
.B1(n_21),
.B2(n_36),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_101),
.B(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_106),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_119),
.B1(n_89),
.B2(n_87),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_66),
.B(n_39),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_109),
.B1(n_116),
.B2(n_118),
.Y(n_135)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_18),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_51),
.B(n_67),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_120),
.C(n_126),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_65),
.B1(n_74),
.B2(n_68),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_113),
.A2(n_115),
.B1(n_117),
.B2(n_95),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_83),
.B1(n_65),
.B2(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_66),
.B1(n_48),
.B2(n_49),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_62),
.B1(n_97),
.B2(n_96),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_64),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_55),
.B(n_64),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_55),
.B1(n_62),
.B2(n_32),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_123),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_35),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_28),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_35),
.C(n_41),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_28),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_129),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_128),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_87),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_132),
.B1(n_151),
.B2(n_107),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_79),
.B1(n_95),
.B2(n_61),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_124),
.C(n_116),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_138),
.C(n_139),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_82),
.C(n_54),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_54),
.C(n_41),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_25),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_145),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_25),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_114),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_17),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_157),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_158),
.B1(n_127),
.B2(n_32),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_63),
.B1(n_92),
.B2(n_19),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_105),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_152),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_125),
.Y(n_165)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_109),
.A2(n_78),
.B1(n_19),
.B2(n_23),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_159),
.B(n_161),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_117),
.B(n_104),
.C(n_108),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_152),
.B(n_108),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_186),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_168),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_128),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_112),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_177),
.C(n_148),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_133),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_172),
.Y(n_202)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_183),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_182),
.B1(n_168),
.B2(n_186),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_115),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_140),
.A2(n_111),
.B(n_102),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_145),
.B(n_147),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_111),
.B(n_127),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_181),
.B(n_28),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_135),
.A2(n_111),
.B(n_127),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_106),
.B1(n_122),
.B2(n_118),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_184),
.A2(n_157),
.B1(n_156),
.B2(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_84),
.B1(n_23),
.B2(n_32),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_187),
.A2(n_141),
.B1(n_154),
.B2(n_131),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_188),
.A2(n_198),
.B(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_190),
.B(n_191),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_194),
.Y(n_223)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_208),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_142),
.B(n_137),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_156),
.B1(n_139),
.B2(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_153),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_203),
.C(n_207),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_143),
.B1(n_23),
.B2(n_33),
.Y(n_204)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_29),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_210),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_31),
.B(n_24),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_213),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_90),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_215),
.C(n_164),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_175),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_166),
.B1(n_159),
.B2(n_162),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_167),
.C(n_178),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_242),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_164),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_193),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_199),
.C(n_209),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_179),
.C(n_184),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_225),
.C(n_231),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_174),
.C(n_161),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_191),
.A2(n_185),
.B1(n_172),
.B2(n_187),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_229),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_185),
.B1(n_26),
.B2(n_90),
.Y(n_230)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_78),
.C(n_24),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_192),
.B1(n_210),
.B2(n_211),
.Y(n_232)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_26),
.B1(n_34),
.B2(n_24),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_233),
.Y(n_244)
);

XNOR2x2_ASAP7_75t_SL g237 ( 
.A(n_188),
.B(n_206),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_237),
.B(n_204),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_24),
.C(n_29),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_200),
.C(n_198),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_240),
.A2(n_196),
.B(n_189),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_190),
.A2(n_26),
.B1(n_34),
.B2(n_24),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_224),
.B1(n_228),
.B2(n_217),
.Y(n_262)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_255),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_249),
.C(n_252),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_240),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_258),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_208),
.C(n_24),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_242),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_24),
.C(n_31),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_256),
.C(n_257),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_29),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_29),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_29),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_232),
.B(n_29),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_29),
.Y(n_263)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_34),
.B1(n_26),
.B2(n_3),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_230),
.B1(n_234),
.B2(n_241),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_236),
.B(n_31),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_236),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_274),
.B1(n_265),
.B2(n_34),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_222),
.C(n_231),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_280),
.C(n_284),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_229),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_277),
.Y(n_294)
);

OA21x2_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_223),
.B(n_226),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_278),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_239),
.C(n_235),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_220),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_281),
.B(n_282),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_245),
.B(n_233),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_16),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_246),
.B(n_256),
.C(n_248),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_31),
.C(n_22),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_31),
.C(n_22),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_266),
.B1(n_245),
.B2(n_244),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_286),
.A2(n_287),
.B1(n_0),
.B2(n_2),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_263),
.B1(n_258),
.B2(n_253),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_257),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_289),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_251),
.Y(n_289)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_298),
.B(n_285),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_299),
.C(n_272),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_296),
.B(n_301),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_268),
.B(n_31),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_300),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_0),
.C(n_2),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_278),
.B(n_15),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_278),
.A2(n_13),
.B1(n_12),
.B2(n_3),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_273),
.Y(n_302)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_275),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_304),
.B(n_306),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_271),
.C(n_280),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_SL g321 ( 
.A(n_308),
.B(n_288),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_271),
.C(n_272),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_309),
.A2(n_314),
.B(n_315),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_13),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_4),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_297),
.B1(n_5),
.B2(n_6),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_299),
.A2(n_2),
.B(n_3),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_2),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_287),
.B1(n_300),
.B2(n_298),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_316),
.A2(n_321),
.B1(n_322),
.B2(n_324),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_295),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_318),
.B(n_325),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_4),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_4),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_304),
.A2(n_309),
.B1(n_310),
.B2(n_307),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_323),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_4),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_319),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_329),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_311),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_317),
.A2(n_311),
.B(n_6),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_330),
.A2(n_7),
.B(n_8),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_331),
.A2(n_333),
.B(n_7),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_316),
.A2(n_7),
.B(n_8),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_324),
.B(n_8),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_336),
.C(n_338),
.Y(n_340)
);

AOI221xp5_ASAP7_75t_SL g341 ( 
.A1(n_337),
.A2(n_327),
.B1(n_10),
.B2(n_11),
.C(n_9),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_332),
.A2(n_9),
.B(n_10),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_332),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_340),
.C(n_339),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_9),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_11),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_345),
.B(n_11),
.Y(n_346)
);


endmodule