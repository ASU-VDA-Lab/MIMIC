module fake_jpeg_3904_n_332 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_8),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_23),
.Y(n_41)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_44),
.B(n_22),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_48),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_49),
.B(n_27),
.Y(n_90)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_62),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_17),
.B1(n_34),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_56),
.A2(n_61),
.B1(n_79),
.B2(n_85),
.Y(n_129)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_28),
.B1(n_24),
.B2(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_30),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_65),
.B(n_82),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_66),
.Y(n_104)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_17),
.B1(n_34),
.B2(n_28),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_100),
.B1(n_101),
.B2(n_18),
.Y(n_113)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_74),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_75),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_36),
.B(n_22),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_77),
.A2(n_98),
.B(n_29),
.C(n_26),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_39),
.A2(n_17),
.B1(n_15),
.B2(n_14),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_81),
.Y(n_118)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_30),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_16),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_84),
.Y(n_130)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_43),
.A2(n_25),
.B1(n_32),
.B2(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_16),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_92),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_25),
.B1(n_15),
.B2(n_20),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_91),
.B1(n_21),
.B2(n_32),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_37),
.A2(n_14),
.B1(n_15),
.B2(n_19),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_97),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_47),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_37),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_44),
.B(n_21),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_21),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_48),
.A2(n_27),
.B1(n_20),
.B2(n_31),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_48),
.A2(n_32),
.B1(n_31),
.B2(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_105),
.B(n_121),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_107),
.A2(n_74),
.B1(n_59),
.B2(n_29),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_18),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_98),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_77),
.A2(n_26),
.B1(n_33),
.B2(n_29),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_94),
.B1(n_78),
.B2(n_67),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_63),
.A2(n_12),
.B1(n_11),
.B2(n_26),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_53),
.A2(n_29),
.B1(n_12),
.B2(n_11),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_53),
.A2(n_29),
.B(n_2),
.C(n_3),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_93),
.C(n_69),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_135),
.B(n_142),
.C(n_154),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_105),
.B(n_73),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_140),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_85),
.B1(n_71),
.B2(n_72),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_147),
.B1(n_148),
.B2(n_114),
.Y(n_176)
);

AO22x1_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_93),
.B1(n_71),
.B2(n_84),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_138),
.A2(n_152),
.B(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_76),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_60),
.C(n_57),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_151),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_95),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_155),
.Y(n_186)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_128),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_121),
.A2(n_94),
.B1(n_78),
.B2(n_67),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_54),
.B1(n_58),
.B2(n_68),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_164),
.B1(n_114),
.B2(n_104),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_106),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_66),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_75),
.C(n_58),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_75),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_0),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_169),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_0),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_0),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_159),
.B(n_165),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_128),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_167),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_59),
.B1(n_29),
.B2(n_5),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_3),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_89),
.C(n_88),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_103),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_104),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_107),
.B(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_3),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_170),
.B(n_171),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_4),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_111),
.B(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_181),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_176),
.A2(n_164),
.B1(n_202),
.B2(n_207),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_134),
.B1(n_118),
.B2(n_126),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_178),
.A2(n_187),
.B1(n_142),
.B2(n_135),
.Y(n_226)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_192),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_185),
.A2(n_114),
.B1(n_123),
.B2(n_163),
.Y(n_238)
);

AOI22x1_ASAP7_75t_L g187 ( 
.A1(n_138),
.A2(n_104),
.B1(n_134),
.B2(n_132),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_122),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_191),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_117),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_196),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_117),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_195),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_115),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_138),
.B(n_124),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_197),
.Y(n_218)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_198),
.B(n_202),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_115),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_201),
.Y(n_232)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_141),
.A2(n_131),
.B1(n_124),
.B2(n_108),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_140),
.B(n_136),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_151),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_159),
.C(n_157),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_152),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_211),
.A2(n_224),
.B(n_177),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_229),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_160),
.B1(n_150),
.B2(n_162),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_214),
.A2(n_205),
.B1(n_184),
.B2(n_179),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_139),
.B(n_154),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_210),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_162),
.B(n_147),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_176),
.A2(n_139),
.B1(n_154),
.B2(n_148),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_193),
.A2(n_158),
.B1(n_167),
.B2(n_156),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_178),
.A2(n_197),
.B1(n_196),
.B2(n_187),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_185),
.B1(n_195),
.B2(n_177),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_237),
.C(n_204),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_171),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_174),
.B1(n_181),
.B2(n_196),
.Y(n_243)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_244),
.C(n_246),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_233),
.B1(n_220),
.B2(n_232),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_208),
.C(n_186),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_245),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_186),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_252),
.B(n_253),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_249),
.A2(n_251),
.B1(n_216),
.B2(n_215),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_223),
.A2(n_209),
.B1(n_187),
.B2(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_200),
.C(n_191),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_259),
.C(n_219),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_256),
.B(n_231),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_233),
.A2(n_188),
.B(n_192),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_211),
.B(n_206),
.C(n_188),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_SL g278 ( 
.A(n_257),
.B(n_182),
.C(n_173),
.Y(n_278)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_258),
.A2(n_232),
.B1(n_222),
.B2(n_235),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_189),
.C(n_199),
.Y(n_259)
);

A2O1A1O1Ixp25_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_180),
.B(n_165),
.C(n_189),
.D(n_152),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_261),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_224),
.B1(n_220),
.B2(n_234),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_267),
.B1(n_279),
.B2(n_264),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_230),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_240),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_270),
.B(n_252),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_227),
.B1(n_249),
.B2(n_239),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_269),
.A2(n_273),
.B1(n_266),
.B2(n_268),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_248),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_216),
.B1(n_229),
.B2(n_231),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_247),
.A2(n_215),
.A3(n_222),
.B1(n_214),
.B2(n_236),
.C1(n_219),
.C2(n_228),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_277),
.C(n_103),
.Y(n_292)
);

NAND4xp25_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_260),
.C(n_261),
.D(n_253),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_247),
.A2(n_174),
.B1(n_163),
.B2(n_123),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_280),
.A2(n_284),
.B(n_290),
.Y(n_303)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_281),
.A2(n_288),
.B1(n_294),
.B2(n_212),
.Y(n_301)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_270),
.B(n_256),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_283),
.B(n_4),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_264),
.B(n_268),
.Y(n_285)
);

O2A1O1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_293),
.B(n_280),
.C(n_282),
.Y(n_306)
);

NAND4xp25_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_287),
.C(n_108),
.D(n_131),
.Y(n_300)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_262),
.A2(n_244),
.B1(n_250),
.B2(n_242),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_274),
.B1(n_275),
.B2(n_271),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_259),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_292),
.C(n_274),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_272),
.B(n_127),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_277),
.B1(n_269),
.B2(n_265),
.Y(n_295)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_293),
.C(n_5),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_294),
.A2(n_278),
.B1(n_271),
.B2(n_275),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_298),
.B(n_300),
.Y(n_307)
);

AOI21x1_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_175),
.B(n_212),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_283),
.B(n_285),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_304),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_289),
.B(n_88),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_291),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_6),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_299),
.A2(n_281),
.B1(n_286),
.B2(n_287),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_303),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_312),
.A2(n_313),
.B(n_316),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_290),
.B(n_292),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_314),
.A2(n_315),
.B(n_300),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_SL g315 ( 
.A(n_302),
.B(n_4),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_321),
.C(n_6),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_306),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_319),
.A2(n_322),
.B(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_305),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_297),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_314),
.B1(n_307),
.B2(n_295),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_326),
.Y(n_329)
);

AO21x1_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_309),
.B(n_298),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_320),
.B(n_7),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_325),
.B(n_7),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_329),
.B1(n_8),
.B2(n_9),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_6),
.Y(n_332)
);


endmodule