module fake_jpeg_142_n_110 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_110);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_16),
.B(n_4),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_5),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_40),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_7),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_20),
.A2(n_11),
.B(n_9),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_54),
.B(n_55),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_26),
.B(n_9),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_30),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_52),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_21),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_20),
.A2(n_28),
.B1(n_23),
.B2(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_23),
.B(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_22),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_36),
.A2(n_54),
.B1(n_46),
.B2(n_51),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_34),
.B1(n_67),
.B2(n_62),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_45),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_74),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_41),
.C(n_50),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_84),
.C(n_69),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_80),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_85),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_57),
.B1(n_72),
.B2(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_68),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_83),
.B1(n_74),
.B2(n_61),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_58),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_84),
.C(n_75),
.Y(n_94)
);

XNOR2x1_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_96),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_93),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_79),
.B1(n_66),
.B2(n_63),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_102),
.B(n_98),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_92),
.B1(n_88),
.B2(n_93),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_101),
.B(n_63),
.C(n_66),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_103),
.B(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_107),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_101),
.Y(n_110)
);


endmodule