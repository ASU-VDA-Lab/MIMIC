module fake_jpeg_29599_n_121 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_17),
.Y(n_47)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_6),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_21),
.B1(n_22),
.B2(n_15),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_59),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_17),
.B(n_22),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_44),
.B(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_12),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_20),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_46),
.B1(n_59),
.B2(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_70),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_12),
.B(n_15),
.C(n_0),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_51),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_0),
.Y(n_71)
);

NAND2x1_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_3),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_74),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_7),
.B1(n_8),
.B2(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_77),
.Y(n_83)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_60),
.B1(n_58),
.B2(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_58),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_63),
.Y(n_86)
);

AOI32xp33_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_53),
.A3(n_54),
.B1(n_51),
.B2(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_92),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_90),
.B(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_61),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_77),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_74),
.C(n_66),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_96),
.C(n_85),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_72),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_69),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_88),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_105),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_104),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_84),
.C(n_85),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_101),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_101),
.A2(n_90),
.B(n_83),
.C(n_98),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_98),
.B(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_113),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_109),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_91),
.C(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_115),
.B(n_110),
.Y(n_117)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_117),
.B1(n_91),
.B2(n_73),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_80),
.C(n_70),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_80),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_70),
.C(n_116),
.Y(n_121)
);


endmodule