module real_jpeg_13430_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_1),
.A2(n_33),
.B(n_47),
.C(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_1),
.B(n_71),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_1),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_1),
.A2(n_41),
.B(n_54),
.C(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_1),
.B(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_1),
.B(n_25),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_1),
.B(n_83),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_3),
.A2(n_35),
.B1(n_41),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_3),
.A2(n_22),
.B1(n_28),
.B2(n_61),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_5),
.A2(n_35),
.B1(n_41),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_59),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_5),
.A2(n_22),
.B1(n_28),
.B2(n_59),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_6),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_6),
.A2(n_27),
.B1(n_35),
.B2(n_41),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_10),
.A2(n_22),
.B1(n_28),
.B2(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_11),
.A2(n_35),
.B1(n_41),
.B2(n_44),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_11),
.A2(n_22),
.B1(n_28),
.B2(n_44),
.Y(n_116)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_13),
.A2(n_22),
.B1(n_28),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_88),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_86),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_62),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_17),
.B(n_62),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_42),
.C(n_50),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_18),
.B(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_31),
.B2(n_32),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_20),
.B(n_31),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_21),
.A2(n_25),
.B1(n_29),
.B2(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_21),
.A2(n_25),
.B1(n_26),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_21),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_21),
.A2(n_25),
.B1(n_38),
.B2(n_116),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_21),
.A2(n_25),
.B1(n_108),
.B2(n_116),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_22),
.A2(n_28),
.B1(n_54),
.B2(n_55),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_22),
.B(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_24),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_28),
.A2(n_38),
.B(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.A3(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_40),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_33),
.A2(n_34),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_42),
.B(n_50),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B(n_46),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_83),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_58),
.B1(n_83),
.B2(n_95),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_78),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_125),
.B(n_129),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_104),
.B(n_124),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_98),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_101),
.C(n_102),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_113),
.B(n_123),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_111),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_119),
.B(n_122),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_120),
.B(n_121),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_126),
.B(n_127),
.Y(n_129)
);


endmodule