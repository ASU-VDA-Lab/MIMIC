module fake_jpeg_8473_n_23 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_23);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_23;

wire n_13;
wire n_21;
wire n_10;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

AOI22xp33_ASAP7_75t_SL g10 ( 
.A1(n_7),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_3),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_11),
.B(n_13),
.Y(n_14)
);

AND2x6_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_15),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_0),
.C(n_1),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_8),
.Y(n_21)
);

BUFx24_ASAP7_75t_SL g22 ( 
.A(n_21),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_19),
.C(n_20),
.Y(n_23)
);


endmodule