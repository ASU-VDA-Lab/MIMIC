module fake_ariane_1168_n_1758 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1758);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1758;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_15),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_80),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_105),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_29),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_10),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_110),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_40),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_59),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_15),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_49),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_10),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_107),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_65),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_148),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_130),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_12),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_2),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_123),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_103),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_98),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_74),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_40),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_45),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_50),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_18),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_13),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_118),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_149),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_132),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_64),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_49),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_100),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_138),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_82),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_104),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_2),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_135),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_119),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_89),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_42),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_55),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_150),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_71),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_139),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_34),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_22),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_11),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_38),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_86),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_44),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_3),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_102),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_52),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_128),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_75),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_33),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_27),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_76),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_16),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_57),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_61),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_25),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_127),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_39),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_9),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_95),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_22),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_97),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_113),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_18),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_19),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_94),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_66),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_111),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_154),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_83),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_32),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_53),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_85),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_142),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_26),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_70),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_17),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_143),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_151),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_131),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_3),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_36),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_29),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_35),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_1),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_101),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_112),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_6),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_84),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_31),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_19),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_48),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_152),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_133),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_8),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_140),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_121),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_62),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_108),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_12),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_43),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_48),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_69),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_67),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_73),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_6),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_78),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_47),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_9),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_41),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_13),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_43),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_91),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_26),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_106),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_124),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_109),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_120),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_35),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_16),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_90),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_51),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_4),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_31),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_96),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_68),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_114),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_99),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_45),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_1),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_30),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_145),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_28),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_144),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_56),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_153),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_47),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_27),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_146),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_32),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_92),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_160),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_158),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_184),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_182),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_171),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_163),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_184),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_184),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_234),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_184),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_163),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_184),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_184),
.Y(n_326)
);

BUFx2_ASAP7_75t_SL g327 ( 
.A(n_202),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_184),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_167),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_248),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_277),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_184),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_215),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_293),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_215),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_215),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_296),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_215),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_215),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_225),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_225),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_167),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_250),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_162),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_186),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_202),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_194),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_237),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_237),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_229),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_211),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_214),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_229),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_232),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_212),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_232),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_235),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_292),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_213),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_171),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_222),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_235),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_297),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_228),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_297),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_230),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_247),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_169),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_193),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_233),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_187),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_199),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_205),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_236),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_202),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_292),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_210),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_216),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_247),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_223),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_284),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_231),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_254),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_243),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_193),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_262),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_251),
.Y(n_388)
);

INVxp33_ASAP7_75t_SL g389 ( 
.A(n_170),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_321),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_316),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_370),
.B(n_388),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_316),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_353),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_353),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_R g397 ( 
.A(n_347),
.B(n_189),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_361),
.B(n_284),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_320),
.A2(n_164),
.B(n_159),
.Y(n_400)
);

BUFx8_ASAP7_75t_L g401 ( 
.A(n_361),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_337),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_353),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_388),
.B(n_165),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_314),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_321),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_320),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_323),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_323),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_325),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_325),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_346),
.B(n_157),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_339),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_326),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_317),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_326),
.B(n_227),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_315),
.B(n_251),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_328),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_328),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_332),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_333),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_333),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_345),
.B(n_318),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_370),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_382),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_327),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_335),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_338),
.Y(n_433)
);

NAND2xp33_ASAP7_75t_R g434 ( 
.A(n_348),
.B(n_170),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_368),
.B(n_266),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_338),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_377),
.A2(n_178),
.B1(n_312),
.B2(n_291),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_330),
.A2(n_282),
.B1(n_312),
.B2(n_176),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_351),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_351),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_354),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_380),
.B(n_369),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_354),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_355),
.Y(n_444)
);

OA21x2_ASAP7_75t_L g445 ( 
.A1(n_355),
.A2(n_177),
.B(n_173),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_327),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_329),
.Y(n_447)
);

AND2x6_ASAP7_75t_L g448 ( 
.A(n_357),
.B(n_227),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_357),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_358),
.B(n_185),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_358),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_363),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_363),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_352),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_364),
.B(n_188),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_R g456 ( 
.A(n_356),
.B(n_176),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_364),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_343),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_376),
.A2(n_273),
.B1(n_178),
.B2(n_281),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_366),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_422),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_342),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_422),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_360),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_390),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_427),
.A2(n_389),
.B1(n_386),
.B2(n_263),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_431),
.A2(n_291),
.B1(n_273),
.B2(n_183),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_390),
.Y(n_470)
);

AOI21x1_ASAP7_75t_L g471 ( 
.A1(n_391),
.A2(n_366),
.B(n_206),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_427),
.B(n_369),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_420),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_390),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_446),
.B(n_362),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_432),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_359),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_407),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_446),
.B(n_365),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_401),
.B(n_322),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_420),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_436),
.Y(n_483)
);

INVxp33_ASAP7_75t_L g484 ( 
.A(n_438),
.Y(n_484)
);

OAI22xp33_ASAP7_75t_L g485 ( 
.A1(n_459),
.A2(n_344),
.B1(n_319),
.B2(n_324),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_407),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_407),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_407),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_436),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_407),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_397),
.B(n_367),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_391),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_407),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_428),
.B(n_371),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_425),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_447),
.B(n_331),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_425),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_437),
.B(n_334),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_425),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_393),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_426),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_426),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_415),
.B(n_375),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_409),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_428),
.B(n_385),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_406),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_428),
.B(n_372),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_419),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_437),
.A2(n_281),
.B1(n_183),
.B2(n_286),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_442),
.B(n_157),
.Y(n_512)
);

BUFx4f_ASAP7_75t_L g513 ( 
.A(n_419),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_428),
.B(n_372),
.Y(n_514)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_409),
.B(n_413),
.C(n_410),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_410),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_435),
.B(n_442),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_435),
.B(n_373),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_435),
.B(n_373),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_426),
.Y(n_520)
);

AO21x2_ASAP7_75t_L g521 ( 
.A1(n_413),
.A2(n_417),
.B(n_414),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_429),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_392),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_414),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_417),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_405),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_435),
.B(n_374),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_442),
.B(n_374),
.Y(n_529)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_454),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_406),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_443),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_421),
.Y(n_533)
);

NOR2x1p5_ASAP7_75t_L g534 ( 
.A(n_434),
.B(n_282),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_421),
.Y(n_535)
);

OAI22xp33_ASAP7_75t_L g536 ( 
.A1(n_459),
.A2(n_309),
.B1(n_286),
.B2(n_272),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_429),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_423),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_423),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_419),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_454),
.B(n_161),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_420),
.B(n_378),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_438),
.B(n_378),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_424),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_430),
.B(n_379),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_424),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_408),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_443),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_406),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_443),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_392),
.B(n_379),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_443),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_418),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_445),
.A2(n_278),
.B1(n_274),
.B2(n_280),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_443),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_408),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_443),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_430),
.B(n_381),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_399),
.B(n_161),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_443),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_L g561 ( 
.A1(n_456),
.A2(n_309),
.B1(n_249),
.B2(n_256),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_419),
.B(n_168),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_460),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_399),
.B(n_381),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_460),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_460),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_408),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_460),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_411),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_460),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g571 ( 
.A1(n_430),
.A2(n_257),
.B1(n_302),
.B2(n_303),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_460),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_392),
.B(n_383),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_392),
.B(n_383),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_439),
.B(n_168),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_460),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_445),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_402),
.Y(n_578)
);

AND3x2_ASAP7_75t_L g579 ( 
.A(n_458),
.B(n_264),
.C(n_301),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_439),
.B(n_172),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_406),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_453),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_406),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_439),
.B(n_172),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_445),
.A2(n_283),
.B1(n_267),
.B2(n_295),
.Y(n_585)
);

OAI22x1_ASAP7_75t_L g586 ( 
.A1(n_458),
.A2(n_260),
.B1(n_255),
.B2(n_253),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_406),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_406),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_453),
.Y(n_589)
);

AO21x2_ASAP7_75t_L g590 ( 
.A1(n_404),
.A2(n_290),
.B(n_201),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_453),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_457),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_439),
.B(n_384),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_411),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_445),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_411),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_416),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_457),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_457),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_433),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_404),
.B(n_384),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_445),
.A2(n_310),
.B1(n_305),
.B2(n_387),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_416),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_416),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_433),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_433),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_448),
.A2(n_387),
.B1(n_166),
.B2(n_313),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_433),
.Y(n_608)
);

OAI22xp33_ASAP7_75t_L g609 ( 
.A1(n_450),
.A2(n_350),
.B1(n_349),
.B2(n_341),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_433),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_484),
.A2(n_448),
.B1(n_419),
.B2(n_400),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_477),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_513),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_473),
.B(n_440),
.Y(n_614)
);

OAI22x1_ASAP7_75t_R g615 ( 
.A1(n_526),
.A2(n_401),
.B1(n_341),
.B2(n_349),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_466),
.B(n_440),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_518),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_538),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_475),
.B(n_419),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_473),
.B(n_419),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_482),
.B(n_419),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_498),
.B(n_441),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_463),
.B(n_401),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_482),
.A2(n_448),
.B1(n_452),
.B2(n_451),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_498),
.B(n_472),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_517),
.B(n_472),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_593),
.B(n_441),
.Y(n_627)
);

INVxp33_ASAP7_75t_L g628 ( 
.A(n_478),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_480),
.B(n_444),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_593),
.B(n_545),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_558),
.B(n_444),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_559),
.B(n_449),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_539),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_526),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_530),
.B(n_401),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_512),
.B(n_449),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_601),
.B(n_451),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_601),
.B(n_452),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_601),
.B(n_448),
.Y(n_639)
);

OAI221xp5_ASAP7_75t_L g640 ( 
.A1(n_511),
.A2(n_455),
.B1(n_450),
.B2(n_340),
.C(n_350),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_530),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_530),
.B(n_174),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_553),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_553),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_601),
.B(n_448),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_530),
.Y(n_646)
);

BUFx6f_ASAP7_75t_SL g647 ( 
.A(n_543),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_478),
.B(n_455),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_601),
.B(n_448),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_519),
.B(n_528),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_523),
.B(n_203),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_539),
.Y(n_652)
);

BUFx5_ASAP7_75t_L g653 ( 
.A(n_587),
.Y(n_653)
);

NAND3xp33_ASAP7_75t_L g654 ( 
.A(n_511),
.B(n_469),
.C(n_496),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_513),
.B(n_174),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_542),
.B(n_448),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_564),
.B(n_340),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_523),
.B(n_306),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_R g659 ( 
.A(n_578),
.B(n_175),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_574),
.B(n_448),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_529),
.B(n_448),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_513),
.B(n_465),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_564),
.B(n_400),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_546),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_546),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_483),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_465),
.B(n_175),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_507),
.B(n_400),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_543),
.B(n_400),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_483),
.Y(n_670)
);

NOR3xp33_ASAP7_75t_L g671 ( 
.A(n_536),
.B(n_217),
.C(n_245),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_578),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_509),
.B(n_400),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_465),
.B(n_179),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_547),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_468),
.B(n_500),
.Y(n_676)
);

OAI22xp33_ASAP7_75t_L g677 ( 
.A1(n_543),
.A2(n_166),
.B1(n_313),
.B2(n_180),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_534),
.A2(n_181),
.B1(n_180),
.B2(n_311),
.Y(n_678)
);

NAND2x1_ASAP7_75t_L g679 ( 
.A(n_465),
.B(n_394),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_489),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_554),
.A2(n_266),
.B1(n_294),
.B2(n_412),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_L g682 ( 
.A(n_492),
.B(n_181),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_500),
.B(n_412),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_573),
.Y(n_684)
);

AND2x6_ASAP7_75t_L g685 ( 
.A(n_607),
.B(n_227),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_531),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_540),
.B(n_275),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_489),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_SL g689 ( 
.A1(n_543),
.A2(n_275),
.B1(n_276),
.B2(n_287),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_531),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_L g691 ( 
.A(n_492),
.B(n_276),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_494),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_514),
.B(n_412),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_540),
.B(n_287),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_585),
.A2(n_294),
.B1(n_412),
.B2(n_433),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_494),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_547),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_540),
.B(n_288),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_543),
.A2(n_289),
.B1(n_311),
.B2(n_308),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_505),
.B(n_288),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_556),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_573),
.B(n_289),
.Y(n_702)
);

AO22x2_ASAP7_75t_L g703 ( 
.A1(n_577),
.A2(n_220),
.B1(n_221),
.B2(n_226),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_461),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_502),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_541),
.B(n_308),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_502),
.B(n_190),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_575),
.B(n_238),
.Y(n_708)
);

INVx8_ASAP7_75t_L g709 ( 
.A(n_531),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_531),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_506),
.A2(n_544),
.B1(n_535),
.B2(n_533),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_506),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_516),
.B(n_191),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_516),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_524),
.B(n_269),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_579),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_524),
.A2(n_300),
.B(n_252),
.C(n_268),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_525),
.B(n_192),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_525),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_551),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_533),
.B(n_535),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_L g722 ( 
.A(n_544),
.B(n_269),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_590),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_515),
.A2(n_285),
.B(n_299),
.C(n_242),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_607),
.A2(n_279),
.B1(n_304),
.B2(n_307),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_540),
.B(n_195),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_470),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_510),
.B(n_196),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_470),
.B(n_197),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_474),
.B(n_198),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_474),
.B(n_200),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_510),
.B(n_204),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_485),
.B(n_0),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_582),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_481),
.B(n_433),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_510),
.B(n_207),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_580),
.B(n_0),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_556),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_567),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_467),
.B(n_208),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_467),
.B(n_209),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_476),
.B(n_259),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_571),
.B(n_561),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_567),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_590),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_476),
.B(n_261),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_584),
.B(n_4),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_462),
.B(n_258),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_L g749 ( 
.A(n_515),
.B(n_600),
.Y(n_749)
);

OAI22xp33_ASAP7_75t_L g750 ( 
.A1(n_586),
.A2(n_244),
.B1(n_218),
.B2(n_219),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_462),
.B(n_224),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_491),
.B(n_5),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_582),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_488),
.B(n_239),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_569),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_589),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_586),
.B(n_5),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_464),
.B(n_270),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_609),
.B(n_271),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_521),
.B(n_7),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_488),
.B(n_7),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_531),
.B(n_240),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_464),
.B(n_298),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_569),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_589),
.B(n_241),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_591),
.B(n_265),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_594),
.Y(n_767)
);

BUFx5_ASAP7_75t_L g768 ( 
.A(n_587),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_549),
.B(n_246),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_591),
.B(n_403),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_592),
.B(n_403),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_488),
.B(n_8),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_592),
.B(n_403),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_602),
.B(n_11),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_594),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_590),
.B(n_14),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_596),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_598),
.B(n_394),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_612),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_628),
.B(n_495),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_676),
.A2(n_599),
.B1(n_598),
.B2(n_461),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_634),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_617),
.B(n_549),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_L g784 ( 
.A(n_654),
.B(n_562),
.C(n_599),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_634),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_671),
.A2(n_521),
.B1(n_532),
.B2(n_572),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_709),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_617),
.B(n_495),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_704),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_704),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_616),
.B(n_521),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_644),
.Y(n_792)
);

O2A1O1Ixp5_ASAP7_75t_L g793 ( 
.A1(n_668),
.A2(n_471),
.B(n_486),
.C(n_493),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_619),
.B(n_495),
.Y(n_794)
);

NAND2x1p5_ASAP7_75t_L g795 ( 
.A(n_613),
.B(n_532),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_641),
.B(n_549),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_672),
.B(n_577),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_616),
.B(n_595),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_613),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_666),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_648),
.B(n_581),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_709),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_709),
.Y(n_803)
);

OR2x6_ASAP7_75t_L g804 ( 
.A(n_643),
.B(n_595),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_613),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_675),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_657),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_697),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_625),
.B(n_497),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_659),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_626),
.B(n_497),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_622),
.B(n_499),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_684),
.B(n_499),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_650),
.B(n_501),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_630),
.B(n_501),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_774),
.A2(n_537),
.B1(n_503),
.B2(n_504),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_683),
.Y(n_817)
);

AND2x6_ASAP7_75t_SL g818 ( 
.A(n_752),
.B(n_548),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_670),
.B(n_680),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_688),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_743),
.B(n_581),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_643),
.B(n_503),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_692),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_646),
.B(n_549),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_615),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_696),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_635),
.B(n_532),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_705),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_712),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_714),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_719),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_727),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_721),
.B(n_504),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_734),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_701),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_720),
.B(n_520),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_720),
.B(n_520),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_753),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_756),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_647),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_677),
.B(n_613),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_647),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_627),
.B(n_522),
.Y(n_843)
);

NAND2x1p5_ASAP7_75t_L g844 ( 
.A(n_760),
.B(n_550),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_677),
.B(n_549),
.Y(n_845)
);

OR2x4_ASAP7_75t_L g846 ( 
.A(n_706),
.B(n_548),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_711),
.B(n_522),
.Y(n_847)
);

INVx5_ASAP7_75t_L g848 ( 
.A(n_686),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_663),
.B(n_527),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_738),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_739),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_631),
.B(n_527),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_671),
.A2(n_537),
.B1(n_596),
.B2(n_597),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_623),
.B(n_550),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_744),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_733),
.B(n_604),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_614),
.B(n_581),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_614),
.B(n_583),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_661),
.B(n_583),
.Y(n_859)
);

INVx5_ASAP7_75t_L g860 ( 
.A(n_686),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_651),
.B(n_604),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_699),
.A2(n_572),
.B1(n_550),
.B2(n_570),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_618),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_752),
.B(n_600),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_629),
.B(n_600),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_633),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_669),
.B(n_572),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_668),
.B(n_583),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_706),
.B(n_588),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_652),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_664),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_636),
.B(n_588),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_665),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_636),
.B(n_588),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_656),
.B(n_479),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_637),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_638),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_716),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_735),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_755),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_673),
.A2(n_508),
.B(n_479),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_629),
.B(n_600),
.Y(n_882)
);

NOR2x1p5_ASAP7_75t_L g883 ( 
.A(n_757),
.B(n_702),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_686),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_760),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_764),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_767),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_632),
.B(n_486),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_700),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_632),
.B(n_493),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_686),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_690),
.Y(n_892)
);

AOI221xp5_ASAP7_75t_SL g893 ( 
.A1(n_640),
.A2(n_566),
.B1(n_563),
.B2(n_565),
.C(n_560),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_703),
.A2(n_597),
.B1(n_603),
.B2(n_576),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_775),
.B(n_490),
.Y(n_895)
);

CKINVDCx11_ASAP7_75t_R g896 ( 
.A(n_669),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_700),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_737),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_651),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_690),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_689),
.B(n_600),
.Y(n_901)
);

OAI22xp33_ASAP7_75t_L g902 ( 
.A1(n_678),
.A2(n_563),
.B1(n_557),
.B2(n_560),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_777),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_770),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_658),
.B(n_669),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_658),
.B(n_490),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_737),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_660),
.B(n_487),
.Y(n_908)
);

O2A1O1Ixp5_ASAP7_75t_L g909 ( 
.A1(n_761),
.A2(n_487),
.B(n_565),
.C(n_552),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_747),
.A2(n_557),
.B1(n_552),
.B2(n_555),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_771),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_642),
.B(n_605),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_723),
.B(n_568),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_776),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_747),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_690),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_690),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_749),
.A2(n_693),
.B(n_621),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_708),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_639),
.B(n_605),
.Y(n_920)
);

AO22x1_ASAP7_75t_L g921 ( 
.A1(n_685),
.A2(n_570),
.B1(n_566),
.B2(n_568),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_708),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_750),
.B(n_576),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_645),
.B(n_610),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_710),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_SL g926 ( 
.A1(n_611),
.A2(n_214),
.B1(n_608),
.B2(n_606),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_SL g927 ( 
.A(n_717),
.B(n_610),
.C(n_608),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_745),
.B(n_603),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_710),
.Y(n_929)
);

NAND2x1p5_ASAP7_75t_L g930 ( 
.A(n_710),
.B(n_606),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_649),
.B(n_269),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_773),
.Y(n_932)
);

NOR3xp33_ASAP7_75t_SL g933 ( 
.A(n_761),
.B(n_14),
.C(n_17),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_620),
.B(n_394),
.Y(n_934)
);

BUFx4f_ASAP7_75t_L g935 ( 
.A(n_685),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_778),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_681),
.B(n_20),
.Y(n_937)
);

NOR3xp33_ASAP7_75t_SL g938 ( 
.A(n_772),
.B(n_20),
.C(n_21),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_707),
.B(n_269),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_703),
.A2(n_214),
.B1(n_269),
.B2(n_396),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_748),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_710),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_751),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_611),
.B(n_396),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_772),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_758),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_662),
.B(n_398),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_763),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_765),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_653),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_L g951 ( 
.A(n_653),
.B(n_768),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_624),
.B(n_396),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_703),
.A2(n_685),
.B1(n_725),
.B2(n_681),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_653),
.B(n_768),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_685),
.A2(n_214),
.B1(n_269),
.B2(n_395),
.Y(n_955)
);

OR2x2_ASAP7_75t_SL g956 ( 
.A(n_713),
.B(n_214),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_766),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_718),
.B(n_269),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_740),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_682),
.B(n_21),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_685),
.B(n_23),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_653),
.B(n_768),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_741),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_679),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_691),
.A2(n_269),
.B1(n_395),
.B2(n_398),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_899),
.B(n_725),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_806),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_779),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_885),
.B(n_844),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_919),
.B(n_759),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_SL g971 ( 
.A1(n_788),
.A2(n_754),
.B(n_730),
.C(n_731),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_915),
.A2(n_729),
.B(n_724),
.C(n_746),
.Y(n_972)
);

OR2x6_ASAP7_75t_L g973 ( 
.A(n_844),
.B(n_655),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_922),
.B(n_695),
.Y(n_974)
);

INVx5_ASAP7_75t_L g975 ( 
.A(n_787),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_807),
.B(n_856),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_953),
.A2(n_695),
.B1(n_674),
.B2(n_687),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_933),
.A2(n_742),
.B(n_694),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_787),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_787),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_802),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_821),
.A2(n_722),
.B(n_715),
.C(n_698),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_889),
.B(n_653),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_897),
.B(n_653),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_937),
.A2(n_667),
.B1(n_762),
.B2(n_769),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_898),
.A2(n_726),
.B(n_736),
.C(n_732),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_802),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_822),
.B(n_728),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_798),
.A2(n_768),
.B(n_398),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_808),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_941),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_802),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_943),
.A2(n_946),
.B(n_949),
.C(n_948),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_907),
.B(n_810),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_957),
.A2(n_24),
.B(n_28),
.C(n_30),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_792),
.B(n_768),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_798),
.A2(n_768),
.B(n_398),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_835),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_878),
.Y(n_999)
);

AND3x1_ASAP7_75t_SL g1000 ( 
.A(n_883),
.B(n_33),
.C(n_34),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_868),
.A2(n_791),
.B(n_864),
.Y(n_1001)
);

OAI21xp33_ASAP7_75t_SL g1002 ( 
.A1(n_819),
.A2(n_791),
.B(n_847),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_945),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_793),
.A2(n_398),
.B(n_39),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_868),
.A2(n_398),
.B(n_395),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_812),
.B(n_37),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_951),
.A2(n_398),
.B(n_395),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_850),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_809),
.B(n_41),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_800),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_782),
.B(n_42),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_785),
.B(n_44),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_954),
.A2(n_395),
.B(n_54),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_959),
.A2(n_46),
.B(n_395),
.C(n_60),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_954),
.A2(n_395),
.B(n_58),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_817),
.B(n_46),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_819),
.A2(n_63),
.B1(n_72),
.B2(n_77),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_820),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_926),
.A2(n_79),
.B1(n_81),
.B2(n_87),
.Y(n_1019)
);

NOR2xp67_ASAP7_75t_SL g1020 ( 
.A(n_803),
.B(n_88),
.Y(n_1020)
);

OAI21xp33_ASAP7_75t_SL g1021 ( 
.A1(n_847),
.A2(n_126),
.B(n_136),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_963),
.A2(n_137),
.B(n_141),
.C(n_156),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_938),
.A2(n_801),
.B(n_822),
.C(n_960),
.Y(n_1023)
);

NOR3xp33_ASAP7_75t_L g1024 ( 
.A(n_902),
.B(n_901),
.C(n_841),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_823),
.Y(n_1025)
);

BUFx2_ASAP7_75t_SL g1026 ( 
.A(n_961),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_826),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_876),
.B(n_877),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_962),
.A2(n_852),
.B(n_794),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_935),
.A2(n_831),
.B1(n_829),
.B2(n_830),
.Y(n_1030)
);

OA21x2_ASAP7_75t_L g1031 ( 
.A1(n_909),
.A2(n_793),
.B(n_881),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_840),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_SL g1033 ( 
.A(n_842),
.B(n_828),
.C(n_780),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_825),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_846),
.B(n_818),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_797),
.Y(n_1036)
);

AND2x4_ASAP7_75t_SL g1037 ( 
.A(n_803),
.B(n_797),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_803),
.B(n_935),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_852),
.A2(n_833),
.B(n_843),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_822),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_861),
.B(n_836),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_851),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_833),
.A2(n_843),
.B(n_918),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_834),
.A2(n_838),
.B1(n_839),
.B2(n_846),
.Y(n_1044)
);

AO32x2_ASAP7_75t_L g1045 ( 
.A1(n_879),
.A2(n_891),
.A3(n_942),
.B1(n_893),
.B2(n_909),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_918),
.A2(n_814),
.B(n_869),
.Y(n_1046)
);

AO21x1_ASAP7_75t_L g1047 ( 
.A1(n_923),
.A2(n_905),
.B(n_845),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_914),
.B(n_813),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_814),
.A2(n_815),
.B(n_859),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_912),
.A2(n_786),
.B(n_784),
.C(n_872),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_836),
.B(n_837),
.Y(n_1051)
);

AOI21x1_ASAP7_75t_L g1052 ( 
.A1(n_881),
.A2(n_958),
.B(n_939),
.Y(n_1052)
);

BUFx12f_ASAP7_75t_L g1053 ( 
.A(n_896),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_815),
.A2(n_859),
.B(n_908),
.Y(n_1054)
);

O2A1O1Ixp5_ASAP7_75t_L g1055 ( 
.A1(n_783),
.A2(n_865),
.B(n_882),
.C(n_824),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_837),
.B(n_832),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_904),
.B(n_932),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_804),
.A2(n_874),
.B(n_858),
.C(n_857),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_884),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_936),
.B(n_811),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_855),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_908),
.A2(n_849),
.B(n_875),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_849),
.A2(n_875),
.B(n_811),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_886),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_797),
.B(n_804),
.Y(n_1065)
);

O2A1O1Ixp5_ASAP7_75t_L g1066 ( 
.A1(n_796),
.A2(n_931),
.B(n_906),
.C(n_950),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_867),
.B(n_860),
.Y(n_1067)
);

O2A1O1Ixp5_ASAP7_75t_L g1068 ( 
.A1(n_921),
.A2(n_942),
.B(n_891),
.C(n_892),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_R g1069 ( 
.A(n_848),
.B(n_860),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_854),
.B(n_789),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_884),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_888),
.A2(n_890),
.B(n_910),
.C(n_854),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_863),
.B(n_866),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_961),
.A2(n_781),
.B1(n_858),
.B2(n_940),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_911),
.B(n_890),
.Y(n_1075)
);

OAI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_888),
.A2(n_862),
.B(n_853),
.Y(n_1076)
);

O2A1O1Ixp5_ASAP7_75t_L g1077 ( 
.A1(n_892),
.A2(n_900),
.B(n_827),
.C(n_952),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_929),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_934),
.A2(n_895),
.B(n_913),
.Y(n_1079)
);

AO32x2_ASAP7_75t_L g1080 ( 
.A1(n_956),
.A2(n_927),
.A3(n_894),
.B1(n_944),
.B2(n_913),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_870),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_867),
.B(n_848),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_790),
.A2(n_927),
.B(n_920),
.C(n_827),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_920),
.A2(n_799),
.B(n_805),
.C(n_952),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_871),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_873),
.B(n_900),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_880),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_887),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_799),
.A2(n_805),
.B(n_965),
.C(n_955),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_903),
.Y(n_1090)
);

INVx4_ASAP7_75t_L g1091 ( 
.A(n_884),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_924),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_934),
.A2(n_795),
.B(n_924),
.C(n_895),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_795),
.A2(n_924),
.B(n_930),
.C(n_947),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_816),
.B(n_916),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_928),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_930),
.A2(n_944),
.B(n_928),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_916),
.B(n_917),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_916),
.A2(n_917),
.B(n_925),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_917),
.B(n_925),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_925),
.B(n_964),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_964),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_964),
.A2(n_654),
.B(n_821),
.C(n_747),
.Y(n_1103)
);

O2A1O1Ixp5_ASAP7_75t_L g1104 ( 
.A1(n_947),
.A2(n_939),
.B(n_958),
.C(n_909),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_798),
.A2(n_868),
.B(n_951),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_779),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_899),
.B(n_625),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_806),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_787),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_806),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_919),
.B(n_899),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_1067),
.B(n_1082),
.Y(n_1113)
);

NOR2x1_ASAP7_75t_SL g1114 ( 
.A(n_996),
.B(n_1026),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_966),
.B(n_1107),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1105),
.A2(n_1046),
.B(n_1039),
.Y(n_1116)
);

INVx8_ASAP7_75t_L g1117 ( 
.A(n_975),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1067),
.B(n_1082),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1029),
.A2(n_1043),
.B(n_1002),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1052),
.A2(n_1097),
.B(n_1062),
.Y(n_1120)
);

OA21x2_ASAP7_75t_L g1121 ( 
.A1(n_1004),
.A2(n_1050),
.B(n_1047),
.Y(n_1121)
);

AOI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1001),
.A2(n_1079),
.B(n_1054),
.Y(n_1122)
);

NAND2xp33_ASAP7_75t_R g1123 ( 
.A(n_1069),
.B(n_1033),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1041),
.B(n_1075),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1056),
.A2(n_970),
.B1(n_1103),
.B2(n_1057),
.Y(n_1125)
);

AO31x2_ASAP7_75t_L g1126 ( 
.A1(n_1063),
.A2(n_1049),
.A3(n_1072),
.B(n_1044),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1028),
.B(n_1096),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1005),
.A2(n_1104),
.B(n_989),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1073),
.Y(n_1129)
);

AOI31xp67_ASAP7_75t_L g1130 ( 
.A1(n_1102),
.A2(n_983),
.A3(n_984),
.B(n_988),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_1034),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1091),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1111),
.B(n_976),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_997),
.A2(n_1093),
.B(n_1015),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_1035),
.B(n_994),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1013),
.A2(n_1004),
.B(n_1066),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1007),
.A2(n_1094),
.B(n_1030),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_969),
.B(n_1040),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_975),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1048),
.B(n_1011),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_1012),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1076),
.A2(n_982),
.B(n_1058),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1031),
.A2(n_1055),
.B(n_1083),
.Y(n_1143)
);

BUFx10_ASAP7_75t_L g1144 ( 
.A(n_980),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1078),
.B(n_993),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1068),
.A2(n_1077),
.B(n_1099),
.Y(n_1146)
);

NAND2xp33_ASAP7_75t_L g1147 ( 
.A(n_978),
.B(n_1059),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1076),
.B(n_974),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1010),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_972),
.A2(n_986),
.B(n_977),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1095),
.A2(n_1065),
.B(n_1014),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1032),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_977),
.A2(n_1074),
.A3(n_1019),
.B(n_1084),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1023),
.B(n_975),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1022),
.A2(n_1098),
.B(n_1100),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_978),
.A2(n_1021),
.B(n_1024),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_999),
.B(n_1070),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1074),
.A2(n_1019),
.A3(n_1089),
.B(n_1017),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1018),
.B(n_1106),
.Y(n_1159)
);

CKINVDCx11_ASAP7_75t_R g1160 ( 
.A(n_1053),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_988),
.B(n_1059),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_SL g1162 ( 
.A(n_1003),
.B(n_991),
.C(n_995),
.Y(n_1162)
);

NOR4xp25_ASAP7_75t_L g1163 ( 
.A(n_1006),
.B(n_1009),
.C(n_1027),
.D(n_1025),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1059),
.B(n_1071),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_967),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_985),
.A2(n_1038),
.B(n_1036),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_969),
.B(n_1081),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1092),
.A2(n_1087),
.B(n_1085),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_971),
.A2(n_996),
.B(n_1101),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1086),
.A2(n_1110),
.A3(n_1042),
.B(n_1108),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1016),
.A2(n_1008),
.B(n_1090),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_990),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_998),
.A2(n_1061),
.B(n_1064),
.Y(n_1173)
);

OA21x2_ASAP7_75t_L g1174 ( 
.A1(n_1045),
.A2(n_1088),
.B(n_1080),
.Y(n_1174)
);

NOR2xp67_ASAP7_75t_SL g1175 ( 
.A(n_980),
.B(n_981),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_979),
.A2(n_1109),
.B(n_992),
.Y(n_1176)
);

NAND3xp33_ASAP7_75t_SL g1177 ( 
.A(n_1000),
.B(n_1091),
.C(n_996),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1037),
.A2(n_992),
.B(n_1109),
.C(n_979),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_969),
.B(n_1071),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_973),
.A2(n_1071),
.B(n_1045),
.Y(n_1180)
);

BUFx4_ASAP7_75t_SL g1181 ( 
.A(n_973),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_973),
.A2(n_1045),
.B(n_987),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_987),
.A2(n_980),
.B(n_981),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_981),
.B(n_1080),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1080),
.B(n_1020),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_975),
.Y(n_1186)
);

OR2x6_ASAP7_75t_L g1187 ( 
.A(n_1026),
.B(n_885),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1043),
.A2(n_1052),
.B(n_1029),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_976),
.B(n_625),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_976),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1047),
.A2(n_1062),
.A3(n_1063),
.B(n_1097),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_976),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1105),
.A2(n_951),
.B(n_1046),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1046),
.A2(n_1052),
.B(n_1043),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1067),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1067),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_976),
.B(n_625),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_1111),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1050),
.A2(n_791),
.B(n_1072),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_976),
.B(n_625),
.Y(n_1204)
);

AO32x2_ASAP7_75t_L g1205 ( 
.A1(n_1044),
.A2(n_1030),
.A3(n_1074),
.B1(n_1019),
.B2(n_926),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1043),
.A2(n_1052),
.B(n_1029),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1207)
);

NAND2x1_ASAP7_75t_L g1208 ( 
.A(n_996),
.B(n_891),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_976),
.B(n_625),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1043),
.A2(n_1052),
.B(n_1029),
.Y(n_1210)
);

OAI22x1_ASAP7_75t_L g1211 ( 
.A1(n_1035),
.A2(n_919),
.B1(n_699),
.B2(n_459),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1041),
.A2(n_953),
.B1(n_654),
.B2(n_919),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_1111),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1214)
);

NOR2xp67_ASAP7_75t_L g1215 ( 
.A(n_975),
.B(n_810),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1043),
.A2(n_1052),
.B(n_1029),
.Y(n_1216)
);

NOR2x1_ASAP7_75t_L g1217 ( 
.A(n_1032),
.B(n_644),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_976),
.Y(n_1218)
);

AOI221x1_ASAP7_75t_L g1219 ( 
.A1(n_1024),
.A2(n_1019),
.B1(n_703),
.B2(n_1103),
.C(n_1004),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_968),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_976),
.Y(n_1221)
);

INVx5_ASAP7_75t_L g1222 ( 
.A(n_996),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1032),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1105),
.A2(n_951),
.B(n_1046),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1034),
.Y(n_1225)
);

INVx3_ASAP7_75t_SL g1226 ( 
.A(n_1034),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1041),
.A2(n_953),
.B1(n_654),
.B2(n_919),
.Y(n_1227)
);

BUFx2_ASAP7_75t_R g1228 ( 
.A(n_1034),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1105),
.A2(n_951),
.B(n_1046),
.Y(n_1229)
);

AOI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1046),
.A2(n_1052),
.B(n_1043),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_SL g1231 ( 
.A1(n_1030),
.A2(n_1023),
.B(n_1044),
.Y(n_1231)
);

AND2x6_ASAP7_75t_L g1232 ( 
.A(n_1067),
.B(n_961),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1233)
);

AOI221x1_ASAP7_75t_L g1234 ( 
.A1(n_1024),
.A2(n_1019),
.B1(n_703),
.B2(n_1103),
.C(n_1004),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1051),
.B(n_1060),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1067),
.B(n_1082),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1046),
.A2(n_1052),
.B(n_1043),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_966),
.B(n_1107),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1111),
.B(n_919),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1067),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_968),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1067),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1032),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1050),
.A2(n_791),
.B(n_1072),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1002),
.A2(n_654),
.B(n_907),
.C(n_898),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1043),
.A2(n_1052),
.B(n_1029),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1032),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1043),
.A2(n_1052),
.B(n_1029),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_976),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1050),
.A2(n_791),
.B(n_1072),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1047),
.A2(n_1062),
.A3(n_1063),
.B(n_1097),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1111),
.B(n_919),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_968),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_SL g1254 ( 
.A1(n_1019),
.A2(n_1072),
.B(n_1030),
.Y(n_1254)
);

BUFx2_ASAP7_75t_R g1255 ( 
.A(n_1131),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1245),
.A2(n_1156),
.B(n_1125),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1159),
.Y(n_1257)
);

NAND3xp33_ASAP7_75t_L g1258 ( 
.A(n_1150),
.B(n_1156),
.C(n_1125),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1189),
.B(n_1201),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1141),
.A2(n_1254),
.B1(n_1213),
.B2(n_1202),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1115),
.B(n_1238),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1212),
.A2(n_1227),
.B1(n_1150),
.B2(n_1211),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1212),
.A2(n_1227),
.B1(n_1162),
.B2(n_1250),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1170),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1117),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1124),
.B(n_1112),
.Y(n_1266)
);

OAI221xp5_ASAP7_75t_L g1267 ( 
.A1(n_1163),
.A2(n_1140),
.B1(n_1145),
.B2(n_1142),
.C(n_1252),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1159),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1170),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_1160),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1225),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1223),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1228),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1237),
.A2(n_1206),
.B(n_1188),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1218),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1226),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1152),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1117),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1190),
.B(n_1192),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1119),
.A2(n_1116),
.B(n_1248),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1190),
.B(n_1192),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1219),
.A2(n_1234),
.B(n_1142),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1149),
.Y(n_1283)
);

BUFx2_ASAP7_75t_SL g1284 ( 
.A(n_1215),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1170),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1221),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1210),
.A2(n_1216),
.B(n_1246),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1249),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1203),
.A2(n_1250),
.B1(n_1244),
.B2(n_1231),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1133),
.B(n_1239),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1203),
.A2(n_1244),
.B1(n_1121),
.B2(n_1204),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1147),
.A2(n_1154),
.B(n_1163),
.C(n_1135),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1222),
.B(n_1113),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1120),
.A2(n_1229),
.B(n_1224),
.Y(n_1294)
);

OAI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1194),
.A2(n_1214),
.B1(n_1207),
.B2(n_1199),
.Y(n_1295)
);

BUFx8_ASAP7_75t_L g1296 ( 
.A(n_1209),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1194),
.A2(n_1235),
.B(n_1199),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1148),
.A2(n_1182),
.A3(n_1196),
.B(n_1180),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1220),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1134),
.A2(n_1122),
.B(n_1136),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1207),
.B(n_1214),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1233),
.A2(n_1235),
.B(n_1169),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1191),
.Y(n_1303)
);

INVx4_ASAP7_75t_L g1304 ( 
.A(n_1139),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1123),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1146),
.A2(n_1143),
.B(n_1137),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1233),
.B(n_1127),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1174),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1193),
.Y(n_1309)
);

NOR2x1_ASAP7_75t_L g1310 ( 
.A(n_1177),
.B(n_1186),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1155),
.A2(n_1151),
.B(n_1168),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1195),
.B(n_1157),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1148),
.A2(n_1185),
.B(n_1127),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1171),
.A2(n_1208),
.B(n_1166),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1121),
.A2(n_1164),
.B(n_1130),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1232),
.A2(n_1187),
.B1(n_1161),
.B2(n_1167),
.Y(n_1316)
);

CKINVDCx11_ASAP7_75t_R g1317 ( 
.A(n_1144),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1241),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1129),
.B(n_1253),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1184),
.A2(n_1173),
.B(n_1172),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1176),
.A2(n_1179),
.B(n_1183),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1179),
.A2(n_1174),
.B(n_1132),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1205),
.A2(n_1158),
.B(n_1153),
.C(n_1222),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1217),
.A2(n_1187),
.B1(n_1243),
.B2(n_1247),
.Y(n_1324)
);

NOR2x1_ASAP7_75t_SL g1325 ( 
.A(n_1187),
.B(n_1139),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1165),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1181),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1118),
.B(n_1236),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1132),
.A2(n_1198),
.B(n_1251),
.Y(n_1329)
);

AND2x6_ASAP7_75t_L g1330 ( 
.A(n_1138),
.B(n_1205),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1198),
.A2(n_1251),
.B(n_1193),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1193),
.A2(n_1251),
.B(n_1126),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1118),
.B(n_1236),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1114),
.A2(n_1158),
.B(n_1205),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1158),
.A2(n_1126),
.B(n_1153),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_SL g1336 ( 
.A1(n_1178),
.A2(n_1153),
.B(n_1126),
.C(n_1175),
.Y(n_1336)
);

NAND2xp33_ASAP7_75t_L g1337 ( 
.A(n_1232),
.B(n_1139),
.Y(n_1337)
);

NOR2x1_ASAP7_75t_SL g1338 ( 
.A(n_1186),
.B(n_1200),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1240),
.B(n_1242),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1232),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1242),
.B(n_1144),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1232),
.A2(n_654),
.B(n_899),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1170),
.Y(n_1343)
);

AOI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1197),
.A2(n_1237),
.B(n_1230),
.Y(n_1344)
);

NAND2x1p5_ASAP7_75t_L g1345 ( 
.A(n_1222),
.B(n_1175),
.Y(n_1345)
);

OA21x2_ASAP7_75t_L g1346 ( 
.A1(n_1119),
.A2(n_1116),
.B(n_1188),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1170),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1128),
.A2(n_1230),
.B(n_1197),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1128),
.A2(n_1230),
.B(n_1197),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1232),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1125),
.B(n_919),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1245),
.A2(n_654),
.B(n_899),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1159),
.Y(n_1353)
);

OA21x2_ASAP7_75t_L g1354 ( 
.A1(n_1119),
.A2(n_1116),
.B(n_1188),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1159),
.Y(n_1355)
);

AOI222xp33_ASAP7_75t_L g1356 ( 
.A1(n_1212),
.A2(n_676),
.B1(n_484),
.B2(n_438),
.C1(n_647),
.C2(n_677),
.Y(n_1356)
);

BUFx4_ASAP7_75t_SL g1357 ( 
.A(n_1223),
.Y(n_1357)
);

AOI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1197),
.A2(n_1237),
.B(n_1230),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1128),
.A2(n_1230),
.B(n_1197),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1152),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1170),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1218),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1218),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1128),
.A2(n_1230),
.B(n_1197),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1160),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1115),
.B(n_1238),
.Y(n_1366)
);

CKINVDCx16_ASAP7_75t_R g1367 ( 
.A(n_1223),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1128),
.A2(n_1230),
.B(n_1197),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1218),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1160),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1128),
.A2(n_1230),
.B(n_1197),
.Y(n_1371)
);

AO31x2_ASAP7_75t_L g1372 ( 
.A1(n_1219),
.A2(n_1234),
.A3(n_1047),
.B(n_1148),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1212),
.A2(n_1227),
.B1(n_733),
.B2(n_1219),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1128),
.A2(n_1230),
.B(n_1197),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1128),
.A2(n_1230),
.B(n_1197),
.Y(n_1375)
);

INVx6_ASAP7_75t_L g1376 ( 
.A(n_1117),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1119),
.A2(n_1116),
.B(n_1188),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1150),
.A2(n_1163),
.B(n_1004),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1212),
.A2(n_676),
.B1(n_1227),
.B2(n_484),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1351),
.A2(n_1267),
.B(n_1352),
.C(n_1260),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1307),
.B(n_1301),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1256),
.A2(n_1258),
.B(n_1351),
.Y(n_1382)
);

O2A1O1Ixp5_ASAP7_75t_L g1383 ( 
.A1(n_1373),
.A2(n_1282),
.B(n_1315),
.C(n_1342),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1307),
.B(n_1301),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1262),
.A2(n_1263),
.B(n_1289),
.C(n_1323),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1288),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1295),
.B(n_1266),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1356),
.A2(n_1263),
.B(n_1292),
.C(n_1373),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1303),
.B(n_1362),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1304),
.Y(n_1390)
);

AOI21x1_ASAP7_75t_SL g1391 ( 
.A1(n_1309),
.A2(n_1378),
.B(n_1259),
.Y(n_1391)
);

AOI221x1_ASAP7_75t_SL g1392 ( 
.A1(n_1290),
.A2(n_1295),
.B1(n_1324),
.B2(n_1261),
.C(n_1366),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1262),
.A2(n_1289),
.B1(n_1379),
.B2(n_1291),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1363),
.Y(n_1394)
);

AOI211xp5_ASAP7_75t_L g1395 ( 
.A1(n_1323),
.A2(n_1302),
.B(n_1334),
.C(n_1297),
.Y(n_1395)
);

O2A1O1Ixp5_ASAP7_75t_L g1396 ( 
.A1(n_1344),
.A2(n_1358),
.B(n_1290),
.C(n_1309),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1379),
.A2(n_1291),
.B1(n_1305),
.B2(n_1369),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1378),
.A2(n_1336),
.B(n_1279),
.C(n_1281),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1312),
.B(n_1275),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1305),
.A2(n_1286),
.B1(n_1327),
.B2(n_1277),
.Y(n_1400)
);

OAI31xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1310),
.A2(n_1330),
.A3(n_1329),
.B(n_1340),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1340),
.B(n_1322),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1257),
.B(n_1268),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1328),
.B(n_1333),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1296),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1283),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1353),
.B(n_1355),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1357),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1319),
.B(n_1299),
.Y(n_1409)
);

NOR2xp67_ASAP7_75t_L g1410 ( 
.A(n_1360),
.B(n_1304),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1318),
.Y(n_1411)
);

BUFx8_ASAP7_75t_SL g1412 ( 
.A(n_1370),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1326),
.Y(n_1413)
);

NOR2xp67_ASAP7_75t_L g1414 ( 
.A(n_1327),
.B(n_1270),
.Y(n_1414)
);

NOR2xp67_ASAP7_75t_L g1415 ( 
.A(n_1270),
.B(n_1271),
.Y(n_1415)
);

AOI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1336),
.A2(n_1308),
.B1(n_1313),
.B2(n_1273),
.C(n_1284),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1341),
.A2(n_1337),
.B(n_1278),
.C(n_1265),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1345),
.A2(n_1350),
.B(n_1325),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1367),
.A2(n_1316),
.B1(n_1276),
.B2(n_1272),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1280),
.A2(n_1377),
.B(n_1354),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1348),
.A2(n_1349),
.B(n_1364),
.Y(n_1421)
);

INVx3_ASAP7_75t_SL g1422 ( 
.A(n_1365),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1320),
.Y(n_1423)
);

CKINVDCx6p67_ASAP7_75t_R g1424 ( 
.A(n_1370),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1293),
.B(n_1335),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1293),
.B(n_1335),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1335),
.B(n_1372),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1264),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1331),
.Y(n_1429)
);

AOI21x1_ASAP7_75t_SL g1430 ( 
.A1(n_1306),
.A2(n_1317),
.B(n_1300),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1298),
.Y(n_1431)
);

O2A1O1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1337),
.A2(n_1278),
.B(n_1345),
.C(n_1272),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1339),
.B(n_1273),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1317),
.B(n_1298),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1372),
.B(n_1332),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1377),
.Y(n_1436)
);

O2A1O1Ixp5_ASAP7_75t_L g1437 ( 
.A1(n_1264),
.A2(n_1343),
.B(n_1269),
.C(n_1285),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1296),
.B(n_1372),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1372),
.Y(n_1439)
);

AOI21x1_ASAP7_75t_SL g1440 ( 
.A1(n_1359),
.A2(n_1375),
.B(n_1374),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1276),
.A2(n_1376),
.B1(n_1365),
.B2(n_1255),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1271),
.A2(n_1376),
.B1(n_1377),
.B2(n_1280),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1280),
.A2(n_1346),
.B(n_1354),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1338),
.B(n_1321),
.Y(n_1444)
);

AOI21x1_ASAP7_75t_SL g1445 ( 
.A1(n_1368),
.A2(n_1371),
.B(n_1274),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1285),
.B(n_1361),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1346),
.B(n_1354),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_SL g1448 ( 
.A1(n_1346),
.A2(n_1294),
.B(n_1347),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1311),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1314),
.B(n_1294),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1287),
.A2(n_1347),
.B(n_1361),
.Y(n_1451)
);

BUFx4f_ASAP7_75t_L g1452 ( 
.A(n_1294),
.Y(n_1452)
);

AOI21x1_ASAP7_75t_SL g1453 ( 
.A1(n_1309),
.A2(n_1133),
.B(n_1009),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1256),
.A2(n_1254),
.B(n_1258),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1351),
.A2(n_1263),
.B1(n_1267),
.B2(n_1258),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1312),
.B(n_1259),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1340),
.B(n_1322),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1307),
.B(n_1301),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1351),
.A2(n_1234),
.B(n_1219),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1351),
.A2(n_1267),
.B(n_1352),
.C(n_743),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1351),
.A2(n_1267),
.B(n_1352),
.C(n_743),
.Y(n_1461)
);

O2A1O1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1351),
.A2(n_1267),
.B(n_1352),
.C(n_743),
.Y(n_1462)
);

NOR2xp67_ASAP7_75t_L g1463 ( 
.A(n_1260),
.B(n_1305),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1303),
.B(n_1288),
.Y(n_1464)
);

BUFx12f_ASAP7_75t_L g1465 ( 
.A(n_1365),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1452),
.B(n_1436),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1423),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1420),
.A2(n_1443),
.B(n_1445),
.Y(n_1468)
);

INVx4_ASAP7_75t_L g1469 ( 
.A(n_1444),
.Y(n_1469)
);

OR2x6_ASAP7_75t_L g1470 ( 
.A(n_1459),
.B(n_1418),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1431),
.B(n_1434),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1406),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1427),
.B(n_1435),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1387),
.B(n_1398),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1439),
.B(n_1389),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1411),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1429),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1464),
.B(n_1438),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1402),
.B(n_1457),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1448),
.A2(n_1447),
.B(n_1385),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1455),
.B(n_1382),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1457),
.B(n_1425),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1426),
.B(n_1450),
.Y(n_1483)
);

AO21x1_ASAP7_75t_SL g1484 ( 
.A1(n_1449),
.A2(n_1385),
.B(n_1430),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1413),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1386),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1393),
.A2(n_1454),
.B1(n_1397),
.B2(n_1388),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1442),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1403),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1407),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1451),
.B(n_1456),
.Y(n_1491)
);

AO21x2_ASAP7_75t_L g1492 ( 
.A1(n_1380),
.A2(n_1460),
.B(n_1461),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1381),
.B(n_1458),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1395),
.B(n_1421),
.Y(n_1494)
);

BUFx2_ASAP7_75t_SL g1495 ( 
.A(n_1463),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1421),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1421),
.B(n_1396),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1462),
.A2(n_1383),
.B(n_1396),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1409),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1399),
.B(n_1394),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1428),
.B(n_1383),
.Y(n_1501)
);

AO21x2_ASAP7_75t_L g1502 ( 
.A1(n_1446),
.A2(n_1384),
.B(n_1391),
.Y(n_1502)
);

AO21x2_ASAP7_75t_L g1503 ( 
.A1(n_1391),
.A2(n_1453),
.B(n_1432),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1401),
.B(n_1416),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1437),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1437),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1483),
.B(n_1404),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1467),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1474),
.B(n_1392),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1475),
.B(n_1494),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1469),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1474),
.B(n_1390),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1491),
.B(n_1419),
.Y(n_1513)
);

AO21x2_ASAP7_75t_L g1514 ( 
.A1(n_1498),
.A2(n_1430),
.B(n_1453),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1481),
.B(n_1400),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1498),
.A2(n_1410),
.B(n_1440),
.Y(n_1516)
);

AOI21xp33_ASAP7_75t_L g1517 ( 
.A1(n_1481),
.A2(n_1492),
.B(n_1487),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1494),
.B(n_1405),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1494),
.B(n_1433),
.Y(n_1519)
);

INVx5_ASAP7_75t_L g1520 ( 
.A(n_1470),
.Y(n_1520)
);

INVx4_ASAP7_75t_L g1521 ( 
.A(n_1492),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1482),
.B(n_1408),
.Y(n_1522)
);

OAI211xp5_ASAP7_75t_SL g1523 ( 
.A1(n_1487),
.A2(n_1441),
.B(n_1417),
.C(n_1424),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1502),
.B(n_1489),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1480),
.B(n_1408),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1488),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1488),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1502),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1480),
.B(n_1415),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1480),
.B(n_1422),
.Y(n_1530)
);

INVx1_ASAP7_75t_SL g1531 ( 
.A(n_1530),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1517),
.A2(n_1492),
.B(n_1488),
.Y(n_1532)
);

OAI221xp5_ASAP7_75t_SL g1533 ( 
.A1(n_1509),
.A2(n_1504),
.B1(n_1470),
.B2(n_1501),
.C(n_1478),
.Y(n_1533)
);

OAI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1517),
.A2(n_1504),
.B1(n_1470),
.B2(n_1473),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1517),
.A2(n_1504),
.B1(n_1492),
.B2(n_1484),
.Y(n_1535)
);

NAND3xp33_ASAP7_75t_SL g1536 ( 
.A(n_1515),
.B(n_1493),
.C(n_1478),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1515),
.A2(n_1492),
.B(n_1480),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1511),
.B(n_1469),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1512),
.B(n_1493),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1526),
.A2(n_1495),
.B1(n_1470),
.B2(n_1486),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1521),
.A2(n_1484),
.B1(n_1470),
.B2(n_1480),
.Y(n_1541)
);

OA21x2_ASAP7_75t_L g1542 ( 
.A1(n_1528),
.A2(n_1496),
.B(n_1468),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1521),
.B(n_1495),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1512),
.Y(n_1544)
);

BUFx6f_ASAP7_75t_L g1545 ( 
.A(n_1520),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1508),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1525),
.B(n_1500),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1510),
.B(n_1475),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1530),
.Y(n_1549)
);

OAI211xp5_ASAP7_75t_L g1550 ( 
.A1(n_1521),
.A2(n_1486),
.B(n_1497),
.C(n_1469),
.Y(n_1550)
);

AOI211xp5_ASAP7_75t_SL g1551 ( 
.A1(n_1523),
.A2(n_1414),
.B(n_1497),
.C(n_1466),
.Y(n_1551)
);

AOI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1521),
.A2(n_1506),
.B1(n_1505),
.B2(n_1490),
.C(n_1489),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1510),
.B(n_1475),
.Y(n_1553)
);

OAI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1526),
.A2(n_1505),
.B1(n_1490),
.B2(n_1499),
.C(n_1485),
.Y(n_1554)
);

AOI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1528),
.A2(n_1497),
.B1(n_1485),
.B2(n_1499),
.C(n_1472),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1526),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1526),
.A2(n_1471),
.B1(n_1479),
.B2(n_1503),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1510),
.B(n_1486),
.Y(n_1558)
);

OAI321xp33_ASAP7_75t_L g1559 ( 
.A1(n_1523),
.A2(n_1530),
.A3(n_1525),
.B1(n_1529),
.B2(n_1510),
.C(n_1518),
.Y(n_1559)
);

OAI211xp5_ASAP7_75t_L g1560 ( 
.A1(n_1530),
.A2(n_1469),
.B(n_1476),
.C(n_1477),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1559),
.B(n_1527),
.Y(n_1561)
);

BUFx12f_ASAP7_75t_L g1562 ( 
.A(n_1556),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1543),
.B(n_1529),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1546),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1542),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1546),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1548),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1548),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1553),
.Y(n_1569)
);

INVx4_ASAP7_75t_L g1570 ( 
.A(n_1556),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1553),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1542),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1542),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1544),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1543),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1554),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1537),
.B(n_1495),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1532),
.A2(n_1524),
.B(n_1496),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1545),
.Y(n_1579)
);

AND2x6_ASAP7_75t_SL g1580 ( 
.A(n_1539),
.B(n_1412),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1558),
.Y(n_1581)
);

INVx4_ASAP7_75t_SL g1582 ( 
.A(n_1545),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1552),
.B(n_1527),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1559),
.A2(n_1527),
.B(n_1514),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1558),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1543),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1536),
.B(n_1527),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1555),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_SL g1589 ( 
.A1(n_1540),
.A2(n_1514),
.B(n_1516),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1547),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1562),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1567),
.B(n_1533),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1588),
.B(n_1513),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1574),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1567),
.B(n_1519),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1568),
.B(n_1569),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1582),
.B(n_1518),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1565),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1588),
.B(n_1513),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1574),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1576),
.A2(n_1535),
.B1(n_1534),
.B2(n_1541),
.Y(n_1601)
);

BUFx12f_ASAP7_75t_L g1602 ( 
.A(n_1580),
.Y(n_1602)
);

OR2x6_ASAP7_75t_L g1603 ( 
.A(n_1589),
.B(n_1545),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1582),
.B(n_1538),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1564),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1582),
.B(n_1538),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1569),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1576),
.B(n_1513),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1564),
.Y(n_1609)
);

INVx5_ASAP7_75t_L g1610 ( 
.A(n_1579),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1566),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1571),
.B(n_1531),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1566),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1565),
.Y(n_1614)
);

NOR2x1_ASAP7_75t_L g1615 ( 
.A(n_1570),
.B(n_1560),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1582),
.B(n_1538),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1587),
.Y(n_1617)
);

OAI21xp33_ASAP7_75t_L g1618 ( 
.A1(n_1583),
.A2(n_1584),
.B(n_1561),
.Y(n_1618)
);

NAND2x1p5_ASAP7_75t_SL g1619 ( 
.A(n_1589),
.B(n_1522),
.Y(n_1619)
);

NOR2x1_ASAP7_75t_L g1620 ( 
.A(n_1570),
.B(n_1540),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1581),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1583),
.B(n_1531),
.Y(n_1622)
);

NAND4xp25_ASAP7_75t_L g1623 ( 
.A(n_1584),
.B(n_1551),
.C(n_1557),
.D(n_1550),
.Y(n_1623)
);

AND2x4_ASAP7_75t_SL g1624 ( 
.A(n_1570),
.B(n_1522),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1593),
.B(n_1599),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1594),
.Y(n_1626)
);

NAND2x2_ASAP7_75t_L g1627 ( 
.A(n_1591),
.B(n_1575),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1619),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1597),
.B(n_1582),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1593),
.B(n_1587),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1619),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1600),
.Y(n_1632)
);

NOR2x1_ASAP7_75t_L g1633 ( 
.A(n_1620),
.B(n_1570),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1597),
.B(n_1590),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1624),
.B(n_1590),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1599),
.B(n_1585),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1605),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1608),
.B(n_1549),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1603),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1609),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1611),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1624),
.B(n_1563),
.Y(n_1642)
);

XNOR2xp5_ASAP7_75t_L g1643 ( 
.A(n_1601),
.B(n_1580),
.Y(n_1643)
);

NAND2x1p5_ASAP7_75t_L g1644 ( 
.A(n_1610),
.B(n_1520),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1617),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1613),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1604),
.B(n_1563),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1621),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1603),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1596),
.Y(n_1650)
);

A2O1A1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1618),
.A2(n_1551),
.B(n_1575),
.C(n_1586),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1608),
.B(n_1578),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1604),
.B(n_1575),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1602),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1607),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1595),
.B(n_1578),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1617),
.B(n_1507),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1598),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1598),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1645),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1652),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1625),
.B(n_1592),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1637),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1654),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1640),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1652),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1654),
.B(n_1412),
.Y(n_1667)
);

NOR2x1_ASAP7_75t_L g1668 ( 
.A(n_1643),
.B(n_1623),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1641),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1633),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1628),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1646),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_1643),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1628),
.Y(n_1674)
);

OAI21x1_ASAP7_75t_L g1675 ( 
.A1(n_1631),
.A2(n_1615),
.B(n_1614),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1647),
.B(n_1606),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1647),
.B(n_1629),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1636),
.B(n_1612),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1650),
.B(n_1601),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1653),
.Y(n_1680)
);

OAI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1631),
.A2(n_1603),
.B1(n_1577),
.B2(n_1622),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1648),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1626),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1629),
.B(n_1606),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1664),
.B(n_1422),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1664),
.B(n_1653),
.Y(n_1686)
);

OAI322xp33_ASAP7_75t_L g1687 ( 
.A1(n_1679),
.A2(n_1662),
.A3(n_1674),
.B1(n_1671),
.B2(n_1683),
.C1(n_1660),
.C2(n_1670),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1671),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1668),
.B(n_1655),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1668),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1671),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1662),
.B(n_1630),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1674),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1674),
.Y(n_1694)
);

XOR2x2_ASAP7_75t_L g1695 ( 
.A(n_1673),
.B(n_1644),
.Y(n_1695)
);

NAND2x1p5_ASAP7_75t_L g1696 ( 
.A(n_1664),
.B(n_1680),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1661),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1680),
.B(n_1673),
.Y(n_1698)
);

AOI21xp33_ASAP7_75t_SL g1699 ( 
.A1(n_1675),
.A2(n_1651),
.B(n_1629),
.Y(n_1699)
);

NOR2x1_ASAP7_75t_L g1700 ( 
.A(n_1680),
.B(n_1667),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1660),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1676),
.B(n_1653),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1673),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1690),
.A2(n_1651),
.B1(n_1627),
.B2(n_1679),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1702),
.B(n_1677),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1690),
.B(n_1677),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1703),
.A2(n_1666),
.B1(n_1661),
.B2(n_1577),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1697),
.A2(n_1666),
.B1(n_1661),
.B2(n_1577),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1700),
.B(n_1684),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1697),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1698),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_L g1712 ( 
.A(n_1687),
.B(n_1681),
.C(n_1670),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1688),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1686),
.B(n_1684),
.Y(n_1714)
);

OAI221xp5_ASAP7_75t_L g1715 ( 
.A1(n_1712),
.A2(n_1699),
.B1(n_1689),
.B2(n_1666),
.C(n_1693),
.Y(n_1715)
);

OAI21xp33_ASAP7_75t_SL g1716 ( 
.A1(n_1710),
.A2(n_1675),
.B(n_1686),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1704),
.A2(n_1695),
.B1(n_1694),
.B2(n_1691),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1706),
.A2(n_1675),
.B(n_1685),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1709),
.B(n_1676),
.Y(n_1719)
);

AND5x1_ASAP7_75t_L g1720 ( 
.A(n_1714),
.B(n_1685),
.C(n_1696),
.D(n_1692),
.E(n_1681),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1707),
.A2(n_1627),
.B1(n_1659),
.B2(n_1658),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1711),
.B(n_1696),
.Y(n_1722)
);

OAI21xp33_ASAP7_75t_SL g1723 ( 
.A1(n_1705),
.A2(n_1701),
.B(n_1683),
.Y(n_1723)
);

NOR3xp33_ASAP7_75t_L g1724 ( 
.A(n_1711),
.B(n_1665),
.C(n_1663),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1713),
.B(n_1663),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1719),
.B(n_1665),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1715),
.A2(n_1708),
.B1(n_1682),
.B2(n_1669),
.C(n_1672),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1716),
.A2(n_1639),
.B1(n_1649),
.B2(n_1614),
.Y(n_1728)
);

AOI322xp5_ASAP7_75t_L g1729 ( 
.A1(n_1717),
.A2(n_1622),
.A3(n_1682),
.B1(n_1669),
.B2(n_1672),
.C1(n_1573),
.C2(n_1572),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1722),
.Y(n_1730)
);

XNOR2xp5_ASAP7_75t_L g1731 ( 
.A(n_1730),
.B(n_1721),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1726),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1728),
.B(n_1678),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1729),
.B(n_1678),
.Y(n_1734)
);

AOI21xp33_ASAP7_75t_SL g1735 ( 
.A1(n_1727),
.A2(n_1723),
.B(n_1724),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1730),
.B(n_1718),
.Y(n_1736)
);

XNOR2x1_ASAP7_75t_L g1737 ( 
.A(n_1731),
.B(n_1720),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1736),
.A2(n_1725),
.B(n_1632),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1732),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1733),
.Y(n_1740)
);

INVx2_ASAP7_75t_SL g1741 ( 
.A(n_1734),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1740),
.B(n_1735),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1739),
.B(n_1635),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1741),
.B(n_1635),
.Y(n_1744)
);

NAND3xp33_ASAP7_75t_L g1745 ( 
.A(n_1742),
.B(n_1740),
.C(n_1737),
.Y(n_1745)
);

AOI322xp5_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1744),
.A3(n_1743),
.B1(n_1738),
.B2(n_1639),
.C1(n_1649),
.C2(n_1573),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1746),
.A2(n_1638),
.B1(n_1656),
.B2(n_1657),
.Y(n_1747)
);

NAND3xp33_ASAP7_75t_SL g1748 ( 
.A(n_1746),
.B(n_1656),
.C(n_1644),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1747),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1748),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1749),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1750),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1751),
.Y(n_1753)
);

OA22x2_ASAP7_75t_L g1754 ( 
.A1(n_1753),
.A2(n_1752),
.B1(n_1642),
.B2(n_1634),
.Y(n_1754)
);

AOI222xp33_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1465),
.B1(n_1634),
.B2(n_1610),
.C1(n_1642),
.C2(n_1562),
.Y(n_1755)
);

XNOR2xp5_ASAP7_75t_L g1756 ( 
.A(n_1755),
.B(n_1465),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1756),
.A2(n_1638),
.B1(n_1610),
.B2(n_1644),
.Y(n_1757)
);

AOI211xp5_ASAP7_75t_L g1758 ( 
.A1(n_1757),
.A2(n_1586),
.B(n_1616),
.C(n_1573),
.Y(n_1758)
);


endmodule