module fake_jpeg_11844_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_39),
.Y(n_109)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_47),
.Y(n_114)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx6p67_ASAP7_75t_R g100 ( 
.A(n_55),
.Y(n_100)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx2_ASAP7_75t_SL g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_20),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_62),
.Y(n_78)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_66),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_31),
.A2(n_15),
.B1(n_14),
.B2(n_2),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_65),
.A2(n_27),
.B1(n_22),
.B2(n_18),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_18),
.B(n_14),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_71),
.Y(n_85)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_70),
.Y(n_101)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_38),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_33),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_23),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_38),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_36),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_93),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_36),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_35),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_32),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_40),
.A2(n_25),
.B1(n_34),
.B2(n_28),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_97),
.A2(n_104),
.B1(n_38),
.B2(n_32),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_33),
.C(n_35),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_102),
.A2(n_80),
.B(n_101),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_41),
.A2(n_25),
.B1(n_34),
.B2(n_28),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_27),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_37),
.B1(n_22),
.B2(n_16),
.Y(n_116)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_116),
.A2(n_118),
.B1(n_134),
.B2(n_114),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_113),
.A2(n_73),
.B1(n_67),
.B2(n_39),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_55),
.B(n_37),
.C(n_16),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_120),
.B(n_80),
.Y(n_166)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_123),
.Y(n_159)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_126),
.A2(n_144),
.B1(n_151),
.B2(n_154),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_128),
.B(n_98),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_129),
.B(n_87),
.Y(n_164)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_53),
.B1(n_69),
.B2(n_54),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_114),
.B1(n_100),
.B2(n_84),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_34),
.B1(n_25),
.B2(n_28),
.Y(n_132)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_80),
.B(n_17),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_77),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_152),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_85),
.A2(n_44),
.B1(n_52),
.B2(n_51),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_87),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_149),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_96),
.A2(n_16),
.B1(n_64),
.B2(n_33),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_0),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_0),
.Y(n_156)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_153),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_81),
.A2(n_47),
.B1(n_66),
.B2(n_17),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_81),
.A2(n_17),
.B1(n_21),
.B2(n_2),
.Y(n_154)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_100),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_156),
.B(n_166),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_158),
.A2(n_112),
.B1(n_107),
.B2(n_115),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_78),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_167),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_164),
.B(n_193),
.C(n_0),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_108),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_108),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_180),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_95),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_176),
.B(n_187),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_137),
.B1(n_136),
.B2(n_79),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_95),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_123),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_192),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_182),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_92),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_149),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_121),
.B(n_145),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_0),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_146),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_129),
.B(n_103),
.C(n_86),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_132),
.B1(n_135),
.B2(n_139),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_195),
.A2(n_203),
.B1(n_205),
.B2(n_216),
.Y(n_240)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

AOI32xp33_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_136),
.A3(n_120),
.B1(n_155),
.B2(n_147),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_197),
.A2(n_208),
.B(n_159),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_198),
.Y(n_263)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_136),
.B(n_148),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_201),
.A2(n_159),
.B(n_172),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_188),
.A2(n_109),
.B1(n_84),
.B2(n_130),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_170),
.B(n_190),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_204),
.B(n_212),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_167),
.A2(n_112),
.B1(n_107),
.B2(n_122),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_161),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_231),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_164),
.A2(n_152),
.B(n_150),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_213),
.B(n_160),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_164),
.A2(n_143),
.B1(n_103),
.B2(n_86),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_209),
.A2(n_221),
.B1(n_226),
.B2(n_183),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_223),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_157),
.B(n_141),
.Y(n_212)
);

AND2x2_ASAP7_75t_SL g213 ( 
.A(n_193),
.B(n_140),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_178),
.A2(n_124),
.B1(n_21),
.B2(n_14),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_169),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_229),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_184),
.B1(n_169),
.B2(n_156),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_21),
.B1(n_3),
.B2(n_4),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_179),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_5),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_160),
.C(n_186),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_160),
.B(n_5),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_162),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_162),
.B(n_8),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_186),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_8),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_194),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_232),
.B(n_243),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_234),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_238),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_158),
.B1(n_174),
.B2(n_173),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_242),
.A2(n_247),
.B1(n_264),
.B2(n_245),
.Y(n_286)
);

NOR2x1_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_172),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_246),
.A2(n_249),
.B(n_228),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_215),
.A2(n_174),
.B1(n_171),
.B2(n_173),
.Y(n_247)
);

AOI22x1_ASAP7_75t_SL g249 ( 
.A1(n_197),
.A2(n_191),
.B1(n_174),
.B2(n_189),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_258),
.B(n_266),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_252),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_191),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_175),
.C(n_189),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_257),
.Y(n_278)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_213),
.B(n_175),
.C(n_177),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_201),
.A2(n_183),
.B(n_168),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_196),
.Y(n_259)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_260),
.A2(n_203),
.B1(n_216),
.B2(n_220),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_213),
.B(n_177),
.C(n_10),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_9),
.Y(n_284)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_205),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_222),
.A2(n_204),
.B1(n_202),
.B2(n_195),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_206),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_265),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_207),
.A2(n_9),
.B(n_10),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_234),
.A2(n_208),
.B(n_222),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_267),
.A2(n_275),
.B(n_246),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_214),
.B1(n_217),
.B2(n_200),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_271),
.A2(n_277),
.B1(n_280),
.B2(n_285),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_199),
.B(n_223),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_240),
.A2(n_202),
.B1(n_221),
.B2(n_211),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_240),
.A2(n_263),
.B1(n_262),
.B2(n_251),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_239),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_284),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_283),
.A2(n_292),
.B1(n_293),
.B2(n_266),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_263),
.A2(n_226),
.B1(n_224),
.B2(n_210),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_254),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_287),
.A2(n_258),
.B(n_243),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_244),
.B(n_227),
.Y(n_288)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_288),
.Y(n_298)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_248),
.Y(n_289)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_229),
.B1(n_218),
.B2(n_12),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_294),
.B1(n_259),
.B2(n_235),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_242),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_293)
);

OAI22x1_ASAP7_75t_SL g294 ( 
.A1(n_236),
.A2(n_13),
.B1(n_245),
.B2(n_241),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_237),
.B(n_247),
.Y(n_295)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_295),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_281),
.B(n_241),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_297),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_269),
.B(n_236),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_299),
.B(n_310),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_233),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_304),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_291),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_303),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_268),
.B(n_233),
.Y(n_304)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_305),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_287),
.Y(n_328)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_270),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_309),
.A2(n_282),
.B(n_275),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_255),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_286),
.A2(n_257),
.B1(n_261),
.B2(n_238),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_311),
.A2(n_312),
.B1(n_278),
.B2(n_285),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_286),
.A2(n_283),
.B1(n_295),
.B2(n_273),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_273),
.A2(n_248),
.B(n_256),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_313),
.A2(n_316),
.B(n_282),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_314),
.A2(n_318),
.B1(n_283),
.B2(n_279),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_276),
.A2(n_235),
.B(n_255),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_291),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_317),
.A2(n_319),
.B1(n_320),
.B2(n_272),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_280),
.A2(n_271),
.B1(n_277),
.B2(n_267),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_289),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_278),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_330),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_313),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_299),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_327),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_336),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_331),
.A2(n_332),
.B(n_306),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_288),
.C(n_274),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_298),
.C(n_315),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_274),
.Y(n_336)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_337),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_312),
.A2(n_279),
.B1(n_290),
.B2(n_294),
.Y(n_338)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_338),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_303),
.Y(n_339)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_339),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_308),
.B(n_284),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_341),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_292),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_343),
.A2(n_332),
.B1(n_320),
.B2(n_301),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_334),
.A2(n_309),
.B(n_318),
.Y(n_344)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_344),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_347),
.C(n_355),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_316),
.C(n_315),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_335),
.B(n_307),
.Y(n_352)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_352),
.Y(n_361)
);

OAI221xp5_ASAP7_75t_L g370 ( 
.A1(n_353),
.A2(n_330),
.B1(n_340),
.B2(n_301),
.C(n_319),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_300),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_331),
.A2(n_300),
.B(n_297),
.Y(n_356)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_356),
.Y(n_364)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_324),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_357),
.A2(n_325),
.B1(n_338),
.B2(n_317),
.Y(n_363)
);

FAx1_ASAP7_75t_SL g358 ( 
.A(n_347),
.B(n_333),
.CI(n_322),
.CON(n_358),
.SN(n_358)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_367),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_348),
.B(n_355),
.C(n_345),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_363),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_350),
.A2(n_329),
.B1(n_337),
.B2(n_305),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_365),
.B(n_366),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_350),
.A2(n_329),
.B1(n_341),
.B2(n_328),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_346),
.B(n_296),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_336),
.C(n_323),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_351),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_344),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_370),
.A2(n_354),
.B1(n_352),
.B2(n_342),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_362),
.A2(n_353),
.B(n_343),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_371),
.B(n_372),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_349),
.C(n_342),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_359),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_375),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_359),
.B(n_366),
.C(n_349),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_356),
.C(n_362),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_381),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_380),
.A2(n_364),
.B(n_361),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_351),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_390),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_376),
.B(n_358),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_385),
.B(n_388),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_386),
.B(n_365),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_377),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_374),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_389),
.Y(n_395)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_380),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_389),
.B(n_378),
.C(n_372),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_392),
.A2(n_387),
.B(n_382),
.Y(n_397)
);

O2A1O1Ixp33_ASAP7_75t_SL g393 ( 
.A1(n_386),
.A2(n_375),
.B(n_364),
.C(n_358),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_393),
.B(n_314),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_394),
.B(n_357),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_397),
.B(n_399),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_396),
.B(n_384),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_398),
.A2(n_400),
.B(n_391),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_402),
.A2(n_396),
.B(n_395),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_401),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_404),
.A2(n_272),
.B(n_292),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_405),
.A2(n_294),
.B(n_293),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_293),
.Y(n_407)
);


endmodule