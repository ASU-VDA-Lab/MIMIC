module real_aes_2391_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_379;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_171;
wire n_87;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_0), .Y(n_126) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_1), .A2(n_50), .B1(n_92), .B2(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_2), .B(n_213), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_3), .B(n_228), .Y(n_246) );
INVx1_ASAP7_75t_L g200 ( .A(n_4), .Y(n_200) );
OAI22xp5_ASAP7_75t_SL g182 ( .A1(n_5), .A2(n_70), .B1(n_183), .B2(n_184), .Y(n_182) );
INVx1_ASAP7_75t_L g184 ( .A(n_5), .Y(n_184) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_6), .A2(n_16), .B1(n_92), .B2(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g248 ( .A(n_7), .B(n_237), .Y(n_248) );
AND2x2_ASAP7_75t_L g257 ( .A(n_8), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g234 ( .A(n_9), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_10), .B(n_228), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_11), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_12), .B(n_213), .Y(n_282) );
AOI22xp33_ASAP7_75t_SL g163 ( .A1(n_13), .A2(n_15), .B1(n_164), .B2(n_167), .Y(n_163) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_14), .A2(n_69), .B1(n_213), .B2(n_320), .Y(n_319) );
OAI221xp5_ASAP7_75t_L g192 ( .A1(n_16), .A2(n_50), .B1(n_55), .B2(n_193), .C(n_195), .Y(n_192) );
OR2x2_ASAP7_75t_L g235 ( .A(n_17), .B(n_68), .Y(n_235) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_17), .A2(n_68), .B(n_234), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_18), .A2(n_41), .B1(n_154), .B2(n_158), .Y(n_153) );
INVx3_ASAP7_75t_L g92 ( .A(n_19), .Y(n_92) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_20), .A2(n_258), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_21), .B(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_22), .A2(n_221), .B(n_244), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_23), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_24), .B(n_228), .Y(n_277) );
INVx1_ASAP7_75t_SL g93 ( .A(n_25), .Y(n_93) );
INVx1_ASAP7_75t_L g202 ( .A(n_26), .Y(n_202) );
AND2x2_ASAP7_75t_L g219 ( .A(n_26), .B(n_200), .Y(n_219) );
AND2x2_ASAP7_75t_L g222 ( .A(n_26), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_27), .B(n_213), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_28), .B(n_228), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_29), .B(n_213), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_30), .A2(n_221), .B(n_253), .Y(n_252) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_31), .A2(n_55), .B1(n_92), .B2(n_96), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_32), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_33), .B(n_213), .Y(n_264) );
INVx1_ASAP7_75t_L g216 ( .A(n_34), .Y(n_216) );
INVx1_ASAP7_75t_L g225 ( .A(n_34), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_35), .B(n_228), .Y(n_255) );
AND2x2_ASAP7_75t_L g292 ( .A(n_36), .B(n_232), .Y(n_292) );
INVx1_ASAP7_75t_L g94 ( .A(n_37), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_38), .B(n_230), .Y(n_254) );
INVx1_ASAP7_75t_L g542 ( .A(n_38), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_39), .B(n_230), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_40), .B(n_213), .Y(n_256) );
INVx1_ASAP7_75t_L g557 ( .A(n_40), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_42), .B(n_213), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_43), .A2(n_221), .B(n_275), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_44), .A2(n_63), .B1(n_187), .B2(n_188), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_44), .Y(n_188) );
AND2x2_ASAP7_75t_L g287 ( .A(n_45), .B(n_233), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_46), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_47), .B(n_230), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_48), .B(n_230), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_49), .A2(n_72), .B1(n_221), .B2(n_325), .Y(n_324) );
INVxp33_ASAP7_75t_L g197 ( .A(n_50), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_51), .B(n_228), .Y(n_285) );
INVx1_ASAP7_75t_L g218 ( .A(n_52), .Y(n_218) );
INVx1_ASAP7_75t_L g223 ( .A(n_52), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_53), .B(n_230), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_54), .A2(n_66), .B1(n_171), .B2(n_174), .Y(n_170) );
INVxp67_ASAP7_75t_L g196 ( .A(n_55), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_56), .A2(n_221), .B(n_296), .Y(n_295) );
AOI22xp33_ASAP7_75t_SL g146 ( .A1(n_57), .A2(n_67), .B1(n_147), .B2(n_150), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_58), .A2(n_221), .B(n_226), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_59), .A2(n_221), .B(n_266), .Y(n_265) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_60), .A2(n_81), .B1(n_179), .B2(n_550), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_60), .Y(n_550) );
AND2x2_ASAP7_75t_L g279 ( .A(n_61), .B(n_233), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_62), .B(n_232), .Y(n_317) );
INVx1_ASAP7_75t_L g187 ( .A(n_63), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_64), .Y(n_104) );
AND2x2_ASAP7_75t_L g236 ( .A(n_65), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g183 ( .A(n_70), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_71), .A2(n_221), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_73), .B(n_228), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_74), .Y(n_118) );
BUFx2_ASAP7_75t_L g80 ( .A(n_75), .Y(n_80) );
BUFx2_ASAP7_75t_SL g194 ( .A(n_76), .Y(n_194) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_189), .B1(n_203), .B2(n_535), .C(n_539), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_180), .Y(n_78) );
AOI22xp33_ASAP7_75t_R g79 ( .A1(n_80), .A2(n_81), .B1(n_178), .B2(n_179), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g178 ( .A(n_80), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_80), .B(n_230), .Y(n_286) );
INVx1_ASAP7_75t_L g179 ( .A(n_81), .Y(n_179) );
AOI22xp33_ASAP7_75t_R g540 ( .A1(n_81), .A2(n_179), .B1(n_541), .B2(n_542), .Y(n_540) );
INVxp33_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_144), .Y(n_82) );
NOR3xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_117), .C(n_132), .Y(n_83) );
OAI221xp5_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_104), .B1(n_105), .B2(n_106), .C(n_112), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx3_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
INVx6_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_97), .Y(n_88) );
AND2x4_ASAP7_75t_L g129 ( .A(n_89), .B(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g142 ( .A(n_89), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_95), .Y(n_89) );
AND2x2_ASAP7_75t_L g110 ( .A(n_90), .B(n_111), .Y(n_110) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_90), .Y(n_116) );
INVx2_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
OAI22x1_ASAP7_75t_L g90 ( .A1(n_91), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
INVx2_ASAP7_75t_L g100 ( .A(n_92), .Y(n_100) );
INVx1_ASAP7_75t_L g103 ( .A(n_92), .Y(n_103) );
INVx2_ASAP7_75t_L g111 ( .A(n_95), .Y(n_111) );
AND2x2_ASAP7_75t_L g138 ( .A(n_95), .B(n_139), .Y(n_138) );
BUFx2_ASAP7_75t_L g161 ( .A(n_95), .Y(n_161) );
AND2x4_ASAP7_75t_L g149 ( .A(n_97), .B(n_110), .Y(n_149) );
AND2x4_ASAP7_75t_L g166 ( .A(n_97), .B(n_152), .Y(n_166) );
AND2x2_ASAP7_75t_L g173 ( .A(n_97), .B(n_138), .Y(n_173) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_101), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x4_ASAP7_75t_L g109 ( .A(n_99), .B(n_101), .Y(n_109) );
AND2x2_ASAP7_75t_L g115 ( .A(n_99), .B(n_102), .Y(n_115) );
INVx1_ASAP7_75t_L g125 ( .A(n_99), .Y(n_125) );
INVxp67_ASAP7_75t_L g143 ( .A(n_101), .Y(n_143) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g124 ( .A(n_102), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x4_ASAP7_75t_L g137 ( .A(n_109), .B(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g177 ( .A(n_109), .B(n_152), .Y(n_177) );
AND2x2_ASAP7_75t_L g123 ( .A(n_110), .B(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g152 ( .A(n_111), .B(n_139), .Y(n_152) );
BUFx12f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x4_ASAP7_75t_L g151 ( .A(n_115), .B(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g160 ( .A(n_115), .B(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_119), .B1(n_126), .B2(n_127), .Y(n_117) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g157 ( .A(n_124), .B(n_138), .Y(n_157) );
AND2x4_ASAP7_75t_L g169 ( .A(n_124), .B(n_152), .Y(n_169) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_125), .Y(n_131) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B1(n_140), .B2(n_141), .Y(n_132) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx4f_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx6_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_145), .B(n_162), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_153), .Y(n_145) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx6_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx2_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx5_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_170), .Y(n_162) );
INVx2_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
INVx8_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
INVx8_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_SL g171 ( .A(n_172), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B1(n_185), .B2(n_186), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
AND3x1_ASAP7_75t_SL g191 ( .A(n_192), .B(n_198), .C(n_201), .Y(n_191) );
INVxp67_ASAP7_75t_L g548 ( .A(n_192), .Y(n_548) );
CKINVDCx8_ASAP7_75t_R g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
CKINVDCx16_ASAP7_75t_R g546 ( .A(n_198), .Y(n_546) );
AO21x1_ASAP7_75t_SL g554 ( .A1(n_198), .A2(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g321 ( .A(n_199), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_SL g553 ( .A(n_199), .B(n_201), .Y(n_553) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g224 ( .A(n_200), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_201), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2x1p5_ASAP7_75t_L g326 ( .A(n_202), .B(n_327), .Y(n_326) );
INVx5_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_439), .Y(n_204) );
NOR3xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_364), .C(n_400), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_338), .Y(n_206) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_259), .B(n_288), .C(n_313), .Y(n_207) );
AND2x2_ASAP7_75t_L g429 ( .A(n_208), .B(n_290), .Y(n_429) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_239), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_209), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g462 ( .A(n_209), .B(n_344), .Y(n_462) );
AND2x2_ASAP7_75t_L g478 ( .A(n_209), .B(n_305), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_209), .B(n_488), .Y(n_487) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_209), .B(n_512), .Y(n_511) );
INVx4_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x4_ASAP7_75t_SL g300 ( .A(n_210), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g333 ( .A(n_210), .Y(n_333) );
AND2x2_ASAP7_75t_L g380 ( .A(n_210), .B(n_315), .Y(n_380) );
AND2x2_ASAP7_75t_L g399 ( .A(n_210), .B(n_239), .Y(n_399) );
BUFx2_ASAP7_75t_L g404 ( .A(n_210), .Y(n_404) );
AND2x2_ASAP7_75t_L g448 ( .A(n_210), .B(n_249), .Y(n_448) );
AND2x4_ASAP7_75t_L g520 ( .A(n_210), .B(n_521), .Y(n_520) );
NOR2x1_ASAP7_75t_L g532 ( .A(n_210), .B(n_304), .Y(n_532) );
OR2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_236), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_220), .B(n_232), .Y(n_211) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_213), .Y(n_538) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_219), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_215), .B(n_217), .Y(n_214) );
AND2x6_ASAP7_75t_L g230 ( .A(n_215), .B(n_223), .Y(n_230) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x4_ASAP7_75t_L g228 ( .A(n_217), .B(n_225), .Y(n_228) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx5_ASAP7_75t_L g231 ( .A(n_219), .Y(n_231) );
AND2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_224), .Y(n_221) );
BUFx3_ASAP7_75t_L g323 ( .A(n_222), .Y(n_323) );
INVx2_ASAP7_75t_L g328 ( .A(n_223), .Y(n_328) );
AND2x4_ASAP7_75t_L g325 ( .A(n_224), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g322 ( .A(n_225), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_229), .B(n_231), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_231), .A2(n_245), .B(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_231), .A2(n_254), .B(n_255), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_231), .A2(n_267), .B(n_268), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_231), .A2(n_276), .B(n_277), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_231), .A2(n_285), .B(n_286), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_231), .A2(n_297), .B(n_298), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_232), .Y(n_241) );
AO21x2_ASAP7_75t_L g318 ( .A1(n_232), .A2(n_319), .B(n_324), .Y(n_318) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_SL g233 ( .A(n_234), .B(n_235), .Y(n_233) );
AND2x4_ASAP7_75t_L g269 ( .A(n_234), .B(n_235), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_237), .A2(n_282), .B(n_283), .Y(n_281) );
BUFx4f_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx3_ASAP7_75t_L g250 ( .A(n_238), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_239), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g451 ( .A(n_239), .Y(n_451) );
BUFx2_ASAP7_75t_L g500 ( .A(n_239), .Y(n_500) );
INVx1_ASAP7_75t_L g522 ( .A(n_239), .Y(n_522) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_249), .Y(n_239) );
INVx3_ASAP7_75t_L g301 ( .A(n_240), .Y(n_301) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_240), .Y(n_488) );
AOI21x1_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_248), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_247), .Y(n_242) );
INVx2_ASAP7_75t_L g304 ( .A(n_249), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_249), .B(n_301), .Y(n_305) );
INVx2_ASAP7_75t_L g388 ( .A(n_249), .Y(n_388) );
OR2x2_ASAP7_75t_L g395 ( .A(n_249), .B(n_344), .Y(n_395) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_257), .Y(n_249) );
INVx4_ASAP7_75t_L g258 ( .A(n_250), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_256), .Y(n_251) );
INVx3_ASAP7_75t_L g272 ( .A(n_258), .Y(n_272) );
AND2x2_ASAP7_75t_L g350 ( .A(n_259), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g384 ( .A(n_259), .B(n_347), .Y(n_384) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_270), .Y(n_259) );
AND2x2_ASAP7_75t_L g420 ( .A(n_260), .B(n_311), .Y(n_420) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g377 ( .A(n_261), .B(n_271), .Y(n_377) );
AND2x2_ASAP7_75t_L g496 ( .A(n_261), .B(n_280), .Y(n_496) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g310 ( .A(n_262), .Y(n_310) );
INVx1_ASAP7_75t_L g336 ( .A(n_262), .Y(n_336) );
AND2x2_ASAP7_75t_L g392 ( .A(n_262), .B(n_271), .Y(n_392) );
AND2x2_ASAP7_75t_L g397 ( .A(n_262), .B(n_291), .Y(n_397) );
OR2x2_ASAP7_75t_L g460 ( .A(n_262), .B(n_280), .Y(n_460) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_262), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B(n_269), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_269), .A2(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g290 ( .A(n_270), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g337 ( .A(n_270), .Y(n_337) );
NOR2x1_ASAP7_75t_SL g270 ( .A(n_271), .B(n_280), .Y(n_270) );
AO21x1_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_273), .B(n_279), .Y(n_271) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_272), .A2(n_273), .B(n_279), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_278), .Y(n_273) );
AND2x2_ASAP7_75t_L g307 ( .A(n_280), .B(n_308), .Y(n_307) );
INVx2_ASAP7_75t_SL g363 ( .A(n_280), .Y(n_363) );
NAND2x1_ASAP7_75t_L g373 ( .A(n_280), .B(n_291), .Y(n_373) );
OR2x2_ASAP7_75t_L g378 ( .A(n_280), .B(n_308), .Y(n_378) );
BUFx2_ASAP7_75t_L g434 ( .A(n_280), .Y(n_434) );
AND2x2_ASAP7_75t_L g470 ( .A(n_280), .B(n_349), .Y(n_470) );
AND2x2_ASAP7_75t_L g481 ( .A(n_280), .B(n_311), .Y(n_481) );
OR2x6_ASAP7_75t_L g280 ( .A(n_281), .B(n_287), .Y(n_280) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_299), .B1(n_305), .B2(n_306), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_290), .A2(n_478), .B1(n_528), .B2(n_533), .Y(n_527) );
INVx4_ASAP7_75t_L g308 ( .A(n_291), .Y(n_308) );
INVx2_ASAP7_75t_L g347 ( .A(n_291), .Y(n_347) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_291), .Y(n_418) );
OR2x2_ASAP7_75t_L g433 ( .A(n_291), .B(n_311), .Y(n_433) );
OR2x2_ASAP7_75t_SL g459 ( .A(n_291), .B(n_460), .Y(n_459) );
OR2x6_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_SL g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx2_ASAP7_75t_SL g340 ( .A(n_300), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_300), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g408 ( .A(n_300), .B(n_356), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_300), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g330 ( .A(n_301), .Y(n_330) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_301), .Y(n_355) );
AND2x2_ASAP7_75t_L g411 ( .A(n_301), .B(n_388), .Y(n_411) );
INVx1_ASAP7_75t_L g521 ( .A(n_301), .Y(n_521) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_303), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_303), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g329 ( .A(n_304), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_305), .B(n_462), .Y(n_461) );
AOI321xp33_ASAP7_75t_L g483 ( .A1(n_306), .A2(n_385), .A3(n_453), .B1(n_484), .B2(n_485), .C(n_489), .Y(n_483) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_307), .Y(n_382) );
AND2x2_ASAP7_75t_L g407 ( .A(n_307), .B(n_336), .Y(n_407) );
AND2x2_ASAP7_75t_L g482 ( .A(n_307), .B(n_392), .Y(n_482) );
INVx1_ASAP7_75t_L g351 ( .A(n_308), .Y(n_351) );
BUFx2_ASAP7_75t_L g361 ( .A(n_308), .Y(n_361) );
NOR2xp67_ASAP7_75t_L g468 ( .A(n_308), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_SL g406 ( .A(n_309), .Y(n_406) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
BUFx2_ASAP7_75t_L g413 ( .A(n_310), .Y(n_413) );
INVx2_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_311), .Y(n_372) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AOI21xp33_ASAP7_75t_SL g313 ( .A1(n_314), .A2(n_331), .B(n_334), .Y(n_313) );
NOR2xp67_ASAP7_75t_L g465 ( .A(n_314), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_329), .Y(n_315) );
INVx3_ASAP7_75t_L g356 ( .A(n_316), .Y(n_356) );
AND2x2_ASAP7_75t_L g387 ( .A(n_316), .B(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x4_ASAP7_75t_L g344 ( .A(n_317), .B(n_318), .Y(n_344) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_322), .Y(n_556) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_326), .Y(n_555) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g427 ( .A(n_329), .Y(n_427) );
INVx1_ASAP7_75t_SL g512 ( .A(n_330), .Y(n_512) );
INVxp33_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_333), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g438 ( .A(n_333), .B(n_395), .Y(n_438) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
AND2x2_ASAP7_75t_L g442 ( .A(n_335), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_335), .B(n_457), .Y(n_456) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_336), .B(n_373), .Y(n_428) );
NOR4xp25_ASAP7_75t_L g523 ( .A(n_336), .B(n_367), .C(n_524), .D(n_525), .Y(n_523) );
OR2x2_ASAP7_75t_L g491 ( .A(n_337), .B(n_492), .Y(n_491) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_345), .B1(n_350), .B2(n_352), .C(n_357), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AND2x2_ASAP7_75t_L g366 ( .A(n_341), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g403 ( .A(n_342), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g423 ( .A(n_343), .Y(n_423) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g446 ( .A(n_344), .Y(n_446) );
AND2x2_ASAP7_75t_L g453 ( .A(n_344), .B(n_454), .Y(n_453) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
OR2x2_ASAP7_75t_L g390 ( .A(n_347), .B(n_391), .Y(n_390) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_349), .B(n_363), .Y(n_362) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx2_ASAP7_75t_L g367 ( .A(n_354), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_354), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g359 ( .A(n_356), .Y(n_359) );
OAI321xp33_ASAP7_75t_L g471 ( .A1(n_356), .A2(n_464), .A3(n_472), .B1(n_477), .B2(n_479), .C(n_483), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
OR2x2_ASAP7_75t_L g426 ( .A(n_359), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g526 ( .A(n_362), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_363), .B(n_406), .Y(n_405) );
NAND2xp33_ASAP7_75t_SL g506 ( .A(n_363), .B(n_377), .Y(n_506) );
OAI211xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .B(n_379), .C(n_383), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NOR2x1_ASAP7_75t_L g368 ( .A(n_369), .B(n_374), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g475 ( .A(n_372), .Y(n_475) );
INVx3_ASAP7_75t_L g414 ( .A(n_373), .Y(n_414) );
OR2x2_ASAP7_75t_L g517 ( .A(n_373), .B(n_391), .Y(n_517) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_375), .A2(n_459), .B1(n_461), .B2(n_463), .Y(n_458) );
OR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_SL g457 ( .A(n_378), .Y(n_457) );
OR2x2_ASAP7_75t_L g534 ( .A(n_378), .B(n_391), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI21xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_385), .B(n_389), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_387), .B(n_404), .Y(n_503) );
AND2x2_ASAP7_75t_L g509 ( .A(n_387), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g454 ( .A(n_388), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_393), .B1(n_396), .B2(n_398), .Y(n_389) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_391), .A2(n_434), .B(n_436), .C(n_438), .Y(n_435) );
INVx2_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_394), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_394), .B(n_486), .Y(n_508) );
INVx2_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g480 ( .A(n_397), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_399), .A2(n_431), .B(n_434), .C(n_435), .Y(n_430) );
NAND3xp33_ASAP7_75t_SL g400 ( .A(n_401), .B(n_415), .C(n_430), .Y(n_400) );
AOI222xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B1(n_407), .B2(n_408), .C1(n_409), .C2(n_412), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g464 ( .A(n_404), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_404), .B(n_437), .Y(n_490) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g424 ( .A(n_411), .Y(n_424) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
OR2x2_ASAP7_75t_L g529 ( .A(n_413), .B(n_446), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_414), .A2(n_505), .B1(n_507), .B2(n_509), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_421), .B1(n_425), .B2(n_428), .C(n_429), .Y(n_415) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI21xp5_ASAP7_75t_SL g489 ( .A1(n_422), .A2(n_490), .B(n_491), .Y(n_489) );
OR2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx2_ASAP7_75t_L g437 ( .A(n_423), .Y(n_437) );
AND2x2_ASAP7_75t_L g531 ( .A(n_423), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g515 ( .A(n_427), .Y(n_515) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g444 ( .A(n_433), .B(n_434), .Y(n_444) );
INVx1_ASAP7_75t_L g497 ( .A(n_433), .Y(n_497) );
NOR3xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_471), .C(n_493), .Y(n_439) );
OAI211xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_445), .B(n_447), .C(n_452), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI21xp33_ASAP7_75t_L g447 ( .A1(n_442), .A2(n_448), .B(n_449), .Y(n_447) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AOI211xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_455), .B(n_458), .C(n_465), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g476 ( .A(n_459), .Y(n_476) );
INVxp67_ASAP7_75t_SL g501 ( .A(n_460), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_462), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g524 ( .A(n_462), .Y(n_524) );
AND2x2_ASAP7_75t_L g514 ( .A(n_464), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g484 ( .A(n_466), .Y(n_484) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
INVx1_ASAP7_75t_L g492 ( .A(n_468), .Y(n_492) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_476), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_480), .A2(n_514), .B1(n_516), .B2(n_518), .C(n_523), .Y(n_513) );
OAI21xp33_ASAP7_75t_SL g528 ( .A1(n_485), .A2(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND4xp25_ASAP7_75t_L g493 ( .A(n_494), .B(n_504), .C(n_513), .D(n_527), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .B1(n_501), .B2(n_502), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
INVxp67_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_522), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OAI222xp33_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_543), .B1(n_549), .B2(n_551), .C1(n_554), .C2(n_557), .Y(n_539) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
CKINVDCx16_ASAP7_75t_R g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
endmodule