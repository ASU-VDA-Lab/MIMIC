module fake_aes_12715_n_745 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_745);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_745;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g107 ( .A(n_29), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_82), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_18), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_50), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_18), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_9), .Y(n_112) );
INVx4_ASAP7_75t_R g113 ( .A(n_10), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_23), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_8), .B(n_46), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_56), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_62), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_37), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_95), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_105), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_58), .Y(n_121) );
BUFx2_ASAP7_75t_L g122 ( .A(n_66), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_48), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_39), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_99), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_96), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_70), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_34), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_76), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_67), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_36), .Y(n_132) );
INVxp33_ASAP7_75t_SL g133 ( .A(n_71), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_47), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_15), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_78), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_9), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_102), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_92), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_20), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_42), .Y(n_141) );
INVx1_ASAP7_75t_SL g142 ( .A(n_21), .Y(n_142) );
CKINVDCx14_ASAP7_75t_R g143 ( .A(n_30), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_13), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_98), .Y(n_145) );
BUFx10_ASAP7_75t_L g146 ( .A(n_72), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_32), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_4), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_23), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g150 ( .A1(n_137), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_132), .Y(n_151) );
NOR2x1_ASAP7_75t_L g152 ( .A(n_107), .B(n_0), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_132), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_122), .B(n_1), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_132), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_108), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g158 ( .A1(n_137), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_158) );
NOR2xp33_ASAP7_75t_SL g159 ( .A(n_110), .B(n_106), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_148), .Y(n_160) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_120), .A2(n_53), .B(n_103), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_114), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g163 ( .A(n_110), .B(n_25), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_128), .B(n_3), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_125), .A2(n_54), .B(n_101), .Y(n_167) );
OAI22xp5_ASAP7_75t_SL g168 ( .A1(n_144), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_151), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_151), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_155), .B(n_114), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_155), .B(n_146), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_167), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_162), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_155), .B(n_146), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_162), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
AND2x6_ASAP7_75t_L g183 ( .A(n_154), .B(n_129), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_155), .B(n_154), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_155), .B(n_116), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_154), .A2(n_111), .B1(n_135), .B2(n_140), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_157), .B(n_133), .Y(n_189) );
INVx8_ASAP7_75t_L g190 ( .A(n_154), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_154), .Y(n_191) );
NAND3xp33_ASAP7_75t_L g192 ( .A(n_157), .B(n_147), .C(n_145), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_164), .B(n_116), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_164), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_153), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_169), .B(n_138), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_183), .A2(n_165), .B1(n_169), .B2(n_163), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_195), .B(n_165), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_190), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_191), .B(n_165), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_195), .B(n_165), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_177), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_191), .B(n_165), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_191), .B(n_189), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_191), .B(n_160), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_190), .B(n_183), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_184), .B(n_152), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_170), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_190), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_190), .B(n_160), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_177), .B(n_160), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_176), .Y(n_215) );
NAND2xp33_ASAP7_75t_L g216 ( .A(n_183), .B(n_138), .Y(n_216) );
BUFx2_ASAP7_75t_L g217 ( .A(n_190), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_183), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_188), .B(n_159), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_194), .A2(n_112), .B(n_109), .C(n_142), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_183), .A2(n_159), .B1(n_163), .B2(n_168), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_176), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_183), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_172), .B(n_133), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_183), .B(n_152), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_198), .B(n_139), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_175), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_173), .B(n_139), .Y(n_228) );
NOR2xp67_ASAP7_75t_L g229 ( .A(n_192), .B(n_26), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_180), .B(n_119), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_186), .B(n_143), .Y(n_231) );
NOR2xp67_ASAP7_75t_L g232 ( .A(n_192), .B(n_27), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_175), .B(n_167), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_175), .B(n_167), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_171), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_171), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_181), .B(n_167), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_201), .B(n_130), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_208), .B(n_149), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_208), .B(n_130), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_233), .A2(n_167), .B(n_161), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_233), .A2(n_161), .B(n_115), .Y(n_242) );
INVxp67_ASAP7_75t_L g243 ( .A(n_217), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_201), .B(n_136), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_234), .A2(n_161), .B(n_196), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_206), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_205), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_213), .B(n_136), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_234), .A2(n_196), .B(n_193), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_201), .Y(n_250) );
INVx4_ASAP7_75t_L g251 ( .A(n_217), .Y(n_251) );
OAI22xp5_ASAP7_75t_SL g252 ( .A1(n_204), .A2(n_144), .B1(n_158), .B2(n_150), .Y(n_252) );
AO21x1_ASAP7_75t_L g253 ( .A1(n_237), .A2(n_185), .B(n_182), .Y(n_253) );
INVxp67_ASAP7_75t_L g254 ( .A(n_213), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_210), .A2(n_168), .B1(n_150), .B2(n_158), .Y(n_255) );
OR2x6_ASAP7_75t_L g256 ( .A(n_209), .B(n_134), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_205), .A2(n_193), .B(n_178), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_209), .B(n_117), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_210), .B(n_226), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_214), .A2(n_123), .B1(n_131), .B2(n_127), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_237), .A2(n_182), .B(n_185), .C(n_187), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_210), .B(n_118), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_200), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_200), .A2(n_178), .B(n_179), .Y(n_264) );
AOI21xp33_ASAP7_75t_L g265 ( .A1(n_212), .A2(n_124), .B(n_134), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_214), .Y(n_266) );
OAI21xp33_ASAP7_75t_L g267 ( .A1(n_199), .A2(n_187), .B(n_134), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_203), .A2(n_179), .B(n_178), .Y(n_268) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_199), .B(n_134), .C(n_141), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_219), .A2(n_113), .B(n_179), .C(n_7), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_241), .A2(n_227), .B(n_203), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_247), .Y(n_272) );
AO31x2_ASAP7_75t_L g273 ( .A1(n_253), .A2(n_225), .A3(n_215), .B(n_211), .Y(n_273) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_245), .A2(n_227), .B(n_232), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_242), .A2(n_227), .B(n_202), .Y(n_275) );
AOI22x1_ASAP7_75t_L g276 ( .A1(n_263), .A2(n_227), .B1(n_210), .B2(n_215), .Y(n_276) );
INVx5_ASAP7_75t_L g277 ( .A(n_250), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_240), .B(n_224), .Y(n_278) );
AOI21x1_ASAP7_75t_L g279 ( .A1(n_269), .A2(n_232), .B(n_229), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_250), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_254), .A2(n_221), .B1(n_226), .B2(n_212), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g282 ( .A1(n_261), .A2(n_225), .B(n_207), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_251), .B(n_218), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_251), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_249), .A2(n_257), .B(n_259), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_254), .B(n_221), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_248), .A2(n_218), .B1(n_223), .B2(n_207), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_264), .A2(n_268), .B(n_246), .Y(n_288) );
NOR2xp33_ASAP7_75t_R g289 ( .A(n_266), .B(n_216), .Y(n_289) );
NOR2xp67_ASAP7_75t_SL g290 ( .A(n_250), .B(n_223), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_250), .B(n_206), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_267), .A2(n_228), .B(n_231), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_239), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_255), .B(n_231), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_272), .Y(n_295) );
NOR3xp33_ASAP7_75t_L g296 ( .A(n_278), .B(n_252), .C(n_220), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_271), .A2(n_270), .B(n_256), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_293), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_284), .B(n_243), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_294), .B(n_238), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_286), .B(n_243), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_278), .A2(n_255), .B(n_206), .C(n_211), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_277), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_277), .B(n_284), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_281), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_273), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_282), .B(n_211), .Y(n_307) );
INVx8_ASAP7_75t_L g308 ( .A(n_277), .Y(n_308) );
AOI22xp33_ASAP7_75t_SL g309 ( .A1(n_289), .A2(n_256), .B1(n_262), .B2(n_244), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_277), .B(n_258), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_285), .A2(n_256), .B(n_265), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_280), .Y(n_312) );
OA21x2_ASAP7_75t_L g313 ( .A1(n_274), .A2(n_229), .B(n_215), .Y(n_313) );
AOI21x1_ASAP7_75t_L g314 ( .A1(n_274), .A2(n_222), .B(n_236), .Y(n_314) );
AOI22xp33_ASAP7_75t_SL g315 ( .A1(n_289), .A2(n_230), .B1(n_141), .B2(n_222), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_287), .B(n_260), .Y(n_316) );
AND2x6_ASAP7_75t_L g317 ( .A(n_307), .B(n_280), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_300), .B(n_273), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_307), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_314), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_313), .Y(n_321) );
AO21x2_ASAP7_75t_L g322 ( .A1(n_311), .A2(n_288), .B(n_275), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_306), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_295), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_305), .Y(n_325) );
BUFx2_ASAP7_75t_SL g326 ( .A(n_303), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_312), .B(n_273), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_313), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_313), .A2(n_279), .B(n_276), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_312), .Y(n_330) );
BUFx4f_ASAP7_75t_SL g331 ( .A(n_303), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_299), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_312), .B(n_273), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_299), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_302), .B(n_222), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_299), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_301), .B(n_291), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_302), .B(n_291), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_297), .A2(n_292), .B(n_236), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_299), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_304), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_304), .Y(n_342) );
NAND3xp33_ASAP7_75t_L g343 ( .A(n_296), .B(n_141), .C(n_153), .Y(n_343) );
OA21x2_ASAP7_75t_L g344 ( .A1(n_316), .A2(n_235), .B(n_283), .Y(n_344) );
AO21x2_ASAP7_75t_L g345 ( .A1(n_316), .A2(n_235), .B(n_283), .Y(n_345) );
NOR2x1_ASAP7_75t_SL g346 ( .A(n_326), .B(n_308), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_327), .B(n_141), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_323), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_323), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_320), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_320), .Y(n_351) );
INVxp67_ASAP7_75t_SL g352 ( .A(n_344), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_325), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_319), .A2(n_298), .B1(n_309), .B2(n_315), .Y(n_354) );
INVxp67_ASAP7_75t_SL g355 ( .A(n_344), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_319), .B(n_153), .Y(n_356) );
INVx4_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_342), .B(n_308), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_318), .B(n_308), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_332), .Y(n_360) );
BUFx2_ASAP7_75t_L g361 ( .A(n_332), .Y(n_361) );
AO21x2_ASAP7_75t_L g362 ( .A1(n_320), .A2(n_283), .B(n_166), .Y(n_362) );
AO21x2_ASAP7_75t_L g363 ( .A1(n_320), .A2(n_166), .B(n_310), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_336), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_325), .B(n_308), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_327), .B(n_166), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_327), .B(n_166), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_341), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_327), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_327), .B(n_166), .Y(n_370) );
INVxp33_ASAP7_75t_L g371 ( .A(n_342), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_333), .Y(n_372) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_324), .A2(n_5), .B1(n_6), .B2(n_8), .C1(n_10), .C2(n_11), .Y(n_373) );
INVx2_ASAP7_75t_SL g374 ( .A(n_330), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_328), .Y(n_375) );
AO21x2_ASAP7_75t_L g376 ( .A1(n_343), .A2(n_166), .B(n_310), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_333), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_333), .B(n_166), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_318), .B(n_11), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_333), .B(n_166), .Y(n_380) );
NOR2x1_ASAP7_75t_L g381 ( .A(n_341), .B(n_174), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_333), .B(n_61), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_318), .B(n_12), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_324), .B(n_12), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_336), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_328), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_345), .B(n_13), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_340), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_328), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_328), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_345), .B(n_14), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_345), .A2(n_290), .B1(n_15), .B2(n_16), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_345), .A2(n_197), .B1(n_174), .B2(n_17), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_348), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_369), .B(n_345), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_369), .B(n_344), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_383), .B(n_337), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_353), .B(n_344), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_372), .B(n_344), .Y(n_399) );
INVx6_ASAP7_75t_L g400 ( .A(n_357), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_348), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_353), .B(n_344), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_350), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_357), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_349), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_383), .B(n_337), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_372), .B(n_335), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_377), .B(n_335), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_349), .B(n_338), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_368), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_387), .B(n_335), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_377), .B(n_338), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_347), .B(n_338), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_347), .B(n_334), .Y(n_415) );
AND2x2_ASAP7_75t_SL g416 ( .A(n_357), .B(n_340), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_347), .B(n_334), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_347), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_388), .B(n_337), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_375), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_347), .B(n_334), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_375), .Y(n_422) );
INVxp67_ASAP7_75t_SL g423 ( .A(n_371), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_368), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_387), .B(n_322), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_383), .B(n_341), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_371), .B(n_331), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_366), .B(n_322), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_388), .B(n_341), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_366), .B(n_322), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_387), .B(n_322), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_350), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_350), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_366), .B(n_322), .Y(n_434) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_368), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_367), .B(n_321), .Y(n_436) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_373), .B(n_343), .C(n_321), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_360), .B(n_361), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_367), .B(n_321), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_391), .B(n_317), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_367), .B(n_330), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_351), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_351), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_391), .B(n_317), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_370), .B(n_321), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_386), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_370), .B(n_321), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_386), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_370), .B(n_321), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_360), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_386), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_389), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_389), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_351), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_378), .B(n_321), .Y(n_455) );
INVx5_ASAP7_75t_L g456 ( .A(n_357), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_389), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_361), .B(n_326), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_379), .B(n_331), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_378), .B(n_321), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_378), .B(n_330), .Y(n_461) );
OAI21xp33_ASAP7_75t_L g462 ( .A1(n_373), .A2(n_339), .B(n_330), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_390), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_380), .B(n_330), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_390), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_428), .B(n_380), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_404), .B(n_357), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_394), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_450), .Y(n_469) );
OR2x6_ASAP7_75t_L g470 ( .A(n_400), .B(n_382), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_394), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_401), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_438), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_438), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_456), .B(n_382), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_401), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_463), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_428), .B(n_380), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_419), .B(n_352), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_462), .A2(n_354), .B1(n_317), .B2(n_359), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_430), .B(n_434), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_458), .Y(n_482) );
NAND5xp2_ASAP7_75t_L g483 ( .A(n_462), .B(n_354), .C(n_392), .D(n_393), .E(n_358), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_405), .B(n_379), .Y(n_484) );
INVxp33_ASAP7_75t_L g485 ( .A(n_458), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_430), .B(n_352), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_405), .Y(n_487) );
NAND3xp33_ASAP7_75t_L g488 ( .A(n_437), .B(n_393), .C(n_392), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_397), .B(n_385), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_429), .Y(n_490) );
NOR2xp33_ASAP7_75t_R g491 ( .A(n_416), .B(n_358), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_419), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_434), .B(n_355), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_406), .B(n_385), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_425), .B(n_355), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_412), .B(n_356), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_436), .B(n_390), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_436), .B(n_364), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_409), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_439), .B(n_364), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_439), .B(n_364), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_409), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_445), .B(n_374), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_429), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_445), .B(n_374), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_425), .B(n_431), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_447), .B(n_374), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_463), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_447), .B(n_362), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_412), .B(n_356), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_463), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_403), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_398), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_459), .B(n_384), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_449), .B(n_362), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_449), .B(n_362), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_411), .B(n_356), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_424), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_455), .B(n_362), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_398), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_455), .B(n_382), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_402), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_404), .B(n_382), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_456), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_402), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_431), .B(n_359), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_413), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_411), .B(n_359), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_426), .B(n_363), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_423), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_407), .B(n_384), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_413), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_460), .B(n_382), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_460), .B(n_363), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_407), .B(n_408), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_420), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_420), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_422), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_408), .B(n_365), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_395), .B(n_365), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_456), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_414), .B(n_363), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_422), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_395), .B(n_363), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_403), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_414), .B(n_339), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_396), .B(n_339), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_446), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_396), .B(n_346), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_399), .B(n_346), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_446), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_399), .B(n_317), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_473), .Y(n_553) );
OAI21xp5_ASAP7_75t_SL g554 ( .A1(n_480), .A2(n_427), .B(n_437), .Y(n_554) );
INVxp67_ASAP7_75t_SL g555 ( .A(n_518), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_482), .Y(n_556) );
NAND2x1_ASAP7_75t_L g557 ( .A(n_470), .B(n_400), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_474), .Y(n_558) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_488), .A2(n_416), .B(n_418), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_477), .Y(n_560) );
O2A1O1Ixp33_ASAP7_75t_L g561 ( .A1(n_483), .A2(n_440), .B(n_444), .C(n_404), .Y(n_561) );
OAI21xp33_ASAP7_75t_L g562 ( .A1(n_485), .A2(n_444), .B(n_440), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_492), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_481), .B(n_461), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_469), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_468), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_471), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_481), .B(n_461), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_472), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_514), .A2(n_531), .B1(n_416), .B2(n_502), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_476), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_477), .Y(n_572) );
INVx2_ASAP7_75t_SL g573 ( .A(n_490), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_470), .A2(n_456), .B1(n_400), .B2(n_404), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_513), .B(n_448), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_487), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_508), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_508), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_499), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_535), .B(n_400), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_504), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_506), .B(n_448), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_491), .Y(n_583) );
INVxp33_ASAP7_75t_L g584 ( .A(n_491), .Y(n_584) );
NAND2x1p5_ASAP7_75t_L g585 ( .A(n_524), .B(n_456), .Y(n_585) );
NAND2x1_ASAP7_75t_L g586 ( .A(n_470), .B(n_400), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_520), .B(n_451), .Y(n_587) );
OAI21xp33_ASAP7_75t_SL g588 ( .A1(n_524), .A2(n_541), .B(n_470), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_522), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_525), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_506), .B(n_451), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_526), .B(n_452), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_511), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_495), .B(n_452), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_SL g595 ( .A1(n_530), .A2(n_465), .B(n_453), .C(n_457), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_527), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_466), .B(n_478), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_466), .B(n_464), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_532), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_536), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_537), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_538), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_511), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_526), .B(n_453), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_495), .B(n_457), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_549), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_543), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_548), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_551), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_479), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_479), .B(n_465), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_486), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_541), .B(n_456), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_486), .B(n_403), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_540), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_493), .B(n_432), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_478), .B(n_464), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_539), .Y(n_618) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_512), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_550), .Y(n_620) );
OAI21xp33_ASAP7_75t_L g621 ( .A1(n_485), .A2(n_435), .B(n_415), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_493), .B(n_454), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g623 ( .A1(n_475), .A2(n_410), .B1(n_441), .B2(n_442), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_498), .B(n_415), .Y(n_624) );
NAND4xp25_ASAP7_75t_SL g625 ( .A(n_528), .B(n_421), .C(n_417), .D(n_381), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_497), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_498), .B(n_417), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_512), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_497), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_484), .B(n_454), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_591), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_581), .B(n_489), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_606), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g634 ( .A1(n_584), .A2(n_475), .B1(n_523), .B2(n_552), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_595), .A2(n_467), .B(n_523), .Y(n_635) );
OAI322xp33_ASAP7_75t_L g636 ( .A1(n_583), .A2(n_494), .A3(n_517), .B1(n_496), .B2(n_510), .C1(n_529), .C2(n_544), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_591), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_620), .Y(n_638) );
NOR4xp25_ASAP7_75t_SL g639 ( .A(n_554), .B(n_467), .C(n_523), .D(n_410), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_565), .B(n_500), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_555), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_561), .A2(n_500), .B1(n_501), .B2(n_546), .C(n_542), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_610), .B(n_545), .Y(n_643) );
AOI321xp33_ASAP7_75t_L g644 ( .A1(n_561), .A2(n_546), .A3(n_542), .B1(n_547), .B2(n_533), .C(n_521), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_612), .B(n_529), .Y(n_645) );
AOI322xp5_ASAP7_75t_L g646 ( .A1(n_588), .A2(n_501), .A3(n_547), .B1(n_509), .B2(n_519), .C1(n_516), .C2(n_515), .Y(n_646) );
AOI21xp33_ASAP7_75t_SL g647 ( .A1(n_585), .A2(n_467), .B(n_519), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_594), .Y(n_648) );
OAI222xp33_ASAP7_75t_L g649 ( .A1(n_570), .A2(n_521), .B1(n_533), .B2(n_515), .C1(n_509), .C2(n_516), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_594), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_559), .A2(n_534), .B1(n_410), .B2(n_507), .Y(n_651) );
OAI32xp33_ASAP7_75t_L g652 ( .A1(n_585), .A2(n_534), .A3(n_507), .B1(n_505), .B2(n_503), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_625), .A2(n_441), .B1(n_421), .B2(n_503), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_614), .B(n_505), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_589), .B(n_545), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_559), .A2(n_441), .B1(n_317), .B2(n_442), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_614), .B(n_454), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_605), .Y(n_658) );
OAI21xp33_ASAP7_75t_L g659 ( .A1(n_621), .A2(n_441), .B(n_442), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_618), .A2(n_443), .B1(n_433), .B2(n_432), .C(n_330), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_615), .B(n_14), .Y(n_661) );
INVx2_ASAP7_75t_SL g662 ( .A(n_573), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_605), .Y(n_663) );
INVxp67_ASAP7_75t_SL g664 ( .A(n_555), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_575), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_575), .Y(n_666) );
OAI211xp5_ASAP7_75t_L g667 ( .A1(n_557), .A2(n_381), .B(n_433), .C(n_432), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_587), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_613), .A2(n_317), .B(n_433), .Y(n_669) );
OAI322xp33_ASAP7_75t_L g670 ( .A1(n_553), .A2(n_443), .A3(n_17), .B1(n_19), .B2(n_20), .C1(n_21), .C2(n_22), .Y(n_670) );
XOR2xp5_ASAP7_75t_L g671 ( .A(n_625), .B(n_16), .Y(n_671) );
OAI21xp5_ASAP7_75t_SL g672 ( .A1(n_574), .A2(n_443), .B(n_330), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_560), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_587), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_590), .B(n_376), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_586), .A2(n_330), .B1(n_22), .B2(n_24), .C(n_19), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_564), .B(n_376), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_574), .A2(n_317), .B1(n_376), .B2(n_24), .Y(n_678) );
NAND2xp33_ASAP7_75t_SL g679 ( .A(n_597), .B(n_376), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_568), .B(n_317), .Y(n_680) );
AOI31xp33_ASAP7_75t_L g681 ( .A1(n_671), .A2(n_623), .A3(n_580), .B(n_558), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_631), .B(n_563), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_636), .A2(n_579), .B1(n_562), .B2(n_571), .C(n_576), .Y(n_683) );
OAI22xp5_ASAP7_75t_SL g684 ( .A1(n_633), .A2(n_556), .B1(n_619), .B2(n_616), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_642), .A2(n_629), .B1(n_626), .B2(n_616), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_651), .A2(n_622), .B1(n_566), .B2(n_567), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_639), .A2(n_619), .B(n_630), .Y(n_687) );
OAI221xp5_ASAP7_75t_SL g688 ( .A1(n_646), .A2(n_622), .B1(n_592), .B2(n_604), .C(n_582), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g689 ( .A1(n_651), .A2(n_569), .B1(n_600), .B2(n_596), .C1(n_599), .C2(n_601), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_637), .B(n_598), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_662), .A2(n_617), .B1(n_602), .B2(n_607), .Y(n_691) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_664), .A2(n_630), .B(n_608), .C(n_609), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_647), .B(n_611), .Y(n_693) );
AO22x1_ASAP7_75t_L g694 ( .A1(n_641), .A2(n_627), .B1(n_624), .B2(n_317), .Y(n_694) );
OAI21xp33_ASAP7_75t_SL g695 ( .A1(n_653), .A2(n_628), .B(n_603), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_649), .A2(n_652), .B1(n_670), .B2(n_650), .C(n_658), .Y(n_696) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_644), .A2(n_593), .B1(n_578), .B2(n_577), .C(n_572), .Y(n_697) );
NAND4xp25_ASAP7_75t_L g698 ( .A(n_661), .B(n_28), .C(n_31), .D(n_33), .Y(n_698) );
OA21x2_ASAP7_75t_SL g699 ( .A1(n_638), .A2(n_329), .B(n_38), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_634), .A2(n_329), .B1(n_197), .B2(n_174), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_659), .A2(n_197), .B1(n_174), .B2(n_329), .C(n_43), .Y(n_701) );
AOI32xp33_ASAP7_75t_L g702 ( .A1(n_679), .A2(n_35), .A3(n_40), .B1(n_41), .B2(n_44), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_632), .B(n_45), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_665), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_635), .A2(n_197), .B(n_174), .Y(n_705) );
AOI22x1_ASAP7_75t_L g706 ( .A1(n_669), .A2(n_49), .B1(n_51), .B2(n_52), .Y(n_706) );
AOI311xp33_ASAP7_75t_L g707 ( .A1(n_640), .A2(n_55), .A3(n_57), .B(n_59), .C(n_60), .Y(n_707) );
AOI322xp5_ASAP7_75t_L g708 ( .A1(n_648), .A2(n_63), .A3(n_64), .B1(n_65), .B2(n_68), .C1(n_69), .C2(n_73), .Y(n_708) );
INVxp67_ASAP7_75t_L g709 ( .A(n_666), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g710 ( .A(n_676), .B(n_197), .C(n_75), .Y(n_710) );
OAI21xp5_ASAP7_75t_SL g711 ( .A1(n_672), .A2(n_74), .B(n_77), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_663), .B(n_79), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_668), .Y(n_713) );
AOI221x1_ASAP7_75t_SL g714 ( .A1(n_674), .A2(n_678), .B1(n_643), .B2(n_655), .C(n_675), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_678), .A2(n_80), .B(n_81), .Y(n_715) );
OAI211xp5_ASAP7_75t_SL g716 ( .A1(n_656), .A2(n_84), .B(n_85), .C(n_86), .Y(n_716) );
NOR4xp25_ASAP7_75t_L g717 ( .A(n_667), .B(n_87), .C(n_88), .D(n_89), .Y(n_717) );
NAND5xp2_ASAP7_75t_L g718 ( .A(n_660), .B(n_90), .C(n_91), .D(n_93), .E(n_94), .Y(n_718) );
OAI211xp5_ASAP7_75t_SL g719 ( .A1(n_645), .A2(n_97), .B(n_100), .C(n_104), .Y(n_719) );
OAI32xp33_ASAP7_75t_L g720 ( .A1(n_654), .A2(n_657), .A3(n_643), .B1(n_680), .B2(n_655), .Y(n_720) );
AOI21xp33_ASAP7_75t_L g721 ( .A1(n_675), .A2(n_677), .B(n_673), .Y(n_721) );
NOR2xp67_ASAP7_75t_L g722 ( .A(n_687), .B(n_695), .Y(n_722) );
NAND3x1_ASAP7_75t_L g723 ( .A(n_705), .B(n_683), .C(n_696), .Y(n_723) );
NAND4xp25_ASAP7_75t_SL g724 ( .A(n_683), .B(n_689), .C(n_685), .D(n_686), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_681), .B(n_688), .Y(n_725) );
NOR2xp67_ASAP7_75t_SL g726 ( .A(n_710), .B(n_711), .Y(n_726) );
NAND3xp33_ASAP7_75t_SL g727 ( .A(n_717), .B(n_702), .C(n_715), .Y(n_727) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_707), .B(n_708), .C(n_703), .Y(n_728) );
NAND4xp25_ASAP7_75t_L g729 ( .A(n_725), .B(n_699), .C(n_714), .D(n_698), .Y(n_729) );
NOR2x1_ASAP7_75t_L g730 ( .A(n_727), .B(n_719), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_723), .Y(n_731) );
NAND3xp33_ASAP7_75t_L g732 ( .A(n_722), .B(n_692), .C(n_709), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_731), .Y(n_733) );
NOR3xp33_ASAP7_75t_L g734 ( .A(n_730), .B(n_724), .C(n_728), .Y(n_734) );
NOR2x1_ASAP7_75t_L g735 ( .A(n_729), .B(n_693), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_734), .B(n_732), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_733), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_737), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_736), .A2(n_735), .B1(n_726), .B2(n_684), .Y(n_739) );
OAI22x1_ASAP7_75t_L g740 ( .A1(n_738), .A2(n_706), .B1(n_691), .B2(n_700), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_739), .A2(n_713), .B1(n_704), .B2(n_712), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_741), .A2(n_694), .B1(n_690), .B2(n_682), .Y(n_742) );
AOI21xp33_ASAP7_75t_SL g743 ( .A1(n_742), .A2(n_740), .B(n_720), .Y(n_743) );
OAI21xp5_ASAP7_75t_L g744 ( .A1(n_743), .A2(n_721), .B(n_701), .Y(n_744) );
O2A1O1Ixp33_ASAP7_75t_L g745 ( .A1(n_744), .A2(n_697), .B(n_716), .C(n_718), .Y(n_745) );
endmodule