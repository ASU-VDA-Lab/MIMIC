module fake_netlist_6_3520_n_2020 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2020);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2020;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_202),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_77),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_30),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_193),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_30),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_31),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_45),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_29),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_161),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_22),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_116),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_46),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_134),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_0),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_87),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_113),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_70),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_200),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_111),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_43),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_107),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_184),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_25),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_178),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_142),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_88),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_90),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_137),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_148),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_58),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_3),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_41),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_50),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_175),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_103),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_59),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_163),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_99),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_187),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_192),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_34),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_106),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_171),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_164),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_181),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_143),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_162),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_194),
.Y(n_266)
);

BUFx8_ASAP7_75t_SL g267 ( 
.A(n_196),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_18),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_96),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_149),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_51),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_179),
.Y(n_273)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_158),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_75),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_191),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_70),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_83),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_97),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_45),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_114),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_51),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_41),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_131),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_44),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_133),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_49),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_183),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_78),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_159),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_132),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_118),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_29),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_0),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_152),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_25),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_147),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_141),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_3),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_65),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_32),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_166),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_5),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_61),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_204),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_136),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_110),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_15),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_125),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_112),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_20),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_39),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_169),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_92),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_109),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_210),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_122),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_89),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_95),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_85),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_105),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_81),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_128),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_207),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_59),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_71),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_82),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_119),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_79),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_129),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_138),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_151),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_13),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_57),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_102),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_27),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_145),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_71),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_11),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_127),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_201),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_55),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_115),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_208),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_173),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_21),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_176),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_76),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_120),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_64),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_50),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_60),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_140),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_123),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_117),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_189),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_165),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_172),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_121),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_100),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_75),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_69),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_52),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_62),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_61),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_6),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_68),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_73),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_2),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_74),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_62),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_156),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_26),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_84),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_33),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_33),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_32),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_135),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_48),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_209),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_31),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_76),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_36),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_8),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_6),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_139),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_130),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_211),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_65),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_86),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_124),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_15),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_80),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_10),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_66),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_60),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_205),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_23),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_35),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_63),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_94),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_57),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_126),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_182),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_53),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_91),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_154),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_34),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_58),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_43),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_104),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_174),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_12),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_10),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_168),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_98),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_195),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_12),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_197),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_216),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_267),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_223),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_392),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_392),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_221),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_214),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_214),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_213),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_212),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_220),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_220),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_228),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_225),
.B(n_1),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_215),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_238),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_222),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_228),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_225),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_274),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_227),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_245),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_245),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_229),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_247),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_247),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_405),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_230),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_232),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_383),
.B(n_1),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_256),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_233),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_307),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_265),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_405),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_251),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_251),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_277),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_289),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_277),
.B(n_2),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_235),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_307),
.B(n_401),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_396),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_313),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_401),
.B(n_4),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_241),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_317),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_282),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_249),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_218),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_253),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_337),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_219),
.Y(n_474)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_396),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_231),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_282),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_359),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_293),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_254),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_330),
.B(n_4),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_403),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_293),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_301),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_255),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_319),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_260),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_263),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_301),
.B(n_5),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_333),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_334),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_334),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_234),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_266),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_336),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_250),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_259),
.B(n_261),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_269),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_336),
.B(n_7),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_338),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_270),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_273),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_237),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_276),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_258),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_338),
.B(n_7),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_274),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_278),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_281),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_250),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_363),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_371),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_288),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_371),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_373),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_290),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_259),
.B(n_261),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_217),
.B(n_8),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_284),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_291),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_295),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_373),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_375),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_302),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_431),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_486),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_R g528 ( 
.A(n_423),
.B(n_305),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_463),
.A2(n_226),
.B1(n_224),
.B2(n_339),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_436),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_498),
.B(n_341),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_518),
.B(n_419),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_486),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_486),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_422),
.B(n_437),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_486),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_486),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_428),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_471),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_438),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_442),
.Y(n_541)
);

INVxp67_ASAP7_75t_SL g542 ( 
.A(n_516),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_428),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_429),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_452),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_429),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_445),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_432),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_449),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_450),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_455),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_432),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_433),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_487),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_441),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_433),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_453),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_434),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_434),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_460),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_462),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_441),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_467),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_508),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_508),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_470),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_472),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_511),
.B(n_284),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_480),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_465),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_485),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_439),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_420),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_468),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_488),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_420),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_421),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_439),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_443),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_421),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_474),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_443),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_444),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_444),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_425),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_495),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_425),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_506),
.B(n_258),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_497),
.Y(n_589)
);

INVxp67_ASAP7_75t_SL g590 ( 
.A(n_461),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_426),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_499),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_520),
.B(n_309),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_502),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_426),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_446),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_446),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_447),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_447),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_457),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_494),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_473),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_478),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_482),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_519),
.B(n_318),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_457),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_503),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_497),
.B(n_335),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_458),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_505),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_509),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_531),
.A2(n_590),
.B1(n_500),
.B2(n_605),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_562),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_536),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_536),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_531),
.B(n_435),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_536),
.Y(n_617)
);

NOR2x1p5_ASAP7_75t_L g618 ( 
.A(n_590),
.B(n_440),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_605),
.A2(n_454),
.B1(n_466),
.B2(n_481),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_532),
.B(n_514),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_536),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_536),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_532),
.B(n_593),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_593),
.B(n_246),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_562),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_538),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_589),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_L g628 ( 
.A(n_599),
.B(n_274),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_589),
.B(n_335),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_562),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_589),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_538),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_608),
.B(n_500),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_608),
.B(n_461),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_608),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_543),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_526),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_530),
.B(n_522),
.Y(n_638)
);

BUFx4f_ASAP7_75t_L g639 ( 
.A(n_599),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_540),
.B(n_430),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_599),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_599),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_541),
.B(n_427),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_543),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_599),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_539),
.A2(n_510),
.B1(n_517),
.B2(n_489),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_568),
.A2(n_448),
.B1(n_424),
.B2(n_456),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_547),
.B(n_521),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_568),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_539),
.A2(n_364),
.B1(n_300),
.B2(n_427),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_599),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_599),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_555),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_588),
.B(n_490),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_536),
.Y(n_655)
);

OAI21xp33_ASAP7_75t_SL g656 ( 
.A1(n_542),
.A2(n_451),
.B(n_490),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_555),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_536),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_545),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_544),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_546),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_568),
.B(n_246),
.Y(n_662)
);

INVx4_ASAP7_75t_SL g663 ( 
.A(n_537),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_L g664 ( 
.A(n_609),
.B(n_274),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_555),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_549),
.B(n_525),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_546),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_548),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_SL g669 ( 
.A(n_554),
.B(n_507),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_537),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_537),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_548),
.B(n_217),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_550),
.B(n_475),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_537),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_557),
.B(n_279),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_542),
.B(n_476),
.Y(n_676)
);

OAI22xp33_ASAP7_75t_L g677 ( 
.A1(n_581),
.A2(n_507),
.B1(n_448),
.B2(n_248),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_552),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_552),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_561),
.B(n_464),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_555),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_563),
.B(n_504),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_553),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_551),
.Y(n_684)
);

CKINVDCx16_ASAP7_75t_R g685 ( 
.A(n_560),
.Y(n_685)
);

NAND2x1p5_ASAP7_75t_L g686 ( 
.A(n_609),
.B(n_412),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_537),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_564),
.B(n_321),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_553),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_554),
.B(n_476),
.Y(n_690)
);

BUFx6f_ASAP7_75t_SL g691 ( 
.A(n_556),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_566),
.B(n_279),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_564),
.B(n_327),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_556),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_570),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_567),
.B(n_298),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_609),
.B(n_274),
.Y(n_697)
);

XOR2x2_ASAP7_75t_SL g698 ( 
.A(n_529),
.B(n_375),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_558),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_609),
.A2(n_379),
.B1(n_381),
.B2(n_382),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_569),
.B(n_244),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_537),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_537),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_564),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_571),
.B(n_298),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_575),
.B(n_315),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_586),
.B(n_257),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_564),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_565),
.Y(n_709)
);

INVx5_ASAP7_75t_L g710 ( 
.A(n_565),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_592),
.Y(n_711)
);

AND2x6_ASAP7_75t_L g712 ( 
.A(n_559),
.B(n_315),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_534),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_565),
.B(n_331),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_559),
.B(n_236),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_572),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_528),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_572),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_534),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_SL g720 ( 
.A(n_594),
.B(n_285),
.Y(n_720)
);

NAND2x1p5_ASAP7_75t_L g721 ( 
.A(n_578),
.B(n_236),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_534),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_579),
.B(n_458),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_607),
.B(n_268),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_579),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_534),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_582),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_565),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_591),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_582),
.B(n_239),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_591),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_583),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_581),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_583),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_535),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_610),
.B(n_271),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_584),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_527),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_527),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_584),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_527),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_596),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_596),
.A2(n_598),
.B1(n_600),
.B2(n_597),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_533),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_611),
.B(n_275),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_597),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_591),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_533),
.B(n_332),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_535),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_533),
.B(n_340),
.Y(n_750)
);

AND2x6_ASAP7_75t_L g751 ( 
.A(n_598),
.B(n_316),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_600),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_601),
.B(n_459),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_606),
.B(n_343),
.Y(n_754)
);

BUFx10_ASAP7_75t_L g755 ( 
.A(n_601),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_606),
.B(n_344),
.Y(n_756)
);

NAND3xp33_ASAP7_75t_L g757 ( 
.A(n_580),
.B(n_283),
.C(n_280),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_580),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_580),
.B(n_345),
.Y(n_759)
);

AND2x2_ASAP7_75t_SL g760 ( 
.A(n_573),
.B(n_316),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_627),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_613),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_613),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_649),
.B(n_459),
.Y(n_764)
);

O2A1O1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_616),
.A2(n_385),
.B(n_394),
.C(n_398),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_623),
.B(n_585),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_649),
.B(n_585),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_748),
.A2(n_576),
.B(n_573),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_726),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_625),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_616),
.B(n_294),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_726),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_619),
.A2(n_529),
.B1(n_387),
.B2(n_388),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_750),
.A2(n_576),
.B(n_573),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_723),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_713),
.A2(n_577),
.B(n_576),
.Y(n_776)
);

AND2x6_ASAP7_75t_SL g777 ( 
.A(n_682),
.B(n_409),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_662),
.A2(n_409),
.B(n_413),
.C(n_366),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_723),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_726),
.Y(n_780)
);

NAND2x1p5_ASAP7_75t_L g781 ( 
.A(n_635),
.B(n_239),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_620),
.B(n_585),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_625),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_630),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_676),
.B(n_296),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_612),
.B(n_319),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_635),
.A2(n_323),
.B1(n_356),
.B2(n_353),
.Y(n_787)
);

NAND3xp33_ASAP7_75t_L g788 ( 
.A(n_676),
.B(n_303),
.C(n_299),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_618),
.A2(n_355),
.B1(n_358),
.B2(n_386),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_753),
.B(n_308),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_633),
.B(n_585),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_733),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_633),
.B(n_591),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_633),
.B(n_591),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_760),
.B(n_686),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_760),
.B(n_591),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_686),
.A2(n_323),
.B1(n_353),
.B2(n_374),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_726),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_716),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_630),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_753),
.B(n_311),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_626),
.B(n_591),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_632),
.B(n_240),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_727),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_636),
.B(n_240),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_644),
.B(n_242),
.Y(n_806)
);

NAND3xp33_ASAP7_75t_L g807 ( 
.A(n_656),
.B(n_325),
.C(n_312),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_629),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_660),
.B(n_242),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_634),
.A2(n_324),
.B1(n_349),
.B2(n_347),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_SL g811 ( 
.A1(n_654),
.A2(n_324),
.B1(n_349),
.B2(n_347),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_661),
.B(n_243),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_667),
.B(n_243),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_727),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_675),
.B(n_326),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_624),
.A2(n_413),
.B1(n_368),
.B2(n_356),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_634),
.B(n_469),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_654),
.B(n_252),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_728),
.B(n_319),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_668),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_678),
.B(n_252),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_679),
.B(n_262),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_683),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_728),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_689),
.B(n_262),
.Y(n_825)
);

NOR2x1p5_ASAP7_75t_L g826 ( 
.A(n_717),
.B(n_342),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_694),
.B(n_264),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_699),
.B(n_264),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_672),
.A2(n_328),
.B(n_397),
.C(n_314),
.Y(n_829)
);

INVx8_ASAP7_75t_L g830 ( 
.A(n_691),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_758),
.B(n_319),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_718),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_713),
.A2(n_587),
.B(n_577),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_725),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_732),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_734),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_690),
.B(n_469),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_669),
.A2(n_357),
.B1(n_390),
.B2(n_416),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_738),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_713),
.A2(n_587),
.B(n_577),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_737),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_624),
.A2(n_310),
.B1(n_314),
.B2(n_329),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_740),
.B(n_286),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_629),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_742),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_746),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_627),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_752),
.B(n_286),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_629),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_662),
.B(n_759),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_672),
.Y(n_851)
);

OAI21xp33_ASAP7_75t_L g852 ( 
.A1(n_654),
.A2(n_647),
.B(n_634),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_675),
.B(n_346),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_688),
.B(n_297),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_653),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_693),
.B(n_297),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_653),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_714),
.B(n_306),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_659),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_754),
.B(n_306),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_719),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_756),
.B(n_310),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_634),
.B(n_477),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_719),
.B(n_328),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_672),
.A2(n_730),
.B(n_715),
.C(n_669),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_692),
.B(n_350),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_755),
.B(n_477),
.Y(n_867)
);

NAND2xp33_ASAP7_75t_L g868 ( 
.A(n_712),
.B(n_751),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_657),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_715),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_657),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_717),
.B(n_320),
.Y(n_872)
);

INVx8_ASAP7_75t_L g873 ( 
.A(n_691),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_719),
.B(n_329),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_722),
.B(n_374),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_641),
.B(n_320),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_641),
.B(n_320),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_755),
.B(n_479),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_642),
.B(n_320),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_665),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_755),
.B(n_479),
.Y(n_881)
);

AOI221xp5_ASAP7_75t_L g882 ( 
.A1(n_677),
.A2(n_287),
.B1(n_304),
.B2(n_348),
.C(n_352),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_722),
.B(n_378),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_665),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_722),
.B(n_378),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_715),
.Y(n_886)
);

INVx8_ASAP7_75t_L g887 ( 
.A(n_691),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_681),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_730),
.B(n_380),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_730),
.B(n_380),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_743),
.B(n_397),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_721),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_642),
.B(n_320),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_701),
.B(n_414),
.C(n_361),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_681),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_690),
.Y(n_896)
);

AND2x6_ASAP7_75t_L g897 ( 
.A(n_645),
.B(n_651),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_645),
.B(n_274),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_721),
.B(n_404),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_651),
.B(n_274),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_692),
.B(n_351),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_664),
.A2(n_417),
.B1(n_415),
.B2(n_404),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_704),
.B(n_415),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_654),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_704),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_631),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_708),
.B(n_417),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_708),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_652),
.B(n_274),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_652),
.B(n_274),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_696),
.A2(n_411),
.B1(n_393),
.B2(n_391),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_696),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_709),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_720),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_707),
.Y(n_915)
);

AOI22x1_ASAP7_75t_L g916 ( 
.A1(n_729),
.A2(n_322),
.B1(n_292),
.B2(n_272),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_709),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_614),
.B(n_587),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_614),
.B(n_595),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_614),
.B(n_595),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_664),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_615),
.B(n_595),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_739),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_705),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_659),
.Y(n_925)
);

AOI221xp5_ASAP7_75t_L g926 ( 
.A1(n_650),
.A2(n_369),
.B1(n_410),
.B2(n_370),
.C(n_362),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_705),
.B(n_706),
.Y(n_927)
);

NAND3xp33_ASAP7_75t_L g928 ( 
.A(n_724),
.B(n_377),
.C(n_367),
.Y(n_928)
);

O2A1O1Ixp5_ASAP7_75t_L g929 ( 
.A1(n_786),
.A2(n_706),
.B(n_639),
.C(n_745),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_915),
.B(n_638),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_786),
.A2(n_697),
.B(n_757),
.C(n_628),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_861),
.A2(n_639),
.B(n_697),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_867),
.B(n_736),
.Y(n_933)
);

AOI21x1_ASAP7_75t_L g934 ( 
.A1(n_819),
.A2(n_731),
.B(n_729),
.Y(n_934)
);

AOI21x1_ASAP7_75t_L g935 ( 
.A1(n_819),
.A2(n_747),
.B(n_731),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_861),
.A2(n_639),
.B(n_628),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_SL g937 ( 
.A(n_792),
.B(n_637),
.Y(n_937)
);

CKINVDCx8_ASAP7_75t_R g938 ( 
.A(n_830),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_847),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_878),
.B(n_637),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_861),
.B(n_637),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_766),
.B(n_673),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_824),
.A2(n_747),
.B(n_687),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_921),
.A2(n_646),
.B1(n_648),
.B2(n_666),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_824),
.A2(n_622),
.B(n_670),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_795),
.A2(n_680),
.B1(n_640),
.B2(n_700),
.Y(n_946)
);

NOR2xp67_ASAP7_75t_L g947 ( 
.A(n_894),
.B(n_739),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_912),
.B(n_711),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_896),
.B(n_574),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_769),
.A2(n_687),
.B(n_622),
.Y(n_950)
);

NOR2xp67_ASAP7_75t_L g951 ( 
.A(n_928),
.B(n_739),
.Y(n_951)
);

OAI321xp33_ASAP7_75t_L g952 ( 
.A1(n_771),
.A2(n_698),
.A3(n_491),
.B1(n_483),
.B2(n_484),
.C(n_492),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_814),
.B(n_764),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_769),
.A2(n_670),
.B(n_622),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_762),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_762),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_771),
.A2(n_643),
.B(n_741),
.C(n_744),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_924),
.B(n_711),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_927),
.A2(n_751),
.B1(n_712),
.B2(n_711),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_892),
.B(n_698),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_847),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_772),
.A2(n_674),
.B(n_617),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_852),
.B(n_602),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_881),
.B(n_785),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_796),
.A2(n_674),
.B(n_617),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_850),
.A2(n_658),
.B(n_702),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_820),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_795),
.A2(n_751),
.B1(n_712),
.B2(n_604),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_820),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_791),
.A2(n_658),
.B(n_655),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_897),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_772),
.A2(n_658),
.B(n_702),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_847),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_780),
.A2(n_655),
.B(n_702),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_835),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_780),
.A2(n_655),
.B(n_621),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_815),
.A2(n_866),
.B(n_901),
.C(n_853),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_865),
.A2(n_741),
.B(n_744),
.C(n_523),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_835),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_914),
.B(n_685),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_815),
.A2(n_741),
.B(n_621),
.C(n_354),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_785),
.B(n_603),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_865),
.A2(n_484),
.B(n_491),
.C(n_492),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_780),
.A2(n_703),
.B(n_671),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_782),
.A2(n_751),
.B(n_712),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_851),
.A2(n_751),
.B1(n_712),
.B2(n_407),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_808),
.B(n_360),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_790),
.B(n_735),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_763),
.Y(n_989)
);

NOR2x1_ASAP7_75t_L g990 ( 
.A(n_826),
.B(n_684),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_767),
.A2(n_751),
.B(n_712),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_798),
.A2(n_703),
.B(n_671),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_836),
.B(n_841),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_859),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_847),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_770),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_870),
.A2(n_406),
.B1(n_738),
.B2(n_671),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_798),
.A2(n_794),
.B(n_793),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_798),
.A2(n_703),
.B(n_671),
.Y(n_999)
);

BUFx4f_ASAP7_75t_L g1000 ( 
.A(n_830),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_864),
.A2(n_703),
.B(n_671),
.Y(n_1001)
);

AO21x1_ASAP7_75t_L g1002 ( 
.A1(n_811),
.A2(n_501),
.B(n_524),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_886),
.A2(n_902),
.B1(n_781),
.B2(n_844),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_906),
.B(n_749),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_849),
.A2(n_738),
.B1(n_695),
.B2(n_684),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_902),
.A2(n_738),
.B1(n_389),
.B2(n_384),
.Y(n_1006)
);

NOR3xp33_ASAP7_75t_L g1007 ( 
.A(n_882),
.B(n_395),
.C(n_399),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_841),
.B(n_710),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_853),
.A2(n_402),
.B(n_365),
.C(n_408),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_874),
.A2(n_710),
.B(n_663),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_845),
.B(n_710),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_875),
.A2(n_710),
.B(n_663),
.Y(n_1012)
);

AO21x1_ASAP7_75t_L g1013 ( 
.A1(n_810),
.A2(n_524),
.B(n_523),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_807),
.A2(n_695),
.B1(n_710),
.B2(n_258),
.Y(n_1014)
);

AOI21x1_ASAP7_75t_L g1015 ( 
.A1(n_776),
.A2(n_501),
.B(n_515),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_817),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_883),
.A2(n_663),
.B(n_515),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_863),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_829),
.A2(n_513),
.B(n_512),
.C(n_496),
.Y(n_1019)
);

NAND3xp33_ASAP7_75t_L g1020 ( 
.A(n_926),
.B(n_400),
.C(n_418),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_833),
.A2(n_513),
.B(n_512),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_845),
.B(n_663),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_885),
.A2(n_868),
.B(n_918),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_775),
.B(n_372),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_868),
.A2(n_920),
.B(n_919),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_781),
.A2(n_496),
.B1(n_493),
.B2(n_483),
.Y(n_1026)
);

BUFx4f_ASAP7_75t_L g1027 ( 
.A(n_830),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_840),
.A2(n_922),
.B(n_774),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_837),
.B(n_493),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_779),
.B(n_372),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_846),
.B(n_372),
.Y(n_1031)
);

O2A1O1Ixp5_ASAP7_75t_SL g1032 ( 
.A1(n_797),
.A2(n_9),
.B(n_11),
.C(n_13),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_829),
.A2(n_9),
.B(n_14),
.C(n_16),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_846),
.B(n_14),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_768),
.A2(n_206),
.B(n_199),
.Y(n_1035)
);

AOI21x1_ASAP7_75t_L g1036 ( 
.A1(n_860),
.A2(n_190),
.B(n_180),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_823),
.B(n_16),
.Y(n_1037)
);

NOR3xp33_ASAP7_75t_L g1038 ( 
.A(n_788),
.B(n_17),
.C(n_18),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_802),
.A2(n_170),
.B(n_157),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_897),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_854),
.A2(n_155),
.B(n_153),
.Y(n_1041)
);

BUFx8_ASAP7_75t_L g1042 ( 
.A(n_904),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_856),
.A2(n_150),
.B(n_146),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_790),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_858),
.A2(n_862),
.B(n_889),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_832),
.B(n_17),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_765),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_801),
.B(n_19),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_834),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_801),
.B(n_22),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_799),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_925),
.B(n_23),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_855),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_866),
.A2(n_144),
.B1(n_108),
.B2(n_101),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_839),
.A2(n_93),
.B(n_26),
.Y(n_1055)
);

INVxp67_ASAP7_75t_L g1056 ( 
.A(n_901),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_923),
.A2(n_24),
.B(n_27),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_L g1058 ( 
.A(n_773),
.B(n_872),
.C(n_761),
.Y(n_1058)
);

NAND2x1_ASAP7_75t_L g1059 ( 
.A(n_897),
.B(n_24),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_855),
.A2(n_28),
.B(n_35),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_890),
.A2(n_28),
.B(n_36),
.C(n_37),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_872),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_857),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_SL g1064 ( 
.A1(n_898),
.A2(n_38),
.B(n_40),
.C(n_42),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_873),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_857),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_898),
.A2(n_40),
.B(n_42),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_804),
.B(n_44),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_899),
.B(n_46),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_818),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_818),
.B(n_47),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_761),
.B(n_74),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_818),
.B(n_47),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_SL g1074 ( 
.A(n_838),
.B(n_48),
.C(n_49),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_803),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_891),
.B(n_52),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_789),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1077)
);

NAND3xp33_ASAP7_75t_L g1078 ( 
.A(n_911),
.B(n_54),
.C(n_56),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_897),
.Y(n_1079)
);

BUFx8_ASAP7_75t_L g1080 ( 
.A(n_873),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_805),
.B(n_848),
.Y(n_1081)
);

AOI21xp33_ASAP7_75t_L g1082 ( 
.A1(n_842),
.A2(n_816),
.B(n_778),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_873),
.Y(n_1083)
);

AOI21x1_ASAP7_75t_L g1084 ( 
.A1(n_908),
.A2(n_56),
.B(n_63),
.Y(n_1084)
);

CKINVDCx10_ASAP7_75t_R g1085 ( 
.A(n_777),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_806),
.B(n_64),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_809),
.B(n_66),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_816),
.A2(n_73),
.B(n_68),
.C(n_69),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_812),
.A2(n_67),
.B1(n_72),
.B2(n_813),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_869),
.A2(n_67),
.B(n_72),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_887),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_821),
.B(n_828),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_822),
.B(n_843),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_900),
.A2(n_909),
.B(n_910),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_871),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_825),
.B(n_827),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_842),
.A2(n_917),
.B1(n_888),
.B2(n_905),
.Y(n_1097)
);

NAND2x1p5_ASAP7_75t_L g1098 ( 
.A(n_871),
.B(n_888),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_783),
.A2(n_784),
.B(n_800),
.Y(n_1099)
);

AOI21x1_ASAP7_75t_L g1100 ( 
.A1(n_900),
.A2(n_910),
.B(n_909),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_787),
.B(n_903),
.C(n_907),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_880),
.A2(n_884),
.B(n_913),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_880),
.A2(n_884),
.B(n_913),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_897),
.Y(n_1104)
);

AOI21x1_ASAP7_75t_L g1105 ( 
.A1(n_783),
.A2(n_784),
.B(n_800),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_887),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_964),
.B(n_895),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_977),
.A2(n_887),
.B(n_831),
.C(n_877),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_993),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1105),
.A2(n_935),
.B(n_934),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1056),
.A2(n_831),
.B1(n_876),
.B2(n_877),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_966),
.A2(n_876),
.B(n_879),
.Y(n_1112)
);

AOI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_1048),
.A2(n_916),
.B(n_879),
.Y(n_1113)
);

INVx5_ASAP7_75t_L g1114 ( 
.A(n_1040),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_942),
.B(n_1044),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_929),
.A2(n_893),
.B(n_931),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1049),
.Y(n_1117)
);

XNOR2xp5_ASAP7_75t_L g1118 ( 
.A(n_994),
.B(n_893),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1045),
.A2(n_998),
.B(n_957),
.Y(n_1119)
);

BUFx5_ASAP7_75t_L g1120 ( 
.A(n_1053),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_932),
.A2(n_1023),
.B(n_936),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_952),
.A2(n_1050),
.B(n_1082),
.C(n_930),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_933),
.B(n_1058),
.Y(n_1123)
);

AO31x2_ASAP7_75t_L g1124 ( 
.A1(n_1013),
.A2(n_981),
.A3(n_1002),
.B(n_1097),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_966),
.A2(n_1025),
.B(n_943),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1075),
.B(n_953),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_955),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_956),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1096),
.A2(n_1003),
.B1(n_968),
.B2(n_944),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1045),
.A2(n_1025),
.B(n_1101),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_940),
.B(n_988),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1077),
.A2(n_1062),
.B(n_1071),
.C(n_1035),
.Y(n_1132)
);

O2A1O1Ixp5_ASAP7_75t_L g1133 ( 
.A1(n_1028),
.A2(n_1023),
.B(n_1093),
.C(n_1081),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_959),
.B(n_946),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_943),
.A2(n_945),
.B(n_1102),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_932),
.A2(n_936),
.B(n_985),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1094),
.A2(n_978),
.B(n_1102),
.Y(n_1137)
);

AND2x2_ASAP7_75t_SL g1138 ( 
.A(n_1038),
.B(n_963),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_970),
.A2(n_1092),
.B(n_965),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1063),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_945),
.A2(n_1103),
.B(n_974),
.Y(n_1141)
);

BUFx12f_ASAP7_75t_L g1142 ( 
.A(n_1080),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1103),
.A2(n_974),
.B(n_972),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_960),
.B(n_982),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_967),
.B(n_969),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_975),
.B(n_979),
.Y(n_1146)
);

INVxp67_ASAP7_75t_SL g1147 ( 
.A(n_939),
.Y(n_1147)
);

AO21x1_ASAP7_75t_L g1148 ( 
.A1(n_983),
.A2(n_1069),
.B(n_1041),
.Y(n_1148)
);

AND3x4_ASAP7_75t_L g1149 ( 
.A(n_1007),
.B(n_990),
.C(n_1091),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1016),
.B(n_1018),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1076),
.B(n_1029),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1094),
.A2(n_965),
.B(n_1017),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1037),
.B(n_1046),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_972),
.A2(n_976),
.B(n_1099),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1040),
.B(n_1079),
.Y(n_1155)
);

NOR2x1_ASAP7_75t_SL g1156 ( 
.A(n_1040),
.B(n_1079),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1079),
.Y(n_1157)
);

AO21x2_ASAP7_75t_L g1158 ( 
.A1(n_991),
.A2(n_1017),
.B(n_1001),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1051),
.B(n_1072),
.Y(n_1159)
);

NAND2x1_ASAP7_75t_L g1160 ( 
.A(n_971),
.B(n_973),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1066),
.Y(n_1161)
);

AOI21x1_ASAP7_75t_L g1162 ( 
.A1(n_976),
.A2(n_951),
.B(n_947),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1086),
.B(n_1087),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1104),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1100),
.A2(n_962),
.B(n_954),
.Y(n_1165)
);

CKINVDCx6p67_ASAP7_75t_R g1166 ( 
.A(n_1083),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_950),
.A2(n_999),
.B(n_992),
.Y(n_1167)
);

INVx5_ASAP7_75t_L g1168 ( 
.A(n_1104),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1015),
.A2(n_1021),
.B(n_984),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1008),
.A2(n_1011),
.B(n_941),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_949),
.B(n_1004),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1022),
.A2(n_1010),
.B(n_1012),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_1052),
.Y(n_1173)
);

AO22x1_ASAP7_75t_L g1174 ( 
.A1(n_1073),
.A2(n_1042),
.B1(n_1070),
.B2(n_1080),
.Y(n_1174)
);

NAND2xp33_ASAP7_75t_L g1175 ( 
.A(n_939),
.B(n_995),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1095),
.Y(n_1176)
);

NAND2x1p5_ASAP7_75t_L g1177 ( 
.A(n_973),
.B(n_1104),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_997),
.A2(n_1098),
.B(n_987),
.Y(n_1178)
);

AND2x6_ASAP7_75t_L g1179 ( 
.A(n_971),
.B(n_995),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1020),
.A2(n_1009),
.B(n_1078),
.C(n_1089),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_1042),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_939),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1034),
.B(n_989),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_961),
.Y(n_1184)
);

AOI21x1_ASAP7_75t_SL g1185 ( 
.A1(n_1031),
.A2(n_1032),
.B(n_1036),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1047),
.A2(n_1088),
.B(n_1033),
.C(n_1061),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1060),
.A2(n_1090),
.A3(n_1057),
.B(n_1039),
.Y(n_1187)
);

AOI21xp33_ASAP7_75t_L g1188 ( 
.A1(n_980),
.A2(n_1005),
.B(n_1024),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_996),
.B(n_995),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_986),
.A2(n_948),
.B(n_958),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1039),
.A2(n_1067),
.A3(n_1043),
.B(n_1041),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1043),
.A2(n_1030),
.B(n_1059),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_937),
.B(n_1014),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1055),
.A2(n_1084),
.B(n_1067),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_961),
.Y(n_1195)
);

OA21x2_ASAP7_75t_L g1196 ( 
.A1(n_1068),
.A2(n_1054),
.B(n_1026),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_961),
.A2(n_1064),
.B(n_1006),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1019),
.A2(n_1074),
.B(n_1106),
.Y(n_1198)
);

BUFx12f_ASAP7_75t_L g1199 ( 
.A(n_938),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1000),
.A2(n_1027),
.B(n_1065),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1000),
.A2(n_977),
.A3(n_957),
.B(n_1013),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1027),
.B(n_1085),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_964),
.B(n_942),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1105),
.A2(n_935),
.B(n_934),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_964),
.B(n_942),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_964),
.B(n_933),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_977),
.A2(n_929),
.B(n_931),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_964),
.B(n_942),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1105),
.A2(n_935),
.B(n_934),
.Y(n_1209)
);

AND2x2_ASAP7_75t_SL g1210 ( 
.A(n_1048),
.B(n_1050),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_1080),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_964),
.B(n_942),
.Y(n_1212)
);

NAND3xp33_ASAP7_75t_L g1213 ( 
.A(n_977),
.B(n_1048),
.C(n_882),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1105),
.A2(n_935),
.B(n_934),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_964),
.B(n_933),
.Y(n_1215)
);

NOR2xp67_ASAP7_75t_L g1216 ( 
.A(n_1056),
.B(n_914),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_977),
.A2(n_929),
.B(n_931),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_964),
.B(n_942),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_993),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1105),
.A2(n_935),
.B(n_934),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1080),
.Y(n_1221)
);

NAND3xp33_ASAP7_75t_L g1222 ( 
.A(n_977),
.B(n_1048),
.C(n_882),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_977),
.A2(n_861),
.B(n_824),
.Y(n_1223)
);

NAND2x1_ASAP7_75t_L g1224 ( 
.A(n_971),
.B(n_861),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_977),
.A2(n_861),
.B(n_824),
.Y(n_1225)
);

BUFx8_ASAP7_75t_L g1226 ( 
.A(n_1083),
.Y(n_1226)
);

AO21x2_ASAP7_75t_L g1227 ( 
.A1(n_977),
.A2(n_957),
.B(n_981),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1048),
.A2(n_786),
.B1(n_1074),
.B2(n_1050),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1105),
.A2(n_935),
.B(n_934),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_977),
.A2(n_957),
.A3(n_1013),
.B(n_981),
.Y(n_1230)
);

AND3x1_ASAP7_75t_SL g1231 ( 
.A(n_1049),
.B(n_882),
.C(n_698),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_977),
.A2(n_957),
.A3(n_1013),
.B(n_981),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1016),
.B(n_1018),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_977),
.A2(n_929),
.B(n_931),
.Y(n_1234)
);

OR2x6_ASAP7_75t_L g1235 ( 
.A(n_1083),
.B(n_830),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_977),
.A2(n_1056),
.B1(n_1044),
.B2(n_930),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1040),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_977),
.A2(n_929),
.B(n_931),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1044),
.B(n_1056),
.Y(n_1239)
);

CKINVDCx8_ASAP7_75t_R g1240 ( 
.A(n_1083),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_993),
.Y(n_1241)
);

BUFx8_ASAP7_75t_SL g1242 ( 
.A(n_994),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_SL g1243 ( 
.A1(n_977),
.A2(n_861),
.B(n_772),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_977),
.A2(n_929),
.B(n_931),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1243),
.A2(n_1225),
.B(n_1223),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1203),
.B(n_1205),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1233),
.B(n_1156),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1206),
.B(n_1215),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1144),
.B(n_1171),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1114),
.B(n_1168),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1208),
.B(n_1212),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1150),
.Y(n_1252)
);

OAI21xp33_ASAP7_75t_L g1253 ( 
.A1(n_1171),
.A2(n_1144),
.B(n_1115),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1131),
.B(n_1233),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1218),
.B(n_1151),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1138),
.A2(n_1210),
.B1(n_1193),
.B2(n_1236),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1138),
.B(n_1210),
.Y(n_1257)
);

INVx8_ASAP7_75t_L g1258 ( 
.A(n_1179),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1239),
.B(n_1126),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1114),
.B(n_1168),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1120),
.Y(n_1261)
);

OR2x6_ASAP7_75t_L g1262 ( 
.A(n_1235),
.B(n_1174),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1122),
.A2(n_1228),
.B(n_1132),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1239),
.B(n_1123),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1242),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1120),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1173),
.B(n_1159),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1147),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1114),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1228),
.A2(n_1132),
.B(n_1129),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1134),
.A2(n_1123),
.B1(n_1244),
.B2(n_1207),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1117),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1226),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_1118),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1140),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1114),
.B(n_1168),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_SL g1277 ( 
.A1(n_1180),
.A2(n_1186),
.B(n_1134),
.C(n_1108),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1161),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1217),
.A2(n_1238),
.B(n_1234),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1226),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1153),
.B(n_1188),
.Y(n_1281)
);

OR2x6_ASAP7_75t_L g1282 ( 
.A(n_1235),
.B(n_1199),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1163),
.B(n_1216),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1109),
.B(n_1219),
.Y(n_1284)
);

OAI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1241),
.A2(n_1107),
.B1(n_1146),
.B2(n_1145),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1196),
.A2(n_1148),
.B1(n_1149),
.B2(n_1227),
.Y(n_1286)
);

AO21x1_ASAP7_75t_L g1287 ( 
.A1(n_1190),
.A2(n_1192),
.B(n_1178),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1166),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1181),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1183),
.B(n_1176),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1127),
.B(n_1128),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1157),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1235),
.B(n_1200),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1195),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1157),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1157),
.Y(n_1296)
);

NAND2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1184),
.B(n_1157),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1221),
.Y(n_1298)
);

INVx3_ASAP7_75t_SL g1299 ( 
.A(n_1211),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1130),
.B(n_1120),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1113),
.A2(n_1133),
.B(n_1197),
.C(n_1111),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1184),
.B(n_1182),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1202),
.B(n_1182),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1149),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1189),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1175),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1164),
.B(n_1237),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1164),
.B(n_1237),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1201),
.B(n_1198),
.Y(n_1309)
);

O2A1O1Ixp5_ASAP7_75t_SL g1310 ( 
.A1(n_1119),
.A2(n_1152),
.B(n_1116),
.C(n_1137),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1155),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1164),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1240),
.B(n_1201),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1164),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1196),
.A2(n_1227),
.B1(n_1197),
.B2(n_1231),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1139),
.B(n_1201),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1237),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1136),
.A2(n_1192),
.B(n_1178),
.C(n_1121),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1201),
.B(n_1155),
.Y(n_1319)
);

BUFx4_ASAP7_75t_SL g1320 ( 
.A(n_1142),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1231),
.A2(n_1158),
.B1(n_1194),
.B2(n_1170),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1237),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1124),
.B(n_1232),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1143),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1124),
.B(n_1232),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1177),
.B(n_1232),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1177),
.B(n_1232),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1124),
.B(n_1230),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1162),
.B(n_1160),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1179),
.A2(n_1170),
.B1(n_1158),
.B2(n_1224),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1124),
.B(n_1230),
.Y(n_1331)
);

CKINVDCx8_ASAP7_75t_R g1332 ( 
.A(n_1179),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1167),
.A2(n_1172),
.B(n_1165),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1179),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1172),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1191),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1187),
.Y(n_1337)
);

OAI21xp33_ASAP7_75t_L g1338 ( 
.A1(n_1125),
.A2(n_1154),
.B(n_1112),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1187),
.B(n_1230),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1135),
.A2(n_1141),
.B(n_1110),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1191),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1230),
.B(n_1191),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1204),
.Y(n_1343)
);

INVx4_ASAP7_75t_L g1344 ( 
.A(n_1185),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1209),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1169),
.A2(n_1214),
.B1(n_1220),
.B2(n_1229),
.Y(n_1346)
);

BUFx12f_ASAP7_75t_L g1347 ( 
.A(n_1185),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1233),
.B(n_1156),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1120),
.Y(n_1349)
);

INVx3_ASAP7_75t_SL g1350 ( 
.A(n_1166),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1117),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1120),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1203),
.B(n_1205),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1233),
.Y(n_1354)
);

NAND2x1p5_ASAP7_75t_L g1355 ( 
.A(n_1114),
.B(n_1168),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1203),
.B(n_1205),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1144),
.B(n_1171),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1114),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1144),
.B(n_1171),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1206),
.B(n_1215),
.Y(n_1360)
);

INVx5_ASAP7_75t_L g1361 ( 
.A(n_1179),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1150),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1150),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1213),
.A2(n_977),
.B(n_1222),
.C(n_1048),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1206),
.B(n_1215),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1242),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1233),
.B(n_1016),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1203),
.B(n_1205),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1120),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1203),
.B(n_1205),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1242),
.Y(n_1371)
);

INVx4_ASAP7_75t_L g1372 ( 
.A(n_1114),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1203),
.B(n_1205),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1233),
.B(n_1016),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1203),
.B(n_1205),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_R g1376 ( 
.A(n_1240),
.B(n_659),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1242),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1117),
.Y(n_1378)
);

BUFx4f_ASAP7_75t_L g1379 ( 
.A(n_1199),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1114),
.Y(n_1380)
);

BUFx12f_ASAP7_75t_L g1381 ( 
.A(n_1142),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1206),
.B(n_1215),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1242),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1203),
.B(n_1205),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1206),
.B(n_1215),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1203),
.B(n_1205),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1272),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1357),
.B(n_1359),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1340),
.A2(n_1245),
.B(n_1333),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1351),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1378),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1357),
.A2(n_1359),
.B1(n_1264),
.B2(n_1256),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1275),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1278),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1270),
.A2(n_1263),
.B1(n_1281),
.B2(n_1249),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1284),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1281),
.A2(n_1264),
.B1(n_1253),
.B2(n_1283),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1291),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1283),
.A2(n_1257),
.B1(n_1304),
.B2(n_1255),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1246),
.A2(n_1386),
.B1(n_1353),
.B2(n_1356),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1318),
.A2(n_1338),
.B(n_1286),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1305),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1290),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1254),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1271),
.A2(n_1279),
.B1(n_1373),
.B2(n_1384),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1268),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1268),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1335),
.A2(n_1376),
.B1(n_1259),
.B2(n_1370),
.Y(n_1408)
);

CKINVDCx11_ASAP7_75t_R g1409 ( 
.A(n_1381),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1252),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1335),
.A2(n_1376),
.B1(n_1375),
.B2(n_1251),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1354),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1362),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1367),
.Y(n_1414)
);

BUFx4f_ASAP7_75t_SL g1415 ( 
.A(n_1381),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1363),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1248),
.B(n_1360),
.Y(n_1417)
);

AND2x6_ASAP7_75t_L g1418 ( 
.A(n_1261),
.B(n_1266),
.Y(n_1418)
);

AO21x1_ASAP7_75t_L g1419 ( 
.A1(n_1285),
.A2(n_1344),
.B(n_1301),
.Y(n_1419)
);

INVx4_ASAP7_75t_L g1420 ( 
.A(n_1260),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1363),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1311),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1311),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1294),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1368),
.A2(n_1279),
.B1(n_1313),
.B2(n_1267),
.Y(n_1425)
);

BUFx12f_ASAP7_75t_L g1426 ( 
.A(n_1265),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1365),
.Y(n_1427)
);

INVx4_ASAP7_75t_SL g1428 ( 
.A(n_1260),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1382),
.B(n_1385),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1306),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1247),
.B(n_1348),
.Y(n_1431)
);

CKINVDCx6p67_ASAP7_75t_R g1432 ( 
.A(n_1371),
.Y(n_1432)
);

AO21x1_ASAP7_75t_SL g1433 ( 
.A1(n_1286),
.A2(n_1315),
.B(n_1271),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1279),
.A2(n_1262),
.B1(n_1274),
.B2(n_1273),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1367),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1318),
.A2(n_1277),
.B(n_1364),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1287),
.A2(n_1346),
.B(n_1330),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1374),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1314),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1364),
.A2(n_1303),
.B1(n_1374),
.B2(n_1247),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1265),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1262),
.A2(n_1273),
.B1(n_1280),
.B2(n_1379),
.Y(n_1442)
);

OAI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1262),
.A2(n_1299),
.B1(n_1282),
.B2(n_1350),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1247),
.Y(n_1444)
);

AOI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1316),
.A2(n_1300),
.B(n_1324),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1322),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1348),
.B(n_1285),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1315),
.A2(n_1339),
.B1(n_1347),
.B2(n_1321),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1293),
.A2(n_1282),
.B1(n_1298),
.B2(n_1379),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1293),
.A2(n_1347),
.B1(n_1282),
.B2(n_1361),
.Y(n_1450)
);

NAND2x1p5_ASAP7_75t_L g1451 ( 
.A(n_1361),
.B(n_1276),
.Y(n_1451)
);

INVx11_ASAP7_75t_L g1452 ( 
.A(n_1320),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1350),
.Y(n_1453)
);

CKINVDCx11_ASAP7_75t_R g1454 ( 
.A(n_1299),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1292),
.Y(n_1455)
);

OAI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1288),
.A2(n_1289),
.B1(n_1332),
.B2(n_1361),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1349),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1292),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1366),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1260),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1366),
.Y(n_1461)
);

OR2x6_ASAP7_75t_L g1462 ( 
.A(n_1336),
.B(n_1341),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1361),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1276),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1352),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1276),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1295),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1295),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1352),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1258),
.Y(n_1470)
);

CKINVDCx11_ASAP7_75t_R g1471 ( 
.A(n_1371),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1342),
.B(n_1327),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1296),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1369),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1339),
.A2(n_1321),
.B1(n_1341),
.B2(n_1336),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1369),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1339),
.A2(n_1344),
.B1(n_1337),
.B2(n_1323),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1377),
.A2(n_1383),
.B1(n_1258),
.B2(n_1309),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1302),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1277),
.B(n_1310),
.Y(n_1480)
);

CKINVDCx11_ASAP7_75t_R g1481 ( 
.A(n_1320),
.Y(n_1481)
);

NAND2x1p5_ASAP7_75t_L g1482 ( 
.A(n_1372),
.B(n_1380),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1302),
.B(n_1307),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1308),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1296),
.Y(n_1485)
);

INVx6_ASAP7_75t_L g1486 ( 
.A(n_1258),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1319),
.Y(n_1487)
);

BUFx2_ASAP7_75t_R g1488 ( 
.A(n_1269),
.Y(n_1488)
);

CKINVDCx16_ASAP7_75t_R g1489 ( 
.A(n_1307),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1308),
.B(n_1317),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1337),
.A2(n_1331),
.B1(n_1328),
.B2(n_1325),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1345),
.A2(n_1326),
.B(n_1329),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1334),
.B(n_1380),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1312),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1343),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1312),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1250),
.A2(n_1355),
.B1(n_1297),
.B2(n_1372),
.Y(n_1497)
);

INVx8_ASAP7_75t_L g1498 ( 
.A(n_1312),
.Y(n_1498)
);

CKINVDCx11_ASAP7_75t_R g1499 ( 
.A(n_1343),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1297),
.Y(n_1500)
);

NOR2x1_ASAP7_75t_R g1501 ( 
.A(n_1358),
.B(n_1343),
.Y(n_1501)
);

CKINVDCx6p67_ASAP7_75t_R g1502 ( 
.A(n_1343),
.Y(n_1502)
);

BUFx2_ASAP7_75t_R g1503 ( 
.A(n_1250),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1260),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1258),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1357),
.B(n_1359),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1357),
.A2(n_1359),
.B1(n_1171),
.B2(n_977),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1357),
.B(n_1359),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1260),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1357),
.A2(n_1359),
.B1(n_1144),
.B2(n_720),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1272),
.Y(n_1511)
);

CKINVDCx11_ASAP7_75t_R g1512 ( 
.A(n_1381),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1354),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1272),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1267),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1354),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1248),
.B(n_1360),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1247),
.B(n_1348),
.Y(n_1518)
);

BUFx12f_ASAP7_75t_L g1519 ( 
.A(n_1381),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1354),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1361),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1361),
.Y(n_1522)
);

NAND2x1p5_ASAP7_75t_L g1523 ( 
.A(n_1361),
.B(n_1260),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1254),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1436),
.A2(n_1507),
.B(n_1400),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1472),
.B(n_1487),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1392),
.A2(n_1510),
.B1(n_1395),
.B2(n_1411),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1417),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1517),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1506),
.B(n_1388),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1397),
.B(n_1506),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1472),
.B(n_1395),
.Y(n_1532)
);

OA21x2_ASAP7_75t_L g1533 ( 
.A1(n_1480),
.A2(n_1419),
.B(n_1389),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1445),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1462),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1508),
.B(n_1403),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1462),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1410),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1425),
.B(n_1433),
.Y(n_1539)
);

INVxp33_ASAP7_75t_L g1540 ( 
.A(n_1429),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1462),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1492),
.Y(n_1542)
);

OA21x2_ASAP7_75t_L g1543 ( 
.A1(n_1491),
.A2(n_1475),
.B(n_1448),
.Y(n_1543)
);

OA21x2_ASAP7_75t_L g1544 ( 
.A1(n_1491),
.A2(n_1475),
.B(n_1448),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1405),
.B(n_1422),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_SL g1546 ( 
.A1(n_1501),
.A2(n_1523),
.B(n_1451),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1492),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1515),
.B(n_1404),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1405),
.B(n_1423),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1492),
.B(n_1413),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1408),
.A2(n_1399),
.B(n_1447),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1418),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1401),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1524),
.B(n_1402),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1401),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1416),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_SL g1557 ( 
.A(n_1437),
.B(n_1430),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1401),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1398),
.B(n_1427),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1457),
.B(n_1465),
.Y(n_1560)
);

OR2x6_ASAP7_75t_L g1561 ( 
.A(n_1447),
.B(n_1495),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1469),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1396),
.B(n_1421),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1474),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1476),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1406),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1418),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1463),
.A2(n_1522),
.B(n_1521),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1476),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1414),
.B(n_1435),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1418),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1407),
.B(n_1477),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1418),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1418),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1502),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1502),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1477),
.B(n_1431),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_SL g1578 ( 
.A(n_1488),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1387),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1390),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1391),
.Y(n_1581)
);

AO21x1_ASAP7_75t_L g1582 ( 
.A1(n_1478),
.A2(n_1393),
.B(n_1394),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1438),
.B(n_1424),
.Y(n_1583)
);

BUFx2_ASAP7_75t_R g1584 ( 
.A(n_1459),
.Y(n_1584)
);

AND2x2_ASAP7_75t_SL g1585 ( 
.A(n_1440),
.B(n_1489),
.Y(n_1585)
);

AO21x1_ASAP7_75t_SL g1586 ( 
.A1(n_1449),
.A2(n_1514),
.B(n_1511),
.Y(n_1586)
);

AO31x2_ASAP7_75t_L g1587 ( 
.A1(n_1455),
.A2(n_1485),
.A3(n_1467),
.B(n_1473),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1431),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1493),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1493),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1493),
.Y(n_1591)
);

OA21x2_ASAP7_75t_L g1592 ( 
.A1(n_1458),
.A2(n_1468),
.B(n_1494),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1412),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1496),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1499),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1463),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1521),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1513),
.B(n_1516),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1522),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1499),
.Y(n_1600)
);

AO21x2_ASAP7_75t_L g1601 ( 
.A1(n_1443),
.A2(n_1456),
.B(n_1497),
.Y(n_1601)
);

AOI21x1_ASAP7_75t_L g1602 ( 
.A1(n_1500),
.A2(n_1518),
.B(n_1446),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1490),
.B(n_1444),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1470),
.B(n_1428),
.Y(n_1604)
);

AO21x1_ASAP7_75t_SL g1605 ( 
.A1(n_1439),
.A2(n_1434),
.B(n_1450),
.Y(n_1605)
);

OA21x2_ASAP7_75t_L g1606 ( 
.A1(n_1484),
.A2(n_1505),
.B(n_1479),
.Y(n_1606)
);

AOI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1442),
.A2(n_1454),
.B1(n_1519),
.B2(n_1453),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1498),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1486),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1516),
.B(n_1520),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1520),
.Y(n_1611)
);

AOI21xp33_ASAP7_75t_L g1612 ( 
.A1(n_1505),
.A2(n_1464),
.B(n_1509),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1464),
.B(n_1523),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1454),
.A2(n_1519),
.B1(n_1432),
.B2(n_1415),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1526),
.B(n_1483),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1535),
.B(n_1470),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1606),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1532),
.B(n_1460),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1559),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1606),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1550),
.B(n_1432),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1592),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1577),
.B(n_1460),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1592),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1536),
.B(n_1466),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1606),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1530),
.B(n_1466),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1592),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1592),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1554),
.B(n_1531),
.Y(n_1630)
);

NOR4xp25_ASAP7_75t_SL g1631 ( 
.A(n_1575),
.B(n_1461),
.C(n_1459),
.D(n_1503),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1550),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1579),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1579),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1546),
.B(n_1486),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1606),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1580),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1555),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1561),
.B(n_1466),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1535),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1547),
.B(n_1482),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1580),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1537),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1525),
.B(n_1504),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1581),
.Y(n_1645)
);

NOR2x1_ASAP7_75t_SL g1646 ( 
.A(n_1605),
.B(n_1504),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1527),
.A2(n_1409),
.B1(n_1512),
.B2(n_1471),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1598),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1561),
.B(n_1545),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1548),
.B(n_1420),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1538),
.B(n_1420),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1545),
.B(n_1471),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1556),
.Y(n_1653)
);

NOR2x1_ASAP7_75t_L g1654 ( 
.A(n_1601),
.B(n_1441),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1549),
.B(n_1498),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1587),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1566),
.B(n_1498),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1549),
.B(n_1461),
.Y(n_1658)
);

OAI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1551),
.A2(n_1415),
.B1(n_1426),
.B2(n_1441),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1587),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1583),
.B(n_1540),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1541),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1575),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1541),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1587),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1528),
.B(n_1426),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_1600),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1547),
.B(n_1409),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1542),
.B(n_1512),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1543),
.B(n_1481),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1543),
.B(n_1481),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1590),
.B(n_1452),
.Y(n_1672)
);

AND2x4_ASAP7_75t_SL g1673 ( 
.A(n_1567),
.B(n_1600),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1529),
.B(n_1563),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1590),
.B(n_1573),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1593),
.B(n_1611),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1649),
.B(n_1539),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1648),
.B(n_1539),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1630),
.B(n_1572),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1647),
.A2(n_1607),
.B(n_1614),
.Y(n_1680)
);

AND2x2_ASAP7_75t_SL g1681 ( 
.A(n_1670),
.B(n_1585),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1654),
.B(n_1582),
.Y(n_1682)
);

OA21x2_ASAP7_75t_L g1683 ( 
.A1(n_1622),
.A2(n_1553),
.B(n_1558),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1619),
.B(n_1572),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1649),
.B(n_1542),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1654),
.B(n_1607),
.C(n_1591),
.Y(n_1686)
);

OAI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1668),
.A2(n_1614),
.B1(n_1610),
.B2(n_1570),
.C(n_1595),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_SL g1688 ( 
.A1(n_1659),
.A2(n_1600),
.B(n_1604),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_SL g1689 ( 
.A(n_1635),
.B(n_1584),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1661),
.B(n_1589),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1674),
.A2(n_1582),
.B1(n_1676),
.B2(n_1670),
.C(n_1671),
.Y(n_1691)
);

OA21x2_ASAP7_75t_L g1692 ( 
.A1(n_1622),
.A2(n_1628),
.B(n_1624),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1625),
.B(n_1591),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1631),
.A2(n_1578),
.B1(n_1585),
.B2(n_1595),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_SL g1695 ( 
.A1(n_1671),
.A2(n_1585),
.B1(n_1543),
.B2(n_1544),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1650),
.B(n_1587),
.Y(n_1696)
);

AND2x2_ASAP7_75t_SL g1697 ( 
.A(n_1668),
.B(n_1543),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1666),
.A2(n_1644),
.B1(n_1669),
.B2(n_1652),
.C(n_1627),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1632),
.B(n_1544),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1632),
.B(n_1544),
.Y(n_1700)
);

NAND4xp25_ASAP7_75t_L g1701 ( 
.A(n_1652),
.B(n_1595),
.C(n_1594),
.D(n_1534),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1621),
.B(n_1552),
.Y(n_1702)
);

AOI211xp5_ASAP7_75t_L g1703 ( 
.A1(n_1658),
.A2(n_1546),
.B(n_1600),
.C(n_1612),
.Y(n_1703)
);

NAND3xp33_ASAP7_75t_L g1704 ( 
.A(n_1669),
.B(n_1596),
.C(n_1597),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1621),
.B(n_1587),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_L g1706 ( 
.A(n_1656),
.B(n_1665),
.C(n_1641),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1658),
.A2(n_1600),
.B(n_1604),
.Y(n_1707)
);

OAI21xp33_ASAP7_75t_L g1708 ( 
.A1(n_1617),
.A2(n_1602),
.B(n_1594),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_L g1709 ( 
.A(n_1641),
.B(n_1597),
.C(n_1596),
.Y(n_1709)
);

NAND3xp33_ASAP7_75t_L g1710 ( 
.A(n_1651),
.B(n_1626),
.C(n_1620),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1618),
.B(n_1534),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1618),
.B(n_1601),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1623),
.B(n_1601),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1640),
.B(n_1643),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1623),
.B(n_1560),
.Y(n_1715)
);

NAND3xp33_ASAP7_75t_L g1716 ( 
.A(n_1636),
.B(n_1599),
.C(n_1533),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1640),
.B(n_1557),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1672),
.B(n_1600),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1667),
.A2(n_1552),
.B1(n_1571),
.B2(n_1588),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1662),
.B(n_1533),
.Y(n_1720)
);

OAI21xp33_ASAP7_75t_L g1721 ( 
.A1(n_1615),
.A2(n_1602),
.B(n_1603),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1664),
.B(n_1533),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1653),
.B(n_1562),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1664),
.B(n_1533),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1672),
.A2(n_1605),
.B1(n_1586),
.B2(n_1588),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1657),
.A2(n_1568),
.B(n_1613),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1633),
.B(n_1564),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1633),
.B(n_1565),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1675),
.B(n_1553),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1634),
.B(n_1565),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1634),
.B(n_1569),
.Y(n_1731)
);

OAI221xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1635),
.A2(n_1613),
.B1(n_1571),
.B2(n_1574),
.C(n_1573),
.Y(n_1732)
);

NAND2xp33_ASAP7_75t_SL g1733 ( 
.A(n_1655),
.B(n_1576),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1692),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1685),
.B(n_1624),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1685),
.B(n_1628),
.Y(n_1736)
);

NAND2x1p5_ASAP7_75t_L g1737 ( 
.A(n_1682),
.B(n_1660),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1692),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1696),
.B(n_1629),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1692),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1717),
.B(n_1667),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1729),
.B(n_1629),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1679),
.B(n_1637),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1677),
.B(n_1697),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1683),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1683),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1683),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1705),
.B(n_1712),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1697),
.B(n_1675),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1684),
.B(n_1699),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1720),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1727),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1703),
.B(n_1672),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1720),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1728),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1714),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1722),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1713),
.B(n_1711),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1699),
.B(n_1637),
.Y(n_1759)
);

NOR2x1_ASAP7_75t_R g1760 ( 
.A(n_1682),
.B(n_1667),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1733),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1724),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1730),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1731),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1710),
.B(n_1700),
.Y(n_1765)
);

AND2x4_ASAP7_75t_SL g1766 ( 
.A(n_1725),
.B(n_1635),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1700),
.B(n_1642),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1723),
.Y(n_1768)
);

NAND2x1_ASAP7_75t_L g1769 ( 
.A(n_1717),
.B(n_1714),
.Y(n_1769)
);

AND2x4_ASAP7_75t_SL g1770 ( 
.A(n_1718),
.B(n_1635),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1721),
.B(n_1642),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1726),
.B(n_1639),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1721),
.B(n_1638),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1681),
.B(n_1639),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1709),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1762),
.B(n_1681),
.Y(n_1776)
);

INVx3_ASAP7_75t_L g1777 ( 
.A(n_1734),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1742),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1762),
.B(n_1702),
.Y(n_1779)
);

INVx2_ASAP7_75t_SL g1780 ( 
.A(n_1761),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1744),
.B(n_1678),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1761),
.B(n_1706),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1765),
.B(n_1715),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1765),
.B(n_1690),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1744),
.B(n_1702),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1775),
.B(n_1691),
.Y(n_1786)
);

NAND3xp33_ASAP7_75t_L g1787 ( 
.A(n_1775),
.B(n_1680),
.C(n_1686),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1742),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1734),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1741),
.B(n_1695),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1748),
.B(n_1708),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1742),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1751),
.B(n_1754),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1748),
.B(n_1716),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1771),
.B(n_1694),
.C(n_1703),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1768),
.B(n_1708),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1741),
.Y(n_1797)
);

NAND2x1p5_ASAP7_75t_L g1798 ( 
.A(n_1769),
.B(n_1567),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1734),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1735),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1735),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1769),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1768),
.B(n_1739),
.Y(n_1803)
);

OAI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1753),
.A2(n_1688),
.B1(n_1689),
.B2(n_1701),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1739),
.B(n_1693),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1735),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1741),
.B(n_1707),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1736),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1736),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1745),
.Y(n_1810)
);

NOR2x1_ASAP7_75t_L g1811 ( 
.A(n_1738),
.B(n_1704),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1751),
.B(n_1754),
.Y(n_1812)
);

NAND2xp67_ASAP7_75t_L g1813 ( 
.A(n_1766),
.B(n_1673),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1760),
.A2(n_1733),
.B(n_1646),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1741),
.B(n_1616),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1745),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1752),
.B(n_1645),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1746),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1749),
.B(n_1616),
.Y(n_1819)
);

INVxp67_ASAP7_75t_L g1820 ( 
.A(n_1787),
.Y(n_1820)
);

NOR2xp67_ASAP7_75t_SL g1821 ( 
.A(n_1787),
.B(n_1687),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1776),
.B(n_1772),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1802),
.B(n_1749),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1817),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1794),
.B(n_1758),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1776),
.B(n_1772),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1786),
.B(n_1752),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1817),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1776),
.B(n_1790),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1777),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1790),
.B(n_1807),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1777),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1777),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_SL g1834 ( 
.A(n_1804),
.B(n_1760),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1786),
.B(n_1755),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1780),
.Y(n_1836)
);

OR4x1_ASAP7_75t_L g1837 ( 
.A(n_1780),
.B(n_1732),
.C(n_1756),
.D(n_1764),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1807),
.B(n_1785),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1810),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1810),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1796),
.B(n_1791),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1796),
.B(n_1755),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1785),
.B(n_1774),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1797),
.B(n_1774),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1780),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1810),
.Y(n_1846)
);

O2A1O1Ixp5_ASAP7_75t_L g1847 ( 
.A1(n_1804),
.A2(n_1771),
.B(n_1743),
.C(n_1773),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1797),
.B(n_1756),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_1782),
.Y(n_1849)
);

INVxp67_ASAP7_75t_SL g1850 ( 
.A(n_1811),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1791),
.B(n_1763),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1816),
.Y(n_1852)
);

BUFx3_ASAP7_75t_L g1853 ( 
.A(n_1782),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1797),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1816),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1811),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1779),
.B(n_1756),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1779),
.B(n_1754),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1794),
.B(n_1783),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1803),
.B(n_1763),
.Y(n_1860)
);

NOR3xp33_ASAP7_75t_SL g1861 ( 
.A(n_1795),
.B(n_1698),
.C(n_1719),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1779),
.B(n_1757),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1803),
.B(n_1764),
.Y(n_1863)
);

INVxp67_ASAP7_75t_L g1864 ( 
.A(n_1795),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1783),
.B(n_1758),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1839),
.Y(n_1866)
);

INVx1_ASAP7_75t_SL g1867 ( 
.A(n_1849),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1864),
.B(n_1784),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1839),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1854),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1820),
.B(n_1781),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1853),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1854),
.Y(n_1873)
);

HB1xp67_ASAP7_75t_L g1874 ( 
.A(n_1836),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1859),
.B(n_1784),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1821),
.B(n_1781),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1840),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1829),
.B(n_1782),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_1821),
.Y(n_1879)
);

OAI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1834),
.A2(n_1814),
.B1(n_1802),
.B2(n_1798),
.C(n_1737),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1859),
.B(n_1805),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1829),
.B(n_1782),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1861),
.B(n_1805),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1825),
.B(n_1778),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1840),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1834),
.A2(n_1766),
.B1(n_1814),
.B2(n_1770),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1853),
.Y(n_1887)
);

NOR2x1_ASAP7_75t_L g1888 ( 
.A(n_1853),
.B(n_1802),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1843),
.B(n_1798),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1846),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1825),
.B(n_1778),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1843),
.B(n_1798),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1850),
.B(n_1802),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1827),
.B(n_1788),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1856),
.A2(n_1798),
.B1(n_1737),
.B2(n_1766),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1846),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1827),
.B(n_1835),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1852),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1836),
.B(n_1815),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1835),
.B(n_1773),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1841),
.B(n_1819),
.Y(n_1901)
);

AOI222xp33_ASAP7_75t_L g1902 ( 
.A1(n_1841),
.A2(n_1773),
.B1(n_1792),
.B2(n_1788),
.C1(n_1719),
.C2(n_1812),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1865),
.B(n_1792),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1830),
.Y(n_1904)
);

OAI221xp5_ASAP7_75t_L g1905 ( 
.A1(n_1879),
.A2(n_1847),
.B1(n_1849),
.B2(n_1831),
.C(n_1845),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1876),
.B(n_1831),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1883),
.B(n_1838),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1871),
.B(n_1838),
.Y(n_1908)
);

NAND2xp33_ASAP7_75t_SL g1909 ( 
.A(n_1878),
.B(n_1837),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1868),
.A2(n_1842),
.B(n_1851),
.Y(n_1910)
);

AOI32xp33_ASAP7_75t_L g1911 ( 
.A1(n_1878),
.A2(n_1882),
.A3(n_1867),
.B1(n_1880),
.B2(n_1886),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_SL g1912 ( 
.A1(n_1882),
.A2(n_1837),
.B1(n_1844),
.B2(n_1826),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1899),
.B(n_1844),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1874),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1901),
.A2(n_1737),
.B1(n_1822),
.B2(n_1826),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1866),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1899),
.B(n_1822),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1875),
.B(n_1865),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1899),
.B(n_1823),
.Y(n_1919)
);

AOI222xp33_ASAP7_75t_L g1920 ( 
.A1(n_1900),
.A2(n_1851),
.B1(n_1842),
.B2(n_1857),
.C1(n_1858),
.C2(n_1862),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1869),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1877),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1885),
.Y(n_1923)
);

INVx3_ASAP7_75t_L g1924 ( 
.A(n_1872),
.Y(n_1924)
);

OAI22xp33_ASAP7_75t_SL g1925 ( 
.A1(n_1872),
.A2(n_1887),
.B1(n_1888),
.B2(n_1875),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1889),
.B(n_1823),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1890),
.Y(n_1927)
);

BUFx2_ASAP7_75t_L g1928 ( 
.A(n_1872),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1902),
.B(n_1823),
.Y(n_1929)
);

OAI21xp33_ASAP7_75t_L g1930 ( 
.A1(n_1897),
.A2(n_1828),
.B(n_1824),
.Y(n_1930)
);

INVx1_ASAP7_75t_SL g1931 ( 
.A(n_1887),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1897),
.B(n_1860),
.Y(n_1932)
);

OAI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1887),
.A2(n_1737),
.B1(n_1635),
.B2(n_1663),
.Y(n_1933)
);

NAND3xp33_ASAP7_75t_SL g1934 ( 
.A(n_1911),
.B(n_1881),
.C(n_1873),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1913),
.B(n_1870),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1924),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1917),
.B(n_1870),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1907),
.B(n_1906),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1907),
.B(n_1873),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1914),
.B(n_1881),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1928),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1926),
.B(n_1893),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1918),
.B(n_1884),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1929),
.B(n_1884),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1924),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_SL g1946 ( 
.A(n_1925),
.B(n_1895),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1919),
.B(n_1893),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1931),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1906),
.B(n_1893),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1908),
.B(n_1889),
.Y(n_1950)
);

AOI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1909),
.A2(n_1892),
.B1(n_1823),
.B2(n_1857),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1912),
.B(n_1892),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1908),
.B(n_1891),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1929),
.B(n_1848),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1905),
.A2(n_1848),
.B1(n_1824),
.B2(n_1828),
.Y(n_1955)
);

INVxp67_ASAP7_75t_L g1956 ( 
.A(n_1932),
.Y(n_1956)
);

AOI221xp5_ASAP7_75t_L g1957 ( 
.A1(n_1934),
.A2(n_1956),
.B1(n_1952),
.B2(n_1954),
.C(n_1938),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1942),
.B(n_1920),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1940),
.B(n_1910),
.Y(n_1959)
);

AOI21xp33_ASAP7_75t_SL g1960 ( 
.A1(n_1944),
.A2(n_1933),
.B(n_1932),
.Y(n_1960)
);

OAI222xp33_ASAP7_75t_L g1961 ( 
.A1(n_1952),
.A2(n_1915),
.B1(n_1933),
.B2(n_1891),
.C1(n_1903),
.C2(n_1894),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_SL g1962 ( 
.A1(n_1955),
.A2(n_1930),
.B(n_1921),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1951),
.A2(n_1940),
.B1(n_1948),
.B2(n_1954),
.Y(n_1963)
);

NOR3xp33_ASAP7_75t_L g1964 ( 
.A(n_1939),
.B(n_1922),
.C(n_1916),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1943),
.B(n_1903),
.Y(n_1965)
);

NAND4xp25_ASAP7_75t_L g1966 ( 
.A(n_1946),
.B(n_1927),
.C(n_1923),
.D(n_1898),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1942),
.A2(n_1896),
.B1(n_1862),
.B2(n_1858),
.Y(n_1967)
);

AOI21xp33_ASAP7_75t_L g1968 ( 
.A1(n_1941),
.A2(n_1945),
.B(n_1949),
.Y(n_1968)
);

AOI221xp5_ASAP7_75t_L g1969 ( 
.A1(n_1953),
.A2(n_1894),
.B1(n_1904),
.B2(n_1852),
.C(n_1855),
.Y(n_1969)
);

XNOR2xp5_ASAP7_75t_L g1970 ( 
.A(n_1949),
.B(n_1813),
.Y(n_1970)
);

NAND2x1p5_ASAP7_75t_L g1971 ( 
.A(n_1959),
.B(n_1945),
.Y(n_1971)
);

NOR4xp25_ASAP7_75t_L g1972 ( 
.A(n_1957),
.B(n_1936),
.C(n_1935),
.D(n_1937),
.Y(n_1972)
);

NAND4xp25_ASAP7_75t_L g1973 ( 
.A(n_1968),
.B(n_1947),
.C(n_1936),
.D(n_1935),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1963),
.B(n_1947),
.Y(n_1974)
);

OAI21xp5_ASAP7_75t_L g1975 ( 
.A1(n_1962),
.A2(n_1937),
.B(n_1950),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1966),
.B(n_1950),
.Y(n_1976)
);

NAND5xp2_ASAP7_75t_L g1977 ( 
.A(n_1958),
.B(n_1855),
.C(n_1863),
.D(n_1860),
.E(n_1815),
.Y(n_1977)
);

NOR3xp33_ASAP7_75t_SL g1978 ( 
.A(n_1961),
.B(n_1970),
.C(n_1969),
.Y(n_1978)
);

NOR2x1_ASAP7_75t_L g1979 ( 
.A(n_1965),
.B(n_1904),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1964),
.B(n_1819),
.Y(n_1980)
);

NAND3x1_ASAP7_75t_L g1981 ( 
.A(n_1967),
.B(n_1863),
.C(n_1777),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1960),
.B(n_1800),
.Y(n_1982)
);

NOR3xp33_ASAP7_75t_SL g1983 ( 
.A(n_1963),
.B(n_1750),
.C(n_1743),
.Y(n_1983)
);

AND4x1_ASAP7_75t_L g1984 ( 
.A(n_1974),
.B(n_1808),
.C(n_1800),
.D(n_1801),
.Y(n_1984)
);

OAI211xp5_ASAP7_75t_SL g1985 ( 
.A1(n_1978),
.A2(n_1975),
.B(n_1976),
.C(n_1983),
.Y(n_1985)
);

AOI211xp5_ASAP7_75t_SL g1986 ( 
.A1(n_1982),
.A2(n_1833),
.B(n_1832),
.C(n_1830),
.Y(n_1986)
);

NAND4xp25_ASAP7_75t_L g1987 ( 
.A(n_1973),
.B(n_1833),
.C(n_1832),
.D(n_1830),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1972),
.B(n_1832),
.Y(n_1988)
);

NOR4xp75_ASAP7_75t_L g1989 ( 
.A(n_1981),
.B(n_1750),
.C(n_1767),
.D(n_1759),
.Y(n_1989)
);

NAND4xp25_ASAP7_75t_SL g1990 ( 
.A(n_1980),
.B(n_1833),
.C(n_1818),
.D(n_1816),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1973),
.B(n_1801),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1988),
.Y(n_1992)
);

NOR2x1_ASAP7_75t_L g1993 ( 
.A(n_1985),
.B(n_1979),
.Y(n_1993)
);

NOR2xp67_ASAP7_75t_SL g1994 ( 
.A(n_1991),
.B(n_1971),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1984),
.B(n_1977),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1987),
.Y(n_1996)
);

NOR2x1_ASAP7_75t_L g1997 ( 
.A(n_1990),
.B(n_1818),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1989),
.A2(n_1818),
.B1(n_1799),
.B2(n_1789),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1995),
.B(n_1986),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1997),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1993),
.Y(n_2001)
);

NOR4xp25_ASAP7_75t_L g2002 ( 
.A(n_1996),
.B(n_1799),
.C(n_1789),
.D(n_1738),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1994),
.B(n_1793),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1992),
.A2(n_1799),
.B(n_1789),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_2001),
.B(n_1998),
.Y(n_2005)
);

NAND4xp75_ASAP7_75t_L g2006 ( 
.A(n_1999),
.B(n_1740),
.C(n_1793),
.D(n_1812),
.Y(n_2006)
);

NOR3xp33_ASAP7_75t_L g2007 ( 
.A(n_2000),
.B(n_1576),
.C(n_1608),
.Y(n_2007)
);

AND2x2_ASAP7_75t_SL g2008 ( 
.A(n_2003),
.B(n_1770),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_2005),
.Y(n_2009)
);

NOR3xp33_ASAP7_75t_L g2010 ( 
.A(n_2009),
.B(n_2007),
.C(n_2006),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_2010),
.Y(n_2011)
);

XNOR2xp5_ASAP7_75t_L g2012 ( 
.A(n_2010),
.B(n_2008),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_2012),
.B(n_2002),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_2011),
.Y(n_2014)
);

OAI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_2013),
.A2(n_2002),
.B(n_2004),
.Y(n_2015)
);

OAI21xp5_ASAP7_75t_L g2016 ( 
.A1(n_2014),
.A2(n_1808),
.B(n_1806),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_2015),
.B(n_1740),
.Y(n_2017)
);

XNOR2xp5_ASAP7_75t_L g2018 ( 
.A(n_2017),
.B(n_2016),
.Y(n_2018)
);

AOI221xp5_ASAP7_75t_L g2019 ( 
.A1(n_2018),
.A2(n_1746),
.B1(n_1747),
.B2(n_1806),
.C(n_1809),
.Y(n_2019)
);

AOI211xp5_ASAP7_75t_L g2020 ( 
.A1(n_2019),
.A2(n_1609),
.B(n_1747),
.C(n_1608),
.Y(n_2020)
);


endmodule