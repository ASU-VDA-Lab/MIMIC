module fake_netlist_6_2056_n_46 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_8, n_46);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_8;

output n_46;

wire n_41;
wire n_16;
wire n_45;
wire n_34;
wire n_42;
wire n_9;
wire n_10;
wire n_21;
wire n_18;
wire n_24;
wire n_37;
wire n_15;
wire n_33;
wire n_27;
wire n_14;
wire n_38;
wire n_39;
wire n_32;
wire n_36;
wire n_22;
wire n_26;
wire n_13;
wire n_35;
wire n_11;
wire n_28;
wire n_23;
wire n_17;
wire n_12;
wire n_20;
wire n_30;
wire n_43;
wire n_19;
wire n_29;
wire n_31;
wire n_25;
wire n_40;
wire n_44;

BUFx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

HB1xp67_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

AND2x4_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_4),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_13),
.Y(n_21)
);

NAND2xp33_ASAP7_75t_SL g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_R g24 ( 
.A(n_22),
.B(n_14),
.Y(n_24)
);

CKINVDCx11_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_14),
.B(n_2),
.Y(n_27)
);

AO21x2_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_23),
.B(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVxp67_ASAP7_75t_SL g31 ( 
.A(n_26),
.Y(n_31)
);

OAI221xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_18),
.B1(n_19),
.B2(n_17),
.C(n_8),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_17),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_17),
.B1(n_25),
.B2(n_8),
.Y(n_34)
);

NAND3xp33_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_1),
.C(n_5),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_31),
.B(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_35),
.A3(n_31),
.B1(n_29),
.B2(n_28),
.C1(n_32),
.C2(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_28),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_28),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_28),
.B1(n_38),
.B2(n_40),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_28),
.B1(n_43),
.B2(n_41),
.Y(n_46)
);


endmodule