module real_jpeg_17161_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_2),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_2),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_3),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_3),
.A2(n_85),
.B1(n_101),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_3),
.A2(n_85),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_85),
.B1(n_181),
.B2(n_184),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_4),
.A2(n_148),
.B1(n_189),
.B2(n_192),
.Y(n_188)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_4),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_5),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_5),
.Y(n_307)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_6),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_6),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g313 ( 
.A(n_6),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_8),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_8),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_8),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_8),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_8),
.Y(n_125)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_9),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_9),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_9),
.A2(n_41),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_9),
.B(n_162),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_9),
.A2(n_54),
.A3(n_209),
.B1(n_211),
.B2(n_214),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_9),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_9),
.B(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_10),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_11),
.Y(n_98)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_294),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_200),
.B(n_292),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_169),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_16),
.B(n_169),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.C(n_159),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_17),
.B(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_89),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_50),
.B2(n_51),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_20),
.B(n_50),
.C(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_38),
.B(n_39),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AO22x2_ASAP7_75t_L g179 ( 
.A1(n_22),
.A2(n_32),
.B1(n_40),
.B2(n_180),
.Y(n_179)
);

AO22x1_ASAP7_75t_L g224 ( 
.A1(n_22),
.A2(n_32),
.B1(n_40),
.B2(n_180),
.Y(n_224)
);

NOR2x1p5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_32),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_26),
.Y(n_234)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AO22x2_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_32),
.B(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_34),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_35),
.Y(n_149)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_35),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_35),
.Y(n_156)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_35),
.Y(n_191)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_35),
.Y(n_306)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B(n_46),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_45),
.Y(n_185)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_45),
.Y(n_217)
);

OAI32xp33_ASAP7_75t_L g230 ( 
.A1(n_46),
.A2(n_231),
.A3(n_235),
.B1(n_237),
.B2(n_242),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_47),
.B(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_50),
.A2(n_51),
.B1(n_179),
.B2(n_196),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_50),
.B(n_179),
.C(n_207),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_68),
.B1(n_74),
.B2(n_81),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_52),
.A2(n_68),
.B1(n_74),
.B2(n_81),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_52),
.A2(n_68),
.B(n_74),
.Y(n_318)
);

NAND2x1p5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_68),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_60),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_68),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_71),
.Y(n_183)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx2_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_89),
.A2(n_90),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_90),
.Y(n_199)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_99),
.B1(n_109),
.B2(n_116),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_91),
.A2(n_99),
.B1(n_109),
.B2(n_116),
.Y(n_173)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_95),
.B(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_95),
.Y(n_265)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21x1_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_105),
.B(n_109),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_109)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_120),
.B(n_159),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_137),
.B2(n_138),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_137),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_137),
.A2(n_138),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_138),
.B(n_223),
.C(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_138),
.B(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_138),
.B(n_264),
.Y(n_266)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_147),
.B1(n_152),
.B2(n_154),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_139),
.A2(n_188),
.B1(n_304),
.B2(n_311),
.Y(n_303)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_155),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_140),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_143),
.Y(n_262)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_144),
.Y(n_236)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_146),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_164),
.B(n_168),
.Y(n_163)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.C(n_163),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_160),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_160),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_160),
.A2(n_172),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_160),
.B(n_173),
.C(n_175),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_161),
.A2(n_163),
.B1(n_268),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_161),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_163),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_163),
.Y(n_268)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_168),
.A2(n_188),
.B(n_193),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_170),
.B(n_178),
.C(n_197),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_173),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_197),
.B2(n_198),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_186),
.B1(n_187),
.B2(n_196),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_179),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_179),
.A2(n_196),
.B1(n_230),
.B2(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_179),
.B(n_187),
.Y(n_315)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_191),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_287),
.B(n_291),
.Y(n_202)
);

AOI21x1_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_274),
.B(n_286),
.Y(n_203)
);

OAI21x1_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_227),
.B(n_273),
.Y(n_204)
);

NOR2xp67_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_222),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_206),
.B(n_222),
.Y(n_273)
);

XOR2x2_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_221),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_208),
.B(n_218),
.Y(n_277)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_223),
.A2(n_224),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_223),
.B(n_277),
.C(n_279),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_223),
.A2(n_224),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_225),
.Y(n_250)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_251),
.B(n_272),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_248),
.Y(n_228)
);

NOR2xp67_ASAP7_75t_SL g272 ( 
.A(n_229),
.B(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21x1_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_267),
.B(n_271),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_263),
.B(n_266),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_285),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_285),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_279),
.B1(n_280),
.B2(n_284),
.Y(n_275)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_276),
.Y(n_284)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_289),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_319),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2x1_ASAP7_75t_SL g320 ( 
.A(n_297),
.B(n_298),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_314),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx6_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2x1_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);


endmodule