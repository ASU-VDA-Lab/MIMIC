module fake_jpeg_19472_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx11_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_21),
.B(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_19),
.C(n_18),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_24),
.C(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_17),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_16),
.B(n_11),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_13),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_10),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_10),
.B1(n_23),
.B2(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_9),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_38),
.C(n_41),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_56),
.C(n_58),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_52),
.B1(n_50),
.B2(n_47),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_53),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_40),
.C(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_52),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_15),
.C(n_12),
.Y(n_65)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_65),
.B(n_6),
.Y(n_70)
);

FAx1_ASAP7_75t_SL g68 ( 
.A(n_67),
.B(n_61),
.CI(n_62),
.CON(n_68),
.SN(n_68)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_3),
.B(n_6),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.C(n_7),
.Y(n_72)
);

AO21x1_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_68),
.B(n_8),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_71),
.Y(n_74)
);


endmodule