module real_jpeg_25180_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_1),
.B(n_73),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_1),
.A2(n_24),
.B1(n_27),
.B2(n_30),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_1),
.B(n_35),
.C(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_1),
.B(n_47),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_1),
.A2(n_32),
.B1(n_120),
.B2(n_127),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx8_ASAP7_75t_SL g74 ( 
.A(n_4),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_5),
.A2(n_24),
.B1(n_30),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_5),
.A2(n_21),
.B1(n_22),
.B2(n_52),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_52),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_24),
.B1(n_30),
.B2(n_40),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_8),
.A2(n_21),
.B1(n_22),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_8),
.A2(n_24),
.B1(n_30),
.B2(n_49),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_49),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_9),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_11),
.A2(n_24),
.B1(n_30),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_61),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_13),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_94),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_93),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_62),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_18),
.B(n_62),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.C(n_50),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_19),
.B(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_20),
.B(n_31),
.Y(n_86)
);

OAI32xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.A3(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_21),
.A2(n_22),
.B1(n_25),
.B2(n_29),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_21),
.A2(n_22),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

HAxp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_27),
.CON(n_26),
.SN(n_26)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_24),
.Y(n_30)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_24),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_24),
.A2(n_30),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_24),
.B(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_27),
.B(n_58),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_27),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_38),
.B(n_41),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_32),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_32),
.A2(n_117),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_33),
.B(n_42),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_33),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_34),
.A2(n_35),
.B1(n_55),
.B2(n_57),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_34),
.B(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_37),
.Y(n_112)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_39),
.B(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_44),
.B(n_50),
.Y(n_141)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_51),
.A2(n_53),
.B1(n_59),
.B2(n_100),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_60),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_59),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_84),
.B2(n_85),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_70),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B(n_83),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_92),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_86),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_138),
.B(n_142),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_113),
.B(n_137),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_97),
.B(n_103),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_101),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_108),
.C(n_109),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_123),
.B(n_136),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_122),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_130),
.B(n_135),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_125),
.B(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_139),
.B(n_140),
.Y(n_142)
);


endmodule