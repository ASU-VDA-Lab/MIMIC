module real_aes_9172_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g190 ( .A1(n_0), .A2(n_191), .B(n_192), .C(n_196), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_1), .B(n_186), .Y(n_197) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_110), .C(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g447 ( .A(n_2), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_3), .B(n_151), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_4), .A2(n_132), .B(n_481), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_5), .A2(n_137), .B(n_142), .C(n_517), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_6), .A2(n_132), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_7), .B(n_186), .Y(n_487) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_8), .A2(n_165), .B(n_215), .Y(n_214) );
AND2x6_ASAP7_75t_L g137 ( .A(n_9), .B(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_10), .A2(n_137), .B(n_142), .C(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g542 ( .A(n_11), .Y(n_542) );
INVx1_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_12), .B(n_39), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_13), .B(n_195), .Y(n_519) );
INVx1_ASAP7_75t_L g161 ( .A(n_14), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_15), .B(n_151), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_16), .A2(n_152), .B(n_527), .C(n_529), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_17), .B(n_186), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_18), .B(n_179), .Y(n_571) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_19), .A2(n_142), .B(n_173), .C(n_178), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_20), .A2(n_194), .B(n_209), .C(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_21), .B(n_195), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_22), .A2(n_76), .B1(n_736), .B2(n_737), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_22), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_23), .B(n_195), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g468 ( .A(n_24), .Y(n_468) );
INVx1_ASAP7_75t_L g493 ( .A(n_25), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_26), .A2(n_142), .B(n_178), .C(n_218), .Y(n_217) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_27), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_28), .Y(n_515) );
INVx1_ASAP7_75t_L g569 ( .A(n_29), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_30), .A2(n_132), .B(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g135 ( .A(n_31), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_32), .A2(n_140), .B(n_145), .C(n_155), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_33), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_34), .A2(n_194), .B(n_484), .C(n_486), .Y(n_483) );
INVxp67_ASAP7_75t_L g570 ( .A(n_35), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_36), .B(n_220), .Y(n_219) );
CKINVDCx14_ASAP7_75t_R g482 ( .A(n_37), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_38), .A2(n_142), .B(n_178), .C(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_39), .B(n_107), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_40), .A2(n_196), .B(n_540), .C(n_541), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_41), .B(n_171), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_42), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_43), .B(n_151), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_44), .B(n_132), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_45), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_46), .Y(n_566) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_47), .A2(n_140), .B(n_155), .C(n_229), .Y(n_228) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_48), .A2(n_87), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_48), .Y(n_123) );
INVx1_ASAP7_75t_L g193 ( .A(n_49), .Y(n_193) );
INVx1_ASAP7_75t_L g230 ( .A(n_50), .Y(n_230) );
INVx1_ASAP7_75t_L g505 ( .A(n_51), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_52), .B(n_132), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_53), .Y(n_182) );
CKINVDCx14_ASAP7_75t_R g538 ( .A(n_54), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_55), .Y(n_450) );
INVx1_ASAP7_75t_L g138 ( .A(n_56), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_57), .B(n_132), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_58), .B(n_186), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_59), .A2(n_177), .B(n_240), .C(n_242), .Y(n_239) );
INVx1_ASAP7_75t_L g160 ( .A(n_60), .Y(n_160) );
INVx1_ASAP7_75t_SL g485 ( .A(n_61), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_62), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_63), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_64), .B(n_186), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_65), .B(n_152), .Y(n_206) );
INVx1_ASAP7_75t_L g471 ( .A(n_66), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_67), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_68), .B(n_148), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_69), .A2(n_142), .B(n_155), .C(n_266), .Y(n_265) );
CKINVDCx16_ASAP7_75t_R g238 ( .A(n_70), .Y(n_238) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_72), .A2(n_132), .B(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_73), .A2(n_102), .B1(n_114), .B2(n_748), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_74), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_75), .A2(n_132), .B(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_76), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_77), .A2(n_171), .B(n_565), .Y(n_564) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_78), .Y(n_490) );
INVx1_ASAP7_75t_L g525 ( .A(n_79), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_80), .B(n_147), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_81), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_82), .A2(n_132), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g528 ( .A(n_83), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_84), .Y(n_747) );
INVx2_ASAP7_75t_L g158 ( .A(n_85), .Y(n_158) );
INVx1_ASAP7_75t_L g518 ( .A(n_86), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_87), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_88), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_89), .B(n_195), .Y(n_207) );
INVx2_ASAP7_75t_L g110 ( .A(n_90), .Y(n_110) );
OR2x2_ASAP7_75t_L g444 ( .A(n_90), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g455 ( .A(n_90), .B(n_446), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_91), .A2(n_142), .B(n_155), .C(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_92), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g146 ( .A(n_93), .Y(n_146) );
INVxp67_ASAP7_75t_L g243 ( .A(n_94), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_95), .B(n_165), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_96), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g202 ( .A(n_97), .Y(n_202) );
INVx1_ASAP7_75t_L g267 ( .A(n_98), .Y(n_267) );
INVx2_ASAP7_75t_L g508 ( .A(n_99), .Y(n_508) );
AND2x2_ASAP7_75t_L g232 ( .A(n_100), .B(n_157), .Y(n_232) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g748 ( .A(n_104), .Y(n_748) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g458 ( .A(n_110), .B(n_446), .Y(n_458) );
NOR2x2_ASAP7_75t_L g746 ( .A(n_110), .B(n_445), .Y(n_746) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OAI21x1_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_119), .B(n_451), .Y(n_114) );
OAI21xp5_ASAP7_75t_SL g451 ( .A1(n_115), .A2(n_449), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_442), .B(n_449), .Y(n_119) );
XOR2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
INVx2_ASAP7_75t_L g456 ( .A(n_124), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_124), .A2(n_739), .B1(n_742), .B2(n_743), .Y(n_738) );
OR3x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_356), .C(n_399), .Y(n_124) );
NAND5xp2_ASAP7_75t_L g125 ( .A(n_126), .B(n_283), .C(n_313), .D(n_330), .E(n_345), .Y(n_125) );
AOI221xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_198), .B1(n_245), .B2(n_251), .C(n_255), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_167), .Y(n_127) );
OR2x2_ASAP7_75t_L g260 ( .A(n_128), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g300 ( .A(n_128), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g318 ( .A(n_128), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_128), .B(n_253), .Y(n_335) );
OR2x2_ASAP7_75t_L g347 ( .A(n_128), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_128), .B(n_306), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_128), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_128), .B(n_284), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_128), .B(n_292), .Y(n_398) );
AND2x2_ASAP7_75t_L g430 ( .A(n_128), .B(n_184), .Y(n_430) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_128), .Y(n_438) );
INVx5_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_129), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g257 ( .A(n_129), .B(n_233), .Y(n_257) );
BUFx2_ASAP7_75t_L g280 ( .A(n_129), .Y(n_280) );
AND2x2_ASAP7_75t_L g309 ( .A(n_129), .B(n_168), .Y(n_309) );
AND2x2_ASAP7_75t_L g364 ( .A(n_129), .B(n_261), .Y(n_364) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_162), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_139), .B(n_157), .Y(n_130) );
BUFx2_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NAND2x1p5_ASAP7_75t_L g203 ( .A(n_133), .B(n_137), .Y(n_203) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
INVx1_ASAP7_75t_L g210 ( .A(n_135), .Y(n_210) );
INVx1_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_136), .Y(n_152) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_136), .Y(n_195) );
INVx1_ASAP7_75t_L g220 ( .A(n_136), .Y(n_220) );
INVx4_ASAP7_75t_SL g156 ( .A(n_137), .Y(n_156) );
BUFx3_ASAP7_75t_L g178 ( .A(n_137), .Y(n_178) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_SL g188 ( .A1(n_141), .A2(n_156), .B(n_189), .C(n_190), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_141), .A2(n_156), .B(n_238), .C(n_239), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_141), .A2(n_156), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_141), .A2(n_156), .B(n_505), .C(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_SL g524 ( .A1(n_141), .A2(n_156), .B(n_525), .C(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_SL g537 ( .A1(n_141), .A2(n_156), .B(n_538), .C(n_539), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_SL g565 ( .A1(n_141), .A2(n_156), .B(n_566), .C(n_567), .Y(n_565) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx3_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_143), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_150), .C(n_153), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_147), .A2(n_153), .B(n_230), .C(n_231), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_147), .A2(n_471), .B(n_472), .C(n_473), .Y(n_470) );
O2A1O1Ixp5_ASAP7_75t_L g517 ( .A1(n_147), .A2(n_473), .B(n_518), .C(n_519), .Y(n_517) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx4_ASAP7_75t_L g241 ( .A(n_149), .Y(n_241) );
INVx2_ASAP7_75t_L g191 ( .A(n_151), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_151), .B(n_243), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_151), .A2(n_176), .B(n_493), .C(n_494), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g568 ( .A1(n_151), .A2(n_241), .B1(n_569), .B2(n_570), .Y(n_568) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_152), .B(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
INVx1_ASAP7_75t_L g529 ( .A(n_154), .Y(n_529) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
INVx1_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_157), .A2(n_227), .B(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_157), .A2(n_203), .B(n_490), .C(n_491), .Y(n_489) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_157), .A2(n_536), .B(n_543), .Y(n_535) );
AND2x2_ASAP7_75t_SL g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AND2x2_ASAP7_75t_L g166 ( .A(n_158), .B(n_159), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
INVx3_ASAP7_75t_L g186 ( .A(n_164), .Y(n_186) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_164), .A2(n_201), .B(n_211), .Y(n_200) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_164), .A2(n_264), .B(n_272), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_164), .B(n_273), .Y(n_272) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_164), .A2(n_467), .B(n_474), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_164), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_164), .B(n_521), .Y(n_520) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_165), .A2(n_216), .B(n_217), .Y(n_215) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_165), .Y(n_235) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_167), .B(n_318), .Y(n_327) );
OAI32xp33_ASAP7_75t_L g341 ( .A1(n_167), .A2(n_277), .A3(n_342), .B1(n_343), .B2(n_344), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_167), .B(n_343), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_167), .B(n_260), .Y(n_384) );
INVx1_ASAP7_75t_SL g413 ( .A(n_167), .Y(n_413) );
NAND4xp25_ASAP7_75t_L g422 ( .A(n_167), .B(n_200), .C(n_364), .D(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_184), .Y(n_167) );
INVx5_ASAP7_75t_L g254 ( .A(n_168), .Y(n_254) );
AND2x2_ASAP7_75t_L g284 ( .A(n_168), .B(n_185), .Y(n_284) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_168), .Y(n_363) );
AND2x2_ASAP7_75t_L g433 ( .A(n_168), .B(n_380), .Y(n_433) );
OR2x6_ASAP7_75t_L g168 ( .A(n_169), .B(n_181), .Y(n_168) );
AOI21xp5_ASAP7_75t_SL g169 ( .A1(n_170), .A2(n_172), .B(n_179), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_176), .Y(n_173) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_177), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_180), .B(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_183), .A2(n_514), .B(n_520), .Y(n_513) );
AND2x4_ASAP7_75t_L g306 ( .A(n_184), .B(n_254), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_184), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g340 ( .A(n_184), .B(n_261), .Y(n_340) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g253 ( .A(n_185), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g292 ( .A(n_185), .B(n_263), .Y(n_292) );
AND2x2_ASAP7_75t_L g301 ( .A(n_185), .B(n_262), .Y(n_301) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_197), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_194), .B(n_485), .Y(n_484) );
INVx4_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g540 ( .A(n_195), .Y(n_540) );
INVx2_ASAP7_75t_L g473 ( .A(n_196), .Y(n_473) );
AOI222xp33_ASAP7_75t_L g369 ( .A1(n_198), .A2(n_370), .B1(n_372), .B2(n_374), .C1(n_377), .C2(n_378), .Y(n_369) );
AND2x4_ASAP7_75t_L g198 ( .A(n_199), .B(n_222), .Y(n_198) );
AND2x2_ASAP7_75t_L g302 ( .A(n_199), .B(n_303), .Y(n_302) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_199), .B(n_280), .C(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_214), .Y(n_199) );
INVx5_ASAP7_75t_SL g250 ( .A(n_200), .Y(n_250) );
OAI322xp33_ASAP7_75t_L g255 ( .A1(n_200), .A2(n_256), .A3(n_258), .B1(n_259), .B2(n_274), .C1(n_277), .C2(n_279), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_200), .B(n_248), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_200), .B(n_234), .Y(n_428) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_204), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_203), .A2(n_468), .B(n_469), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_203), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_208), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_208), .A2(n_219), .B(n_221), .Y(n_218) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
INVx2_ASAP7_75t_L g563 ( .A(n_213), .Y(n_563) );
INVx2_ASAP7_75t_L g248 ( .A(n_214), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_214), .B(n_224), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_222), .B(n_287), .Y(n_342) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OR2x2_ASAP7_75t_L g321 ( .A(n_223), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_233), .Y(n_223) );
OR2x2_ASAP7_75t_L g249 ( .A(n_224), .B(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_224), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g289 ( .A(n_224), .B(n_234), .Y(n_289) );
AND2x2_ASAP7_75t_L g312 ( .A(n_224), .B(n_248), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_224), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g328 ( .A(n_224), .B(n_287), .Y(n_328) );
AND2x2_ASAP7_75t_L g336 ( .A(n_224), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_224), .B(n_296), .Y(n_386) );
INVx5_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g276 ( .A(n_225), .B(n_250), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_225), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g303 ( .A(n_225), .B(n_234), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_225), .B(n_350), .Y(n_391) );
OR2x2_ASAP7_75t_L g407 ( .A(n_225), .B(n_351), .Y(n_407) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_225), .B(n_368), .Y(n_414) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_225), .Y(n_421) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_232), .Y(n_225) );
AND2x2_ASAP7_75t_L g275 ( .A(n_233), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g325 ( .A(n_233), .B(n_248), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_233), .B(n_250), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_233), .B(n_287), .Y(n_409) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_234), .B(n_250), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_234), .B(n_248), .Y(n_297) );
OR2x2_ASAP7_75t_L g351 ( .A(n_234), .B(n_248), .Y(n_351) );
AND2x2_ASAP7_75t_L g368 ( .A(n_234), .B(n_247), .Y(n_368) );
INVxp67_ASAP7_75t_L g390 ( .A(n_234), .Y(n_390) );
AND2x2_ASAP7_75t_L g417 ( .A(n_234), .B(n_287), .Y(n_417) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_234), .Y(n_424) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_244), .Y(n_234) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_235), .A2(n_480), .B(n_487), .Y(n_479) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_235), .A2(n_503), .B(n_509), .Y(n_502) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_235), .A2(n_523), .B(n_530), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_240), .A2(n_267), .B(n_268), .C(n_269), .Y(n_266) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_241), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_241), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_247), .B(n_298), .Y(n_371) );
INVx1_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g287 ( .A(n_248), .B(n_250), .Y(n_287) );
OR2x2_ASAP7_75t_L g354 ( .A(n_248), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g298 ( .A(n_249), .Y(n_298) );
OR2x2_ASAP7_75t_L g359 ( .A(n_249), .B(n_351), .Y(n_359) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g258 ( .A(n_253), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_253), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g259 ( .A(n_254), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_254), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_254), .B(n_261), .Y(n_294) );
INVx2_ASAP7_75t_L g339 ( .A(n_254), .Y(n_339) );
AND2x2_ASAP7_75t_L g352 ( .A(n_254), .B(n_292), .Y(n_352) );
AND2x2_ASAP7_75t_L g377 ( .A(n_254), .B(n_301), .Y(n_377) );
INVx1_ASAP7_75t_L g329 ( .A(n_259), .Y(n_329) );
INVx2_ASAP7_75t_SL g316 ( .A(n_260), .Y(n_316) );
INVx1_ASAP7_75t_L g319 ( .A(n_261), .Y(n_319) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_262), .Y(n_282) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g380 ( .A(n_263), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_271), .Y(n_264) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g486 ( .A(n_270), .Y(n_486) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g349 ( .A(n_276), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g355 ( .A(n_276), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_276), .A2(n_358), .B1(n_360), .B2(n_365), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_276), .B(n_368), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_277), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g311 ( .A(n_278), .Y(n_311) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
OR2x2_ASAP7_75t_L g293 ( .A(n_280), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_280), .B(n_284), .Y(n_344) );
AND2x2_ASAP7_75t_L g367 ( .A(n_280), .B(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g343 ( .A(n_282), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B(n_290), .C(n_304), .Y(n_283) );
INVx1_ASAP7_75t_L g307 ( .A(n_284), .Y(n_307) );
OAI221xp5_ASAP7_75t_SL g415 ( .A1(n_284), .A2(n_416), .B1(n_418), .B2(n_419), .C(n_422), .Y(n_415) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g434 ( .A(n_287), .Y(n_434) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g383 ( .A(n_289), .B(n_322), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_293), .B(n_295), .C(n_299), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OAI32xp33_ASAP7_75t_L g408 ( .A1(n_297), .A2(n_298), .A3(n_361), .B1(n_398), .B2(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
AND2x2_ASAP7_75t_L g440 ( .A(n_300), .B(n_339), .Y(n_440) );
AND2x2_ASAP7_75t_L g387 ( .A(n_301), .B(n_339), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_301), .B(n_309), .Y(n_405) );
AOI31xp33_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_307), .A3(n_308), .B(n_310), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_306), .B(n_318), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_306), .B(n_316), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_306), .A2(n_336), .B1(n_426), .B2(n_429), .C(n_431), .Y(n_425) );
CKINVDCx16_ASAP7_75t_R g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g331 ( .A(n_311), .B(n_332), .Y(n_331) );
AOI222xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_320), .B1(n_323), .B2(n_326), .C1(n_328), .C2(n_329), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g396 ( .A(n_315), .Y(n_396) );
INVx1_ASAP7_75t_L g418 ( .A(n_318), .Y(n_418) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_321), .A2(n_432), .B1(n_434), .B2(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g337 ( .A(n_322), .Y(n_337) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .B1(n_336), .B2(n_338), .C(n_341), .Y(n_330) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g375 ( .A(n_333), .B(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g427 ( .A(n_333), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g402 ( .A(n_338), .Y(n_402) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g366 ( .A(n_339), .Y(n_366) );
INVx1_ASAP7_75t_L g348 ( .A(n_340), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_343), .B(n_430), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_349), .B1(n_352), .B2(n_353), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g439 ( .A(n_352), .Y(n_439) );
INVxp33_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_354), .B(n_398), .Y(n_397) );
OAI32xp33_ASAP7_75t_L g388 ( .A1(n_355), .A2(n_389), .A3(n_390), .B1(n_391), .B2(n_392), .Y(n_388) );
NAND4xp25_ASAP7_75t_L g356 ( .A(n_357), .B(n_369), .C(n_381), .D(n_393), .Y(n_356) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
NAND2xp33_ASAP7_75t_SL g360 ( .A(n_361), .B(n_362), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_364), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
CKINVDCx16_ASAP7_75t_R g374 ( .A(n_375), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_378), .A2(n_394), .B1(n_411), .B2(n_414), .C(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g429 ( .A(n_380), .B(n_430), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B1(n_385), .B2(n_387), .C(n_388), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_390), .B(n_421), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g399 ( .A(n_400), .B(n_410), .C(n_425), .D(n_436), .Y(n_399) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_404), .B(n_406), .C(n_408), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g441 ( .A(n_428), .Y(n_441) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_440), .B(n_441), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
NOR2xp33_ASAP7_75t_SL g449 ( .A(n_444), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
OAI222xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_735), .B1(n_738), .B2(n_744), .C1(n_745), .C2(n_747), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_456), .B1(n_457), .B2(n_459), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g741 ( .A(n_455), .Y(n_741) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx6_ASAP7_75t_L g742 ( .A(n_458), .Y(n_742) );
INVx3_ASAP7_75t_L g743 ( .A(n_459), .Y(n_743) );
AND2x2_ASAP7_75t_SL g459 ( .A(n_460), .B(n_690), .Y(n_459) );
NOR4xp25_ASAP7_75t_L g460 ( .A(n_461), .B(n_627), .C(n_661), .D(n_677), .Y(n_460) );
NAND4xp25_ASAP7_75t_SL g461 ( .A(n_462), .B(n_556), .C(n_591), .D(n_607), .Y(n_461) );
AOI222xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_497), .B1(n_531), .B2(n_544), .C1(n_549), .C2(n_555), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AOI31xp33_ASAP7_75t_L g723 ( .A1(n_464), .A2(n_724), .A3(n_725), .B(n_727), .Y(n_723) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_476), .Y(n_464) );
AND2x2_ASAP7_75t_L g698 ( .A(n_465), .B(n_478), .Y(n_698) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g548 ( .A(n_466), .Y(n_548) );
AND2x2_ASAP7_75t_L g555 ( .A(n_466), .B(n_488), .Y(n_555) );
AND2x2_ASAP7_75t_L g612 ( .A(n_466), .B(n_479), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_476), .B(n_642), .Y(n_641) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_477), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_477), .B(n_559), .Y(n_602) );
AND2x2_ASAP7_75t_L g695 ( .A(n_477), .B(n_635), .Y(n_695) );
OAI321xp33_ASAP7_75t_L g729 ( .A1(n_477), .A2(n_548), .A3(n_702), .B1(n_730), .B2(n_732), .C(n_733), .Y(n_729) );
NAND4xp25_ASAP7_75t_L g733 ( .A(n_477), .B(n_534), .C(n_642), .D(n_734), .Y(n_733) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_488), .Y(n_477) );
AND2x2_ASAP7_75t_L g597 ( .A(n_478), .B(n_546), .Y(n_597) );
AND2x2_ASAP7_75t_L g616 ( .A(n_478), .B(n_548), .Y(n_616) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g547 ( .A(n_479), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g572 ( .A(n_479), .B(n_488), .Y(n_572) );
AND2x2_ASAP7_75t_L g658 ( .A(n_479), .B(n_546), .Y(n_658) );
INVx3_ASAP7_75t_SL g546 ( .A(n_488), .Y(n_546) );
AND2x2_ASAP7_75t_L g590 ( .A(n_488), .B(n_577), .Y(n_590) );
OR2x2_ASAP7_75t_L g623 ( .A(n_488), .B(n_548), .Y(n_623) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_488), .Y(n_630) );
AND2x2_ASAP7_75t_L g659 ( .A(n_488), .B(n_547), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_488), .B(n_632), .Y(n_674) );
AND2x2_ASAP7_75t_L g706 ( .A(n_488), .B(n_698), .Y(n_706) );
AND2x2_ASAP7_75t_L g715 ( .A(n_488), .B(n_560), .Y(n_715) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_495), .Y(n_488) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_510), .Y(n_498) );
INVx1_ASAP7_75t_SL g683 ( .A(n_499), .Y(n_683) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g551 ( .A(n_500), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g533 ( .A(n_501), .B(n_512), .Y(n_533) );
AND2x2_ASAP7_75t_L g619 ( .A(n_501), .B(n_535), .Y(n_619) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g589 ( .A(n_502), .B(n_522), .Y(n_589) );
OR2x2_ASAP7_75t_L g600 ( .A(n_502), .B(n_535), .Y(n_600) );
AND2x2_ASAP7_75t_L g626 ( .A(n_502), .B(n_535), .Y(n_626) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_502), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_510), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_510), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g599 ( .A(n_511), .B(n_600), .Y(n_599) );
AOI322xp5_ASAP7_75t_L g685 ( .A1(n_511), .A2(n_589), .A3(n_595), .B1(n_626), .B2(n_676), .C1(n_686), .C2(n_688), .Y(n_685) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_522), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_512), .B(n_534), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_512), .B(n_535), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_512), .B(n_552), .Y(n_606) );
AND2x2_ASAP7_75t_L g660 ( .A(n_512), .B(n_626), .Y(n_660) );
INVx1_ASAP7_75t_L g664 ( .A(n_512), .Y(n_664) );
AND2x2_ASAP7_75t_L g676 ( .A(n_512), .B(n_522), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_512), .B(n_551), .Y(n_708) );
INVx4_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g573 ( .A(n_513), .B(n_522), .Y(n_573) );
BUFx3_ASAP7_75t_L g587 ( .A(n_513), .Y(n_587) );
AND3x2_ASAP7_75t_L g669 ( .A(n_513), .B(n_649), .C(n_670), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_522), .B(n_533), .C(n_534), .Y(n_532) );
INVx1_ASAP7_75t_SL g552 ( .A(n_522), .Y(n_552) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_522), .Y(n_654) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g648 ( .A(n_533), .B(n_649), .Y(n_648) );
INVxp67_ASAP7_75t_L g655 ( .A(n_533), .Y(n_655) );
AND2x2_ASAP7_75t_L g693 ( .A(n_534), .B(n_671), .Y(n_693) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g574 ( .A(n_535), .Y(n_574) );
AND2x2_ASAP7_75t_L g649 ( .A(n_535), .B(n_552), .Y(n_649) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
OR2x2_ASAP7_75t_L g593 ( .A(n_546), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g712 ( .A(n_546), .B(n_612), .Y(n_712) );
AND2x2_ASAP7_75t_L g726 ( .A(n_546), .B(n_548), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_547), .B(n_560), .Y(n_667) );
AND2x2_ASAP7_75t_L g714 ( .A(n_547), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g577 ( .A(n_548), .B(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g594 ( .A(n_548), .B(n_560), .Y(n_594) );
INVx1_ASAP7_75t_L g604 ( .A(n_548), .Y(n_604) );
AND2x2_ASAP7_75t_L g635 ( .A(n_548), .B(n_560), .Y(n_635) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OAI221xp5_ASAP7_75t_L g677 ( .A1(n_550), .A2(n_678), .B1(n_682), .B2(n_684), .C(n_685), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_551), .B(n_553), .Y(n_550) );
AND2x2_ASAP7_75t_L g581 ( .A(n_551), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_554), .B(n_588), .Y(n_731) );
AOI322xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_573), .A3(n_574), .B1(n_575), .B2(n_581), .C1(n_583), .C2(n_590), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_572), .Y(n_558) );
NAND2x1p5_ASAP7_75t_L g611 ( .A(n_559), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_559), .B(n_622), .Y(n_621) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_559), .A2(n_572), .B(n_646), .C(n_647), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_559), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_559), .B(n_616), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_559), .B(n_698), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_559), .B(n_726), .Y(n_725) );
BUFx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_560), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_560), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g687 ( .A(n_560), .B(n_574), .Y(n_687) );
OA21x2_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .B(n_571), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AO21x2_ASAP7_75t_L g578 ( .A1(n_562), .A2(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g579 ( .A(n_564), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_571), .Y(n_580) );
INVx1_ASAP7_75t_L g662 ( .A(n_572), .Y(n_662) );
OAI31xp33_ASAP7_75t_L g672 ( .A1(n_572), .A2(n_597), .A3(n_673), .B(n_675), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_572), .B(n_578), .Y(n_724) );
INVx1_ASAP7_75t_SL g585 ( .A(n_573), .Y(n_585) );
AND2x2_ASAP7_75t_L g618 ( .A(n_573), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g699 ( .A(n_573), .B(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g584 ( .A(n_574), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g609 ( .A(n_574), .Y(n_609) );
AND2x2_ASAP7_75t_L g636 ( .A(n_574), .B(n_589), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_574), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g728 ( .A(n_574), .B(n_676), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_576), .B(n_646), .Y(n_719) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g615 ( .A(n_578), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g633 ( .A(n_578), .Y(n_633) );
NAND2xp33_ASAP7_75t_SL g583 ( .A(n_584), .B(n_586), .Y(n_583) );
OAI211xp5_ASAP7_75t_SL g627 ( .A1(n_585), .A2(n_628), .B(n_634), .C(n_650), .Y(n_627) );
OR2x2_ASAP7_75t_L g702 ( .A(n_585), .B(n_683), .Y(n_702) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
CKINVDCx16_ASAP7_75t_R g639 ( .A(n_587), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_587), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g608 ( .A(n_589), .B(n_609), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_595), .B(n_598), .C(n_601), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_SL g642 ( .A(n_594), .Y(n_642) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_597), .B(n_635), .Y(n_640) );
INVx1_ASAP7_75t_L g646 ( .A(n_597), .Y(n_646) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g605 ( .A(n_600), .B(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g638 ( .A(n_600), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g700 ( .A(n_600), .Y(n_700) );
AOI21xp33_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_603), .B(n_605), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_603), .A2(n_614), .B(n_617), .Y(n_613) );
AOI211xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B(n_613), .C(n_620), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_608), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_611), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_SL g624 ( .A(n_612), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g679 ( .A1(n_614), .A2(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_619), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g644 ( .A(n_619), .Y(n_644) );
AOI21xp33_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_624), .B(n_625), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g675 ( .A(n_626), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_632), .B(n_658), .Y(n_684) );
AND2x2_ASAP7_75t_L g697 ( .A(n_632), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g711 ( .A(n_632), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g721 ( .A(n_632), .B(n_659), .Y(n_721) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B(n_637), .C(n_645), .Y(n_634) );
INVx1_ASAP7_75t_L g681 ( .A(n_635), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B1(n_641), .B2(n_643), .Y(n_637) );
OR2x2_ASAP7_75t_L g643 ( .A(n_639), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_639), .B(n_700), .Y(n_722) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g716 ( .A(n_649), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_656), .B1(n_659), .B2(n_660), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g734 ( .A(n_654), .Y(n_734) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g680 ( .A(n_658), .Y(n_680) );
OAI211xp5_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_663), .B(n_665), .C(n_672), .Y(n_661) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx2_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_680), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NOR5xp2_ASAP7_75t_L g690 ( .A(n_691), .B(n_709), .C(n_717), .D(n_723), .E(n_729), .Y(n_690) );
OAI211xp5_ASAP7_75t_SL g691 ( .A1(n_692), .A2(n_694), .B(n_696), .C(n_703), .Y(n_691) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_699), .B(n_701), .Y(n_696) );
OAI21xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_706), .B(n_707), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_706), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI21xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_713), .B(n_716), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g732 ( .A(n_712), .Y(n_732) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B(n_722), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
CKINVDCx16_ASAP7_75t_R g744 ( .A(n_735), .Y(n_744) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx3_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
endmodule