module fake_netlist_5_970_n_1710 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1710);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1710;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1439;
wire n_1312;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx10_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_61),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_107),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_110),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_39),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_22),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_53),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_53),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_49),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_70),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_8),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_64),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_93),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_76),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_60),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_28),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_37),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_34),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_39),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_47),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_146),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_145),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_62),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_104),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_32),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_20),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_20),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_117),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_55),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_65),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_119),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_94),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_159),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_136),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_133),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_51),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_144),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_4),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_88),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_150),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_95),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_52),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_139),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_30),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_67),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_59),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_74),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_8),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_168),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_16),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_78),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_2),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_41),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_36),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_35),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_90),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_126),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_7),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_58),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_84),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_114),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_72),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_17),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_46),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_47),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_33),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_165),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_23),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_32),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_54),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_28),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_81),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_131),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_167),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_22),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_138),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_19),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_36),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_151),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_82),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_54),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_77),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_164),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_73),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_33),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_127),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_87),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_1),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_152),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_41),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_38),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_2),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_141),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_158),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_27),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_38),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_75),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_85),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_124),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_0),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_148),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_116),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_15),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_111),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_19),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_153),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_92),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_31),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_50),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_79),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_166),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_56),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_143),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_55),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_142),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_134),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_51),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_34),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_50),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_52),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_108),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_63),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_27),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_7),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_3),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_48),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_123),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_23),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_29),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_12),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_155),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_66),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_25),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_0),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_69),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_101),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_128),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_15),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_106),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_3),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_56),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_135),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_5),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_96),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_105),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_25),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_109),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_11),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_42),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_156),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_35),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_42),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_68),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_251),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_202),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_263),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_251),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_251),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_251),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_203),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_208),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_251),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_205),
.B(n_1),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_206),
.B(n_4),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_176),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_177),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_210),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_227),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_240),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_267),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_270),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_282),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_211),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_178),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_331),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_334),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_207),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_182),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_212),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_214),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_287),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_263),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_215),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_217),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_222),
.B(n_5),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_234),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_236),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_280),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_245),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_280),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_222),
.B(n_6),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_216),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_247),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_218),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_220),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_221),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_266),
.B(n_6),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_288),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_209),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_286),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_224),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_171),
.Y(n_387)
);

BUFx2_ASAP7_75t_SL g388 ( 
.A(n_294),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_177),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_173),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_176),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_300),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_301),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_306),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_311),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_324),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_179),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_327),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_206),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_180),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_294),
.B(n_9),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_177),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_180),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_186),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_186),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_188),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_226),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_188),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_196),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_230),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_232),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_196),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_198),
.B(n_9),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_268),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_198),
.B(n_10),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_175),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_336),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_R g422 ( 
.A(n_348),
.B(n_170),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_341),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_335),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_342),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_338),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_416),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_339),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_339),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_340),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_343),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_350),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_387),
.B(n_390),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_351),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_265),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_416),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_343),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_402),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_404),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_337),
.B(n_170),
.Y(n_443)
);

BUFx8_ASAP7_75t_L g444 ( 
.A(n_348),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_402),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_358),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_405),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_364),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_417),
.A2(n_370),
.B(n_328),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_337),
.B(n_172),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_337),
.B(n_172),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_373),
.B(n_265),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_381),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_SL g454 ( 
.A(n_347),
.B(n_179),
.Y(n_454)
);

INVxp33_ASAP7_75t_SL g455 ( 
.A(n_365),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_337),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_405),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_337),
.B(n_376),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_368),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_367),
.B(n_328),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_352),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_406),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_407),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_367),
.B(n_183),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_391),
.B(n_398),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_407),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_408),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_408),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_410),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_410),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_375),
.B(n_184),
.Y(n_472)
);

NAND2x1p5_ASAP7_75t_L g473 ( 
.A(n_415),
.B(n_237),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_411),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_411),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_347),
.B(n_185),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_414),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_414),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_403),
.B(n_174),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_383),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_353),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_377),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_359),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_379),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_380),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_344),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_355),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_359),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_362),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_412),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_344),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_362),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_413),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_357),
.B(n_223),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_483),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_483),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_456),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_456),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_420),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_436),
.B(n_479),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_488),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_488),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_489),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_458),
.B(n_452),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_466),
.B(n_389),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_422),
.Y(n_506)
);

INVx4_ASAP7_75t_SL g507 ( 
.A(n_476),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_476),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_489),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_492),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_456),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_492),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_420),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_420),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_424),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_473),
.A2(n_366),
.B1(n_386),
.B2(n_409),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_473),
.B(n_189),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_443),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_456),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_436),
.B(n_388),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_479),
.B(n_375),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_432),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_438),
.A2(n_382),
.B1(n_346),
.B2(n_399),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_452),
.B(n_443),
.Y(n_524)
);

INVx4_ASAP7_75t_SL g525 ( 
.A(n_476),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_424),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_L g527 ( 
.A(n_476),
.B(n_268),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_466),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_426),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_429),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_465),
.B(n_371),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_419),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_429),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_450),
.B(n_238),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_473),
.B(n_195),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_473),
.B(n_349),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_428),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_455),
.A2(n_360),
.B1(n_361),
.B2(n_292),
.Y(n_540)
);

NOR2x1p5_ASAP7_75t_L g541 ( 
.A(n_423),
.B(n_382),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_438),
.A2(n_369),
.B1(n_400),
.B2(n_399),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_428),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_451),
.B(n_401),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_476),
.B(n_241),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_427),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_432),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_SL g548 ( 
.A(n_461),
.B(n_250),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_476),
.B(n_253),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_438),
.B(n_442),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_421),
.B(n_273),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_430),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_476),
.A2(n_454),
.B1(n_449),
.B2(n_461),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_465),
.B(n_369),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_430),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_431),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_476),
.B(n_268),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_442),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_476),
.B(n_268),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_421),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_465),
.B(n_372),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_472),
.B(n_254),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_433),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_437),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_429),
.Y(n_565)
);

AND2x6_ASAP7_75t_L g566 ( 
.A(n_472),
.B(n_204),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_429),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_L g568 ( 
.A(n_429),
.B(n_268),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_472),
.B(n_372),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_461),
.B(n_255),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_433),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_429),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_431),
.Y(n_573)
);

BUFx4f_ASAP7_75t_L g574 ( 
.A(n_471),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g575 ( 
.A(n_494),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_435),
.B(n_374),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_429),
.B(n_257),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_439),
.B(n_264),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_471),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_441),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_441),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_439),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_446),
.A2(n_201),
.B1(n_192),
.B2(n_303),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_433),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_434),
.Y(n_585)
);

NAND2x1p5_ASAP7_75t_L g586 ( 
.A(n_449),
.B(n_213),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_439),
.B(n_274),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_471),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_439),
.B(n_278),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_494),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_L g591 ( 
.A(n_471),
.B(n_268),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_448),
.B(n_400),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_425),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_459),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_434),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_482),
.B(n_374),
.Y(n_596)
);

AND2x6_ASAP7_75t_L g597 ( 
.A(n_445),
.B(n_228),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_468),
.B(n_279),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_445),
.Y(n_599)
);

NOR2x1p5_ASAP7_75t_L g600 ( 
.A(n_484),
.B(n_485),
.Y(n_600)
);

BUFx4f_ASAP7_75t_L g601 ( 
.A(n_471),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_490),
.B(n_397),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_493),
.B(n_397),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_449),
.B(n_242),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_457),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_440),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_471),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_457),
.B(n_396),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_460),
.B(n_396),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_486),
.Y(n_610)
);

CKINVDCx11_ASAP7_75t_R g611 ( 
.A(n_462),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_468),
.B(n_478),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_468),
.B(n_283),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_425),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_486),
.B(n_268),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_486),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_460),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_440),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_463),
.B(n_378),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_L g620 ( 
.A1(n_463),
.A2(n_256),
.B1(n_219),
.B2(n_249),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_469),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_453),
.B(n_378),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_481),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_469),
.Y(n_624)
);

INVx4_ASAP7_75t_SL g625 ( 
.A(n_486),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_470),
.B(n_395),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_470),
.B(n_395),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_475),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_468),
.B(n_291),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_SL g630 ( 
.A(n_453),
.B(n_281),
.C(n_284),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_444),
.A2(n_201),
.B1(n_192),
.B2(n_312),
.Y(n_631)
);

AND2x2_ASAP7_75t_SL g632 ( 
.A(n_480),
.B(n_243),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_486),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_486),
.B(n_248),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_475),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_486),
.B(n_260),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_478),
.B(n_323),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_477),
.A2(n_393),
.B1(n_392),
.B2(n_385),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_478),
.B(n_477),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_500),
.B(n_478),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_500),
.B(n_444),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_495),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_518),
.B(n_447),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_622),
.B(n_480),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_576),
.B(n_444),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_551),
.B(n_298),
.Y(n_646)
);

BUFx5_ASAP7_75t_L g647 ( 
.A(n_597),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_518),
.B(n_521),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_553),
.A2(n_504),
.B1(n_557),
.B2(n_527),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_608),
.Y(n_650)
);

INVx8_ASAP7_75t_L g651 ( 
.A(n_566),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_521),
.B(n_447),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_576),
.B(n_444),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_592),
.B(n_259),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_520),
.B(n_174),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_560),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_528),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_582),
.Y(n_658)
);

NOR3xp33_ASAP7_75t_L g659 ( 
.A(n_506),
.B(n_296),
.C(n_308),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_524),
.B(n_464),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_582),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_538),
.B(n_190),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_561),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_538),
.B(n_191),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_554),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_499),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_596),
.B(n_259),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_544),
.B(n_467),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_602),
.B(n_292),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_505),
.B(n_385),
.Y(n_670)
);

AND2x6_ASAP7_75t_SL g671 ( 
.A(n_603),
.B(n_392),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_536),
.B(n_467),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_496),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_501),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_L g675 ( 
.A(n_566),
.B(n_268),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_523),
.B(n_303),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_502),
.B(n_474),
.Y(n_677)
);

AND2x2_ASAP7_75t_SL g678 ( 
.A(n_527),
.B(n_261),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_550),
.B(n_312),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_554),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_503),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_509),
.B(n_474),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_510),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_499),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_512),
.B(n_275),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_609),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_580),
.B(n_285),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_581),
.B(n_302),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_626),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_569),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_517),
.A2(n_326),
.B1(n_325),
.B2(n_318),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_517),
.A2(n_317),
.B1(n_316),
.B2(n_320),
.Y(n_692)
);

AO22x1_ASAP7_75t_L g693 ( 
.A1(n_516),
.A2(n_200),
.B1(n_199),
.B2(n_197),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_550),
.B(n_316),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_531),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_513),
.Y(n_696)
);

BUFx5_ASAP7_75t_L g697 ( 
.A(n_597),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_531),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_513),
.Y(n_699)
);

AND2x4_ASAP7_75t_SL g700 ( 
.A(n_533),
.B(n_487),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_599),
.B(n_313),
.Y(n_701)
);

NOR3xp33_ASAP7_75t_L g702 ( 
.A(n_630),
.B(n_317),
.C(n_318),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_523),
.B(n_259),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_583),
.B(n_320),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_514),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_590),
.B(n_393),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_632),
.B(n_169),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_632),
.B(n_169),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_553),
.A2(n_269),
.B1(n_332),
.B2(n_322),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_557),
.A2(n_252),
.B1(n_187),
.B2(n_181),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_608),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_608),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_542),
.B(n_169),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_531),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_627),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_570),
.B(n_225),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_605),
.B(n_491),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_537),
.A2(n_181),
.B1(n_193),
.B2(n_194),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_627),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_514),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_537),
.A2(n_297),
.B1(n_491),
.B2(n_394),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_562),
.A2(n_545),
.B1(n_549),
.B2(n_586),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_617),
.B(n_491),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_564),
.Y(n_724)
);

INVx5_ASAP7_75t_L g725 ( 
.A(n_597),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_548),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_621),
.B(n_624),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_564),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_559),
.A2(n_187),
.B1(n_244),
.B2(n_193),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_566),
.B(n_229),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_627),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_522),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_628),
.B(n_440),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_635),
.B(n_394),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_533),
.B(n_262),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_515),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_611),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_526),
.B(n_231),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_529),
.B(n_233),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_614),
.B(n_345),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_548),
.A2(n_297),
.B1(n_235),
.B2(n_239),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_534),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_539),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_533),
.B(n_262),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_586),
.A2(n_246),
.B1(n_258),
.B2(n_271),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_543),
.B(n_272),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_522),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_552),
.Y(n_748)
);

NOR2xp67_ASAP7_75t_L g749 ( 
.A(n_540),
.B(n_71),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_546),
.B(n_262),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_555),
.B(n_276),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_532),
.Y(n_752)
);

AND2x2_ASAP7_75t_SL g753 ( 
.A(n_559),
.B(n_356),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_631),
.B(n_289),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_556),
.B(n_290),
.Y(n_755)
);

BUFx2_ASAP7_75t_R g756 ( 
.A(n_558),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_620),
.B(n_305),
.Y(n_757)
);

BUFx5_ASAP7_75t_L g758 ( 
.A(n_597),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_573),
.B(n_356),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_598),
.B(n_354),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_613),
.B(n_194),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_629),
.B(n_354),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_546),
.B(n_305),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_558),
.B(n_99),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_498),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_637),
.B(n_197),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_619),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_593),
.B(n_304),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_639),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_541),
.B(n_345),
.Y(n_770)
);

OR2x6_ASAP7_75t_L g771 ( 
.A(n_600),
.B(n_330),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_578),
.B(n_199),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_587),
.B(n_244),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_604),
.A2(n_589),
.B1(n_577),
.B2(n_612),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_547),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_507),
.B(n_330),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_530),
.B(n_293),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_546),
.B(n_330),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_530),
.B(n_321),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_535),
.B(n_321),
.Y(n_780)
);

OAI22xp33_ASAP7_75t_L g781 ( 
.A1(n_619),
.A2(n_315),
.B1(n_314),
.B2(n_304),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_547),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_623),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_563),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_604),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_634),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_563),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_535),
.B(n_315),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_611),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_579),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_565),
.B(n_314),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_571),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_572),
.B(n_295),
.Y(n_793)
);

OR2x6_ASAP7_75t_L g794 ( 
.A(n_634),
.B(n_310),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_737),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_785),
.A2(n_497),
.B(n_618),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_660),
.A2(n_601),
.B(n_574),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_767),
.B(n_597),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_785),
.A2(n_649),
.B(n_640),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_649),
.A2(n_638),
.B1(n_299),
.B2(n_307),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_767),
.B(n_572),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_665),
.A2(n_606),
.B(n_595),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_655),
.A2(n_636),
.B(n_568),
.C(n_615),
.Y(n_803)
);

CKINVDCx10_ASAP7_75t_R g804 ( 
.A(n_771),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_672),
.A2(n_574),
.B(n_601),
.Y(n_805)
);

INVx5_ASAP7_75t_L g806 ( 
.A(n_651),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_650),
.B(n_507),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_665),
.B(n_571),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_787),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_655),
.A2(n_568),
.B(n_615),
.C(n_633),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_680),
.B(n_575),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_680),
.B(n_584),
.Y(n_812)
);

AO21x1_ASAP7_75t_L g813 ( 
.A1(n_662),
.A2(n_591),
.B(n_616),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_648),
.B(n_584),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_700),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_722),
.A2(n_595),
.B(n_585),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_657),
.B(n_575),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_711),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_657),
.B(n_567),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_753),
.A2(n_610),
.B(n_616),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_787),
.Y(n_821)
);

NAND2x1p5_ASAP7_75t_L g822 ( 
.A(n_650),
.B(n_579),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_666),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_684),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_695),
.B(n_525),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_753),
.A2(n_610),
.B(n_519),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_769),
.B(n_511),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_783),
.Y(n_828)
);

BUFx4f_ASAP7_75t_L g829 ( 
.A(n_771),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_650),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_774),
.A2(n_519),
.B(n_498),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_765),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_698),
.B(n_525),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_714),
.B(n_525),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_668),
.A2(n_588),
.B(n_607),
.Y(n_835)
);

NOR2xp67_ASAP7_75t_L g836 ( 
.A(n_656),
.B(n_638),
.Y(n_836)
);

OAI21x1_ASAP7_75t_L g837 ( 
.A1(n_696),
.A2(n_633),
.B(n_625),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_699),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_678),
.A2(n_607),
.B(n_309),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_678),
.A2(n_607),
.B(n_309),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_716),
.B(n_588),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_690),
.A2(n_607),
.B(n_307),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_705),
.A2(n_732),
.B(n_720),
.Y(n_843)
);

AO22x1_ASAP7_75t_L g844 ( 
.A1(n_703),
.A2(n_299),
.B1(n_310),
.B2(n_12),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_716),
.B(n_625),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_761),
.B(n_10),
.Y(n_846)
);

O2A1O1Ixp5_ASAP7_75t_L g847 ( 
.A1(n_664),
.A2(n_727),
.B(n_766),
.C(n_761),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_790),
.A2(n_112),
.B(n_163),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_SL g849 ( 
.A1(n_707),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_790),
.A2(n_725),
.B(n_765),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_725),
.A2(n_102),
.B(n_147),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_725),
.A2(n_100),
.B(n_132),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_766),
.B(n_13),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_725),
.A2(n_765),
.B(n_762),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_726),
.A2(n_310),
.B(n_130),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_747),
.Y(n_856)
);

AO21x1_ASAP7_75t_L g857 ( 
.A1(n_708),
.A2(n_14),
.B(n_16),
.Y(n_857)
);

CKINVDCx8_ASAP7_75t_R g858 ( 
.A(n_671),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_658),
.Y(n_859)
);

NAND2x1_ASAP7_75t_L g860 ( 
.A(n_765),
.B(n_129),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_726),
.B(n_17),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_644),
.B(n_18),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_679),
.A2(n_694),
.B(n_772),
.C(n_712),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_760),
.A2(n_125),
.B(n_122),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_772),
.B(n_18),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_SL g866 ( 
.A1(n_676),
.A2(n_21),
.B(n_24),
.C(n_26),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_786),
.A2(n_651),
.B(n_661),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_651),
.A2(n_120),
.B(n_98),
.Y(n_868)
);

NOR2x1_ASAP7_75t_R g869 ( 
.A(n_789),
.B(n_21),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_752),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_679),
.A2(n_24),
.B(n_26),
.C(n_29),
.Y(n_871)
);

INVx5_ASAP7_75t_L g872 ( 
.A(n_776),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_677),
.A2(n_97),
.B(n_91),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_770),
.Y(n_874)
);

AOI21x1_ASAP7_75t_L g875 ( 
.A1(n_733),
.A2(n_89),
.B(n_86),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_715),
.A2(n_83),
.B(n_31),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_740),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_719),
.A2(n_731),
.B(n_723),
.Y(n_878)
);

BUFx4f_ASAP7_75t_L g879 ( 
.A(n_771),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_682),
.A2(n_40),
.B(n_43),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_717),
.A2(n_40),
.B(n_43),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_770),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_694),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_663),
.B(n_686),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_689),
.B(n_642),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_675),
.A2(n_44),
.B(n_45),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_724),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_777),
.A2(n_780),
.B(n_779),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_764),
.B(n_49),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_673),
.B(n_57),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_710),
.A2(n_729),
.B1(n_749),
.B2(n_713),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_654),
.B(n_57),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_788),
.A2(n_773),
.B(n_793),
.Y(n_893)
);

O2A1O1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_718),
.A2(n_709),
.B(n_659),
.C(n_781),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_674),
.B(n_681),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_645),
.B(n_653),
.C(n_763),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_683),
.B(n_736),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_742),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_743),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_775),
.A2(n_792),
.B(n_782),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_748),
.Y(n_901)
);

INVx1_ASAP7_75t_SL g902 ( 
.A(n_706),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_784),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_791),
.A2(n_746),
.B(n_659),
.C(n_667),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_730),
.A2(n_685),
.B(n_688),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_687),
.A2(n_701),
.B(n_738),
.Y(n_906)
);

AOI22x1_ASAP7_75t_L g907 ( 
.A1(n_670),
.A2(n_646),
.B1(n_768),
.B2(n_744),
.Y(n_907)
);

AO22x1_ASAP7_75t_L g908 ( 
.A1(n_702),
.A2(n_750),
.B1(n_735),
.B2(n_745),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_740),
.B(n_710),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_739),
.A2(n_751),
.B(n_755),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_759),
.Y(n_911)
);

OAI21xp33_ASAP7_75t_L g912 ( 
.A1(n_729),
.A2(n_746),
.B(n_741),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_734),
.A2(n_669),
.B(n_754),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_721),
.B(n_718),
.Y(n_914)
);

AO21x1_ASAP7_75t_L g915 ( 
.A1(n_641),
.A2(n_757),
.B(n_704),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_647),
.B(n_758),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_728),
.B(n_794),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_794),
.A2(n_781),
.B1(n_692),
.B2(n_691),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_702),
.A2(n_794),
.B(n_776),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_778),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_693),
.B(n_756),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_647),
.A2(n_697),
.B(n_758),
.C(n_776),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_647),
.B(n_697),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_647),
.A2(n_697),
.B1(n_758),
.B2(n_776),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_697),
.Y(n_925)
);

AOI21x1_ASAP7_75t_L g926 ( 
.A1(n_652),
.A2(n_577),
.B(n_643),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_774),
.A2(n_722),
.B(n_787),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_655),
.A2(n_500),
.B1(n_518),
.B2(n_678),
.Y(n_928)
);

OAI21x1_ASAP7_75t_L g929 ( 
.A1(n_774),
.A2(n_722),
.B(n_787),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_L g930 ( 
.A(n_662),
.B(n_655),
.C(n_576),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_660),
.A2(n_508),
.B(n_672),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_660),
.A2(n_508),
.B(n_672),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_660),
.A2(n_508),
.B(n_672),
.Y(n_933)
);

AOI21x1_ASAP7_75t_L g934 ( 
.A1(n_652),
.A2(n_577),
.B(n_643),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_660),
.A2(n_508),
.B(n_672),
.Y(n_935)
);

AND2x2_ASAP7_75t_SL g936 ( 
.A(n_700),
.B(n_703),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_660),
.A2(n_508),
.B(n_672),
.Y(n_937)
);

AOI21xp33_ASAP7_75t_L g938 ( 
.A1(n_655),
.A2(n_500),
.B(n_662),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_660),
.A2(n_508),
.B(n_672),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_660),
.A2(n_508),
.B(n_672),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_767),
.B(n_500),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_650),
.B(n_506),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_767),
.B(n_500),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_660),
.A2(n_508),
.B(n_672),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_650),
.B(n_506),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_654),
.B(n_592),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_767),
.B(n_500),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_665),
.A2(n_680),
.B(n_767),
.C(n_648),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_660),
.A2(n_508),
.B(n_672),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_665),
.B(n_506),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_711),
.Y(n_951)
);

NOR2xp67_ASAP7_75t_L g952 ( 
.A(n_657),
.B(n_594),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_649),
.A2(n_767),
.B1(n_678),
.B2(n_500),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_767),
.B(n_500),
.Y(n_954)
);

CKINVDCx8_ASAP7_75t_R g955 ( 
.A(n_671),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_652),
.A2(n_577),
.B(n_643),
.Y(n_956)
);

NOR2xp67_ASAP7_75t_L g957 ( 
.A(n_657),
.B(n_594),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_644),
.B(n_706),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_650),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_828),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_928),
.A2(n_930),
.B1(n_953),
.B2(n_941),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_903),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_938),
.A2(n_799),
.B(n_863),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_884),
.B(n_874),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_825),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_799),
.A2(n_841),
.B(n_803),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_943),
.B(n_947),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_954),
.B(n_938),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_809),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_795),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_898),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_950),
.B(n_811),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_946),
.B(n_902),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_958),
.B(n_817),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_894),
.A2(n_953),
.B(n_912),
.C(n_914),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_837),
.A2(n_843),
.B(n_831),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_931),
.A2(n_933),
.B(n_932),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_911),
.B(n_948),
.Y(n_978)
);

OA21x2_ASAP7_75t_L g979 ( 
.A1(n_927),
.A2(n_929),
.B(n_816),
.Y(n_979)
);

AOI21xp33_ASAP7_75t_L g980 ( 
.A1(n_891),
.A2(n_918),
.B(n_904),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_935),
.A2(n_939),
.B(n_937),
.Y(n_981)
);

AOI21xp33_ASAP7_75t_L g982 ( 
.A1(n_891),
.A2(n_918),
.B(n_847),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_808),
.B(n_812),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_881),
.A2(n_855),
.B(n_876),
.C(n_853),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_940),
.A2(n_949),
.B(n_944),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_L g986 ( 
.A(n_846),
.B(n_865),
.C(n_907),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_867),
.A2(n_826),
.B(n_926),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_910),
.B(n_915),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_887),
.Y(n_989)
);

OAI21x1_ASAP7_75t_L g990 ( 
.A1(n_934),
.A2(n_956),
.B(n_820),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_808),
.B(n_812),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_881),
.A2(n_855),
.B(n_876),
.C(n_861),
.Y(n_992)
);

AO21x1_ASAP7_75t_L g993 ( 
.A1(n_919),
.A2(n_893),
.B(n_798),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_885),
.B(n_895),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_896),
.A2(n_909),
.B1(n_942),
.B2(n_945),
.Y(n_995)
);

BUFx4f_ASAP7_75t_L g996 ( 
.A(n_874),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_885),
.B(n_897),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_899),
.B(n_901),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_884),
.B(n_908),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_810),
.A2(n_888),
.B(n_796),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_819),
.B(n_818),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_796),
.A2(n_814),
.B(n_878),
.Y(n_1002)
);

AO31x2_ASAP7_75t_L g1003 ( 
.A1(n_871),
.A2(n_922),
.A3(n_857),
.B(n_814),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_832),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_806),
.B(n_830),
.Y(n_1005)
);

O2A1O1Ixp5_ASAP7_75t_L g1006 ( 
.A1(n_905),
.A2(n_797),
.B(n_906),
.C(n_805),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_952),
.B(n_957),
.Y(n_1007)
);

NOR2xp67_ASAP7_75t_L g1008 ( 
.A(n_920),
.B(n_877),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_832),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_924),
.A2(n_872),
.B(n_801),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_883),
.A2(n_919),
.B(n_800),
.C(n_836),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_872),
.A2(n_923),
.B(n_916),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_SL g1013 ( 
.A1(n_913),
.A2(n_886),
.B(n_868),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_842),
.A2(n_951),
.B(n_840),
.C(n_839),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_815),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_874),
.Y(n_1016)
);

AOI21xp33_ASAP7_75t_L g1017 ( 
.A1(n_800),
.A2(n_842),
.B(n_840),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_835),
.A2(n_850),
.B(n_802),
.Y(n_1018)
);

INVx5_ASAP7_75t_L g1019 ( 
.A(n_832),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_806),
.A2(n_872),
.B1(n_959),
.B2(n_827),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_900),
.A2(n_854),
.B(n_822),
.Y(n_1021)
);

NAND2x1p5_ASAP7_75t_L g1022 ( 
.A(n_806),
.B(n_830),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_823),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_959),
.B(n_890),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_830),
.B(n_859),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_821),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_875),
.A2(n_859),
.B(n_807),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_839),
.A2(n_925),
.B(n_856),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_824),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_860),
.A2(n_870),
.B(n_838),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_848),
.A2(n_873),
.B(n_851),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_892),
.B(n_844),
.Y(n_1032)
);

AO31x2_ASAP7_75t_L g1033 ( 
.A1(n_880),
.A2(n_864),
.A3(n_852),
.B(n_877),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_889),
.B(n_882),
.Y(n_1034)
);

AO21x2_ASAP7_75t_L g1035 ( 
.A1(n_866),
.A2(n_849),
.B(n_825),
.Y(n_1035)
);

CKINVDCx6p67_ASAP7_75t_R g1036 ( 
.A(n_804),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_862),
.A2(n_829),
.B(n_879),
.C(n_917),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_833),
.A2(n_834),
.B(n_936),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_882),
.B(n_833),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_882),
.B(n_834),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_921),
.A2(n_829),
.B1(n_879),
.B2(n_858),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_869),
.A2(n_649),
.B(n_799),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_955),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_941),
.B(n_943),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_938),
.A2(n_930),
.B(n_912),
.C(n_894),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_928),
.A2(n_930),
.B1(n_953),
.B2(n_943),
.Y(n_1046)
);

BUFx2_ASAP7_75t_SL g1047 ( 
.A(n_952),
.Y(n_1047)
);

AOI21x1_ASAP7_75t_SL g1048 ( 
.A1(n_845),
.A2(n_853),
.B(n_846),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_941),
.B(n_943),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_938),
.A2(n_930),
.B(n_785),
.Y(n_1050)
);

AOI221xp5_ASAP7_75t_SL g1051 ( 
.A1(n_894),
.A2(n_718),
.B1(n_918),
.B2(n_912),
.C(n_800),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_799),
.A2(n_649),
.B(n_841),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_828),
.Y(n_1053)
);

AOI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_930),
.A2(n_938),
.B(n_912),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_898),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_799),
.A2(n_649),
.B(n_841),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_884),
.B(n_874),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_903),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_898),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_813),
.A2(n_953),
.A3(n_863),
.B(n_803),
.Y(n_1060)
);

AND3x4_ASAP7_75t_L g1061 ( 
.A(n_952),
.B(n_728),
.C(n_724),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_941),
.B(n_943),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_799),
.A2(n_649),
.B(n_841),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_825),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_938),
.A2(n_930),
.B(n_912),
.C(n_894),
.Y(n_1065)
);

AO31x2_ASAP7_75t_L g1066 ( 
.A1(n_813),
.A2(n_953),
.A3(n_863),
.B(n_803),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_837),
.A2(n_843),
.B(n_831),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_837),
.A2(n_843),
.B(n_831),
.Y(n_1068)
);

AO31x2_ASAP7_75t_L g1069 ( 
.A1(n_813),
.A2(n_953),
.A3(n_863),
.B(n_803),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_799),
.A2(n_649),
.B(n_841),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_832),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_837),
.A2(n_843),
.B(n_831),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_799),
.A2(n_649),
.B(n_841),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_799),
.A2(n_649),
.B(n_841),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_941),
.B(n_943),
.Y(n_1075)
);

BUFx4_ASAP7_75t_SL g1076 ( 
.A(n_815),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_837),
.A2(n_843),
.B(n_831),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_825),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_928),
.A2(n_930),
.B1(n_953),
.B2(n_943),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_941),
.B(n_943),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_903),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_828),
.Y(n_1082)
);

BUFx4f_ASAP7_75t_SL g1083 ( 
.A(n_815),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_837),
.A2(n_843),
.B(n_831),
.Y(n_1084)
);

NAND2xp33_ASAP7_75t_L g1085 ( 
.A(n_928),
.B(n_953),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_938),
.A2(n_930),
.B(n_785),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_941),
.B(n_943),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_799),
.A2(n_649),
.B(n_841),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_938),
.A2(n_930),
.B(n_785),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_941),
.B(n_943),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_837),
.A2(n_843),
.B(n_831),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_941),
.B(n_943),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_795),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_941),
.B(n_943),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_832),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_938),
.B(n_953),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_938),
.A2(n_930),
.B(n_785),
.Y(n_1097)
);

AO221x2_ASAP7_75t_L g1098 ( 
.A1(n_844),
.A2(n_918),
.B1(n_693),
.B2(n_891),
.C(n_781),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_837),
.A2(n_843),
.B(n_831),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1000),
.A2(n_988),
.B(n_966),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_964),
.B(n_1057),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_973),
.Y(n_1102)
);

AOI22x1_ASAP7_75t_L g1103 ( 
.A1(n_963),
.A2(n_1013),
.B1(n_1097),
.B2(n_1089),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_960),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_972),
.B(n_974),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_1053),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1010),
.A2(n_1056),
.B(n_1052),
.Y(n_1107)
);

AOI221xp5_ASAP7_75t_L g1108 ( 
.A1(n_1051),
.A2(n_1054),
.B1(n_980),
.B2(n_1017),
.C(n_972),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_964),
.B(n_1057),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_997),
.B(n_999),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_997),
.B(n_994),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_968),
.B(n_989),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_967),
.B(n_1044),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_1009),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1055),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_999),
.B(n_1082),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1007),
.B(n_1032),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_998),
.B(n_1045),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_992),
.A2(n_984),
.B1(n_975),
.B2(n_1080),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1098),
.A2(n_1085),
.B1(n_1061),
.B2(n_995),
.Y(n_1120)
);

NAND3xp33_ASAP7_75t_L g1121 ( 
.A(n_1065),
.B(n_984),
.C(n_992),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_970),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1049),
.B(n_1062),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_975),
.A2(n_1075),
.B1(n_1094),
.B2(n_1092),
.Y(n_1124)
);

INVxp67_ASAP7_75t_SL g1125 ( 
.A(n_1087),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_1083),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1090),
.B(n_983),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_991),
.B(n_961),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1059),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1098),
.A2(n_1061),
.B1(n_1046),
.B2(n_1079),
.Y(n_1130)
);

INVx5_ASAP7_75t_L g1131 ( 
.A(n_1009),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1093),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1050),
.B(n_1086),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1009),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_1009),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1010),
.A2(n_1052),
.B(n_1063),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1023),
.Y(n_1137)
);

NOR2x1_ASAP7_75t_SL g1138 ( 
.A(n_1004),
.B(n_1019),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1011),
.A2(n_1096),
.B1(n_1042),
.B2(n_1014),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1076),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_978),
.B(n_1042),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_993),
.A2(n_977),
.A3(n_981),
.B(n_985),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_996),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1029),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1056),
.A2(n_1063),
.B(n_1070),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1096),
.A2(n_982),
.B1(n_986),
.B2(n_1034),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_969),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1070),
.A2(n_1074),
.B(n_1088),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_1083),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_1016),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1011),
.A2(n_1037),
.B(n_1024),
.C(n_1001),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1073),
.A2(n_1088),
.B(n_1074),
.Y(n_1152)
);

AND2x2_ASAP7_75t_SL g1153 ( 
.A(n_996),
.B(n_1041),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_1076),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1037),
.B(n_1047),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1043),
.B(n_962),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1036),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1073),
.A2(n_1002),
.B(n_1006),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_1025),
.Y(n_1159)
);

INVx5_ASAP7_75t_L g1160 ( 
.A(n_1071),
.Y(n_1160)
);

NOR2x1_ASAP7_75t_SL g1161 ( 
.A(n_1004),
.B(n_1019),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1038),
.A2(n_1028),
.B(n_1030),
.C(n_1012),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1038),
.A2(n_965),
.B1(n_1064),
.B2(n_1078),
.Y(n_1163)
);

BUFx12f_ASAP7_75t_L g1164 ( 
.A(n_1015),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1008),
.B(n_1039),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_1040),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1026),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1064),
.A2(n_1078),
.B1(n_1081),
.B2(n_1058),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1071),
.B(n_1095),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1071),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1005),
.A2(n_1022),
.B1(n_1071),
.B2(n_1095),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1005),
.A2(n_1022),
.B1(n_1095),
.B2(n_1020),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1095),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1035),
.B(n_1060),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_979),
.A2(n_1060),
.B1(n_1069),
.B2(n_1066),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1003),
.Y(n_1176)
);

INVx5_ASAP7_75t_L g1177 ( 
.A(n_1048),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1027),
.Y(n_1178)
);

AND3x1_ASAP7_75t_SL g1179 ( 
.A(n_1048),
.B(n_1069),
.C(n_1003),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1069),
.B(n_1003),
.Y(n_1180)
);

BUFx12f_ASAP7_75t_L g1181 ( 
.A(n_1033),
.Y(n_1181)
);

NOR2x1_ASAP7_75t_L g1182 ( 
.A(n_979),
.B(n_1033),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1033),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1003),
.B(n_1033),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_SL g1185 ( 
.A1(n_1031),
.A2(n_1018),
.B1(n_987),
.B2(n_1021),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_990),
.Y(n_1186)
);

BUFx4f_ASAP7_75t_SL g1187 ( 
.A(n_976),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1067),
.Y(n_1188)
);

BUFx2_ASAP7_75t_SL g1189 ( 
.A(n_1068),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1072),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1077),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1084),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1091),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1099),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_971),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_992),
.A2(n_953),
.B1(n_928),
.B2(n_943),
.Y(n_1196)
);

OAI21xp33_ASAP7_75t_L g1197 ( 
.A1(n_972),
.A2(n_938),
.B(n_902),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_992),
.A2(n_938),
.B(n_930),
.C(n_912),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_973),
.B(n_946),
.Y(n_1199)
);

BUFx12f_ASAP7_75t_L g1200 ( 
.A(n_1015),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_968),
.B(n_941),
.Y(n_1201)
);

AO22x2_ASAP7_75t_L g1202 ( 
.A1(n_1096),
.A2(n_1079),
.B1(n_961),
.B2(n_1046),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_971),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_973),
.B(n_946),
.Y(n_1204)
);

INVx5_ASAP7_75t_SL g1205 ( 
.A(n_1036),
.Y(n_1205)
);

BUFx12f_ASAP7_75t_L g1206 ( 
.A(n_1015),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1053),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1053),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_970),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1053),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_997),
.B(n_994),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_1053),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_992),
.A2(n_984),
.B(n_975),
.Y(n_1213)
);

INVxp67_ASAP7_75t_SL g1214 ( 
.A(n_997),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_973),
.B(n_946),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_997),
.B(n_994),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_964),
.B(n_1057),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_964),
.B(n_1057),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1083),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_973),
.B(n_946),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1053),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_971),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_973),
.B(n_946),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_997),
.B(n_994),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_971),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_992),
.A2(n_953),
.B1(n_928),
.B2(n_943),
.Y(n_1226)
);

BUFx4f_ASAP7_75t_L g1227 ( 
.A(n_1036),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1009),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1176),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1101),
.B(n_1109),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1106),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1131),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1130),
.A2(n_1202),
.B1(n_1120),
.B2(n_1121),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1110),
.B(n_1214),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1125),
.B(n_1111),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1131),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1211),
.A2(n_1224),
.B1(n_1216),
.B2(n_1113),
.Y(n_1237)
);

CKINVDCx11_ASAP7_75t_R g1238 ( 
.A(n_1126),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1181),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1198),
.A2(n_1108),
.B(n_1141),
.Y(n_1240)
);

BUFx2_ASAP7_75t_R g1241 ( 
.A(n_1140),
.Y(n_1241)
);

CKINVDCx16_ASAP7_75t_R g1242 ( 
.A(n_1149),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1222),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1225),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1129),
.Y(n_1245)
);

CKINVDCx8_ASAP7_75t_R g1246 ( 
.A(n_1209),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1105),
.B(n_1113),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1123),
.B(n_1102),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1201),
.B(n_1118),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1195),
.Y(n_1250)
);

NOR2xp67_ASAP7_75t_SL g1251 ( 
.A(n_1121),
.B(n_1123),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1102),
.B(n_1112),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1160),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1203),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1202),
.A2(n_1153),
.B1(n_1213),
.B2(n_1139),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1116),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1213),
.A2(n_1139),
.B1(n_1226),
.B2(n_1196),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1199),
.B(n_1204),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1180),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1180),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1196),
.A2(n_1226),
.B1(n_1117),
.B2(n_1119),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1101),
.B(n_1109),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1158),
.A2(n_1107),
.B(n_1136),
.Y(n_1263)
);

INVx6_ASAP7_75t_L g1264 ( 
.A(n_1160),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1155),
.A2(n_1197),
.B1(n_1223),
.B2(n_1220),
.Y(n_1265)
);

BUFx12f_ASAP7_75t_L g1266 ( 
.A(n_1157),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1133),
.A2(n_1103),
.B1(n_1119),
.B2(n_1124),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1183),
.B(n_1177),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1137),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1201),
.B(n_1127),
.Y(n_1270)
);

BUFx8_ASAP7_75t_SL g1271 ( 
.A(n_1227),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1221),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1215),
.B(n_1124),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1144),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1207),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1158),
.A2(n_1100),
.B(n_1162),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1208),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1148),
.A2(n_1152),
.B(n_1145),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1147),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1227),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1159),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1128),
.A2(n_1146),
.B1(n_1163),
.B2(n_1210),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1167),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1219),
.A2(n_1165),
.B1(n_1218),
.B2(n_1217),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1156),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1104),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1159),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1166),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1122),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1142),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1174),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1114),
.Y(n_1292)
);

NAND2x1p5_ASAP7_75t_L g1293 ( 
.A(n_1177),
.B(n_1186),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1170),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1132),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1173),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1128),
.A2(n_1154),
.B1(n_1165),
.B2(n_1164),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1168),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1212),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1150),
.Y(n_1300)
);

NAND2x1p5_ASAP7_75t_L g1301 ( 
.A(n_1177),
.B(n_1182),
.Y(n_1301)
);

NAND2x1p5_ASAP7_75t_L g1302 ( 
.A(n_1177),
.B(n_1178),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1145),
.A2(n_1184),
.B(n_1151),
.Y(n_1303)
);

AO21x2_ASAP7_75t_L g1304 ( 
.A1(n_1175),
.A2(n_1172),
.B(n_1185),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1169),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1178),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1143),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1178),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1175),
.A2(n_1172),
.B(n_1171),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1200),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1193),
.Y(n_1311)
);

CKINVDCx11_ASAP7_75t_R g1312 ( 
.A(n_1206),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1134),
.B(n_1135),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1194),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1134),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1188),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1192),
.A2(n_1187),
.B1(n_1228),
.B2(n_1135),
.Y(n_1317)
);

OA21x2_ASAP7_75t_L g1318 ( 
.A1(n_1179),
.A2(n_1189),
.B(n_1171),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1205),
.A2(n_1138),
.B1(n_1161),
.B2(n_1228),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1205),
.A2(n_1135),
.B1(n_1188),
.B2(n_1190),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1188),
.A2(n_1190),
.B1(n_1191),
.B2(n_1205),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1191),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1131),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1130),
.A2(n_1098),
.B1(n_930),
.B2(n_912),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1176),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1115),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1176),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1120),
.A2(n_930),
.B1(n_1130),
.B2(n_1111),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1202),
.A2(n_1098),
.B1(n_930),
.B2(n_632),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1176),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1198),
.A2(n_930),
.B(n_938),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1181),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1176),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1101),
.B(n_1109),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1176),
.Y(n_1335)
);

AO21x1_ASAP7_75t_SL g1336 ( 
.A1(n_1267),
.A2(n_1240),
.B(n_1233),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1258),
.B(n_1247),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1291),
.B(n_1255),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1270),
.B(n_1235),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1281),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1270),
.B(n_1235),
.Y(n_1341)
);

AOI221xp5_ASAP7_75t_L g1342 ( 
.A1(n_1328),
.A2(n_1324),
.B1(n_1331),
.B2(n_1329),
.C(n_1257),
.Y(n_1342)
);

NAND2xp33_ASAP7_75t_SL g1343 ( 
.A(n_1280),
.B(n_1252),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1291),
.B(n_1229),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1281),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1242),
.B(n_1231),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1249),
.B(n_1261),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1229),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1237),
.A2(n_1282),
.B(n_1251),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1249),
.B(n_1234),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1325),
.B(n_1327),
.Y(n_1351)
);

AO21x1_ASAP7_75t_SL g1352 ( 
.A1(n_1273),
.A2(n_1335),
.B(n_1333),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1256),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1256),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1330),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1333),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1259),
.B(n_1260),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1311),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1287),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1272),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1248),
.B(n_1285),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1303),
.B(n_1276),
.Y(n_1362)
);

NAND2x1_ASAP7_75t_L g1363 ( 
.A(n_1322),
.B(n_1318),
.Y(n_1363)
);

INVx4_ASAP7_75t_L g1364 ( 
.A(n_1232),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1275),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1263),
.A2(n_1276),
.B(n_1290),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1309),
.A2(n_1290),
.B(n_1298),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1278),
.B(n_1311),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1238),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1263),
.A2(n_1278),
.B(n_1304),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1309),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1314),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1297),
.B(n_1265),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1268),
.B(n_1293),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1278),
.B(n_1304),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1306),
.A2(n_1308),
.B(n_1316),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_1299),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1301),
.A2(n_1302),
.B(n_1268),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1304),
.B(n_1239),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1245),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1250),
.Y(n_1381)
);

NAND2xp33_ASAP7_75t_SL g1382 ( 
.A(n_1280),
.B(n_1236),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1243),
.B(n_1326),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1300),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1244),
.B(n_1269),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1254),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1318),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1318),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1293),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1286),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1301),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1301),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1268),
.Y(n_1393)
);

NAND2xp33_ASAP7_75t_R g1394 ( 
.A(n_1239),
.B(n_1332),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1279),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1294),
.B(n_1296),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1332),
.B(n_1283),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1368),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1363),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1363),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1371),
.B(n_1393),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1367),
.B(n_1274),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1367),
.B(n_1313),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1367),
.B(n_1313),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1387),
.B(n_1288),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1337),
.B(n_1246),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1362),
.B(n_1321),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1348),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1362),
.B(n_1317),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1388),
.B(n_1320),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1388),
.B(n_1315),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1357),
.B(n_1277),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1357),
.B(n_1305),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1375),
.B(n_1379),
.Y(n_1414)
);

OR2x6_ASAP7_75t_L g1415 ( 
.A(n_1374),
.B(n_1264),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1375),
.B(n_1300),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1366),
.B(n_1284),
.Y(n_1417)
);

NOR2x1_ASAP7_75t_L g1418 ( 
.A(n_1379),
.B(n_1295),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1358),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1376),
.Y(n_1420)
);

NOR2x1_ASAP7_75t_SL g1421 ( 
.A(n_1374),
.B(n_1236),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_R g1422 ( 
.A(n_1369),
.B(n_1246),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1376),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1352),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1370),
.A2(n_1307),
.B(n_1334),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1342),
.A2(n_1230),
.B1(n_1334),
.B2(n_1262),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1339),
.B(n_1319),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1374),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1351),
.B(n_1292),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1376),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1426),
.A2(n_1349),
.B(n_1373),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1405),
.B(n_1340),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1406),
.B(n_1343),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1420),
.Y(n_1434)
);

OAI21xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1418),
.A2(n_1378),
.B(n_1338),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1422),
.B(n_1384),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1426),
.A2(n_1336),
.B1(n_1347),
.B2(n_1338),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1405),
.B(n_1345),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1403),
.B(n_1404),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1405),
.B(n_1353),
.Y(n_1440)
);

NAND3xp33_ASAP7_75t_L g1441 ( 
.A(n_1427),
.B(n_1397),
.C(n_1377),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1412),
.B(n_1354),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1421),
.A2(n_1347),
.B1(n_1336),
.B2(n_1350),
.Y(n_1443)
);

OAI21xp33_ASAP7_75t_L g1444 ( 
.A1(n_1427),
.A2(n_1361),
.B(n_1341),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1409),
.B(n_1397),
.C(n_1359),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1412),
.B(n_1360),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1413),
.B(n_1365),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1409),
.B(n_1394),
.C(n_1385),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1403),
.B(n_1352),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1418),
.B(n_1395),
.C(n_1386),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1429),
.B(n_1346),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1404),
.B(n_1355),
.Y(n_1452)
);

NAND3xp33_ASAP7_75t_L g1453 ( 
.A(n_1407),
.B(n_1395),
.C(n_1386),
.Y(n_1453)
);

AOI21xp33_ASAP7_75t_L g1454 ( 
.A1(n_1407),
.A2(n_1389),
.B(n_1392),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1417),
.B(n_1355),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1417),
.B(n_1356),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1424),
.A2(n_1390),
.B1(n_1289),
.B2(n_1295),
.Y(n_1457)
);

NOR3xp33_ASAP7_75t_L g1458 ( 
.A(n_1399),
.B(n_1382),
.C(n_1364),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1414),
.B(n_1344),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1398),
.Y(n_1460)
);

NOR3xp33_ASAP7_75t_SL g1461 ( 
.A(n_1408),
.B(n_1392),
.C(n_1391),
.Y(n_1461)
);

OAI221xp5_ASAP7_75t_L g1462 ( 
.A1(n_1428),
.A2(n_1310),
.B1(n_1289),
.B2(n_1380),
.C(n_1381),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1411),
.B(n_1356),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1419),
.B(n_1372),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1416),
.B(n_1396),
.C(n_1383),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1416),
.B(n_1238),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1439),
.B(n_1420),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1460),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1439),
.B(n_1420),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1452),
.B(n_1402),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1455),
.B(n_1402),
.Y(n_1471)
);

BUFx2_ASAP7_75t_SL g1472 ( 
.A(n_1436),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1462),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1434),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1463),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1434),
.B(n_1400),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1459),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1449),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1449),
.B(n_1456),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1450),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1456),
.B(n_1423),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1459),
.Y(n_1482)
);

NOR2x1p5_ASAP7_75t_L g1483 ( 
.A(n_1448),
.B(n_1310),
.Y(n_1483)
);

AND2x4_ASAP7_75t_SL g1484 ( 
.A(n_1458),
.B(n_1415),
.Y(n_1484)
);

NAND2xp67_ASAP7_75t_L g1485 ( 
.A(n_1446),
.B(n_1396),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1465),
.B(n_1402),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1464),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1435),
.B(n_1430),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1445),
.B(n_1414),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1465),
.B(n_1414),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1453),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1435),
.B(n_1430),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1453),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1461),
.B(n_1400),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1440),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1480),
.B(n_1441),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1467),
.B(n_1410),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1482),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1467),
.B(n_1410),
.Y(n_1499)
);

OR2x6_ASAP7_75t_L g1500 ( 
.A(n_1472),
.B(n_1415),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1467),
.B(n_1410),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1469),
.B(n_1451),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1489),
.B(n_1432),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1478),
.B(n_1399),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1488),
.B(n_1425),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1482),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1488),
.B(n_1425),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1473),
.B(n_1466),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1478),
.B(n_1476),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1488),
.B(n_1425),
.Y(n_1510)
);

AOI322xp5_ASAP7_75t_L g1511 ( 
.A1(n_1480),
.A2(n_1444),
.A3(n_1437),
.B1(n_1433),
.B2(n_1443),
.C1(n_1431),
.C2(n_1454),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1478),
.B(n_1401),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1494),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1493),
.B(n_1441),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1489),
.B(n_1438),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_L g1516 ( 
.A(n_1493),
.B(n_1448),
.C(n_1444),
.Y(n_1516)
);

NOR3xp33_ASAP7_75t_L g1517 ( 
.A(n_1491),
.B(n_1445),
.C(n_1473),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1477),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1474),
.Y(n_1519)
);

INVxp67_ASAP7_75t_SL g1520 ( 
.A(n_1491),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1477),
.Y(n_1521)
);

NOR2xp67_ASAP7_75t_L g1522 ( 
.A(n_1491),
.B(n_1489),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1486),
.B(n_1447),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1474),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1486),
.B(n_1442),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1494),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1474),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1475),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1481),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1487),
.B(n_1411),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1518),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1514),
.B(n_1490),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1518),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1521),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1525),
.B(n_1490),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1519),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1497),
.B(n_1499),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1521),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1514),
.B(n_1470),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1517),
.B(n_1473),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1509),
.Y(n_1541)
);

NAND2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1513),
.B(n_1494),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1522),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1496),
.B(n_1470),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1497),
.B(n_1478),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1519),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1528),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1517),
.B(n_1485),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1525),
.B(n_1523),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1528),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1498),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1498),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1496),
.B(n_1471),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1506),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1513),
.B(n_1484),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1497),
.B(n_1478),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1508),
.B(n_1472),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1506),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1522),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1499),
.B(n_1479),
.Y(n_1560)
);

INVx1_ASAP7_75t_SL g1561 ( 
.A(n_1526),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1520),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1516),
.B(n_1502),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1523),
.B(n_1485),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1526),
.B(n_1487),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1520),
.Y(n_1566)
);

NAND2x1p5_ASAP7_75t_L g1567 ( 
.A(n_1509),
.B(n_1494),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1530),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1516),
.B(n_1495),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1530),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1499),
.B(n_1501),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1503),
.B(n_1495),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1501),
.B(n_1479),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1537),
.B(n_1509),
.Y(n_1574)
);

AO21x2_ASAP7_75t_L g1575 ( 
.A1(n_1540),
.A2(n_1507),
.B(n_1505),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1569),
.B(n_1501),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1537),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1547),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1571),
.B(n_1502),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1550),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1557),
.A2(n_1483),
.B1(n_1500),
.B2(n_1494),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1571),
.B(n_1502),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1560),
.B(n_1573),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1543),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1563),
.B(n_1532),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1532),
.B(n_1503),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1536),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1560),
.B(n_1509),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1573),
.B(n_1509),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1531),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1533),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1561),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1536),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1542),
.Y(n_1594)
);

AOI21xp33_ASAP7_75t_L g1595 ( 
.A1(n_1548),
.A2(n_1559),
.B(n_1557),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1567),
.B(n_1512),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1542),
.Y(n_1597)
);

INVxp67_ASAP7_75t_SL g1598 ( 
.A(n_1567),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1551),
.B(n_1515),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1562),
.A2(n_1500),
.B(n_1450),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1564),
.A2(n_1483),
.B1(n_1500),
.B2(n_1555),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1566),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1564),
.A2(n_1500),
.B(n_1484),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1555),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1555),
.B(n_1512),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1534),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1538),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1565),
.A2(n_1511),
.B(n_1500),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1552),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1608),
.A2(n_1500),
.B1(n_1544),
.B2(n_1553),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1595),
.B(n_1266),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1592),
.B(n_1565),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1592),
.B(n_1539),
.Y(n_1613)
);

AOI32xp33_ASAP7_75t_L g1614 ( 
.A1(n_1604),
.A2(n_1545),
.A3(n_1556),
.B1(n_1505),
.B2(n_1510),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1576),
.B(n_1549),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1584),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1578),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1578),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1580),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1585),
.B(n_1539),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1604),
.Y(n_1621)
);

OAI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1608),
.A2(n_1544),
.B1(n_1553),
.B2(n_1535),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1576),
.B(n_1572),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1580),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1590),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1590),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1595),
.B(n_1266),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1591),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1585),
.B(n_1554),
.Y(n_1629)
);

AOI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1602),
.A2(n_1558),
.B1(n_1570),
.B2(n_1568),
.C(n_1507),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1602),
.A2(n_1511),
.B(n_1492),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1579),
.B(n_1545),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1579),
.B(n_1556),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1581),
.B(n_1515),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1577),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1635),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1612),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1621),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1617),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1611),
.B(n_1627),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1616),
.B(n_1582),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1613),
.B(n_1582),
.Y(n_1642)
);

AOI222xp33_ASAP7_75t_L g1643 ( 
.A1(n_1622),
.A2(n_1586),
.B1(n_1599),
.B2(n_1598),
.C1(n_1597),
.C2(n_1609),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1618),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1631),
.B(n_1609),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1619),
.B(n_1597),
.Y(n_1646)
);

NOR2xp67_ASAP7_75t_L g1647 ( 
.A(n_1631),
.B(n_1594),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1624),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_R g1649 ( 
.A(n_1620),
.B(n_1601),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1625),
.B(n_1626),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1615),
.B(n_1586),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1628),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1629),
.B(n_1312),
.Y(n_1653)
);

AND2x2_ASAP7_75t_SL g1654 ( 
.A(n_1623),
.B(n_1594),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1630),
.B(n_1591),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1630),
.B(n_1606),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1636),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_L g1658 ( 
.A(n_1643),
.B(n_1610),
.C(n_1634),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1645),
.A2(n_1581),
.B1(n_1601),
.B2(n_1597),
.C(n_1600),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1654),
.Y(n_1660)
);

OAI21xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1647),
.A2(n_1614),
.B(n_1594),
.Y(n_1661)
);

NOR2xp67_ASAP7_75t_L g1662 ( 
.A(n_1638),
.B(n_1594),
.Y(n_1662)
);

NAND4xp25_ASAP7_75t_L g1663 ( 
.A(n_1640),
.B(n_1641),
.C(n_1653),
.D(n_1645),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1650),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1650),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1655),
.A2(n_1600),
.B1(n_1633),
.B2(n_1632),
.C(n_1575),
.Y(n_1666)
);

NOR3xp33_ASAP7_75t_L g1667 ( 
.A(n_1637),
.B(n_1655),
.C(n_1656),
.Y(n_1667)
);

NAND3x2_ASAP7_75t_L g1668 ( 
.A(n_1651),
.B(n_1596),
.C(n_1605),
.Y(n_1668)
);

NAND4xp25_ASAP7_75t_L g1669 ( 
.A(n_1658),
.B(n_1656),
.C(n_1642),
.D(n_1644),
.Y(n_1669)
);

AND5x1_ASAP7_75t_L g1670 ( 
.A(n_1666),
.B(n_1649),
.C(n_1603),
.D(n_1646),
.E(n_1639),
.Y(n_1670)
);

NOR4xp25_ASAP7_75t_L g1671 ( 
.A(n_1663),
.B(n_1652),
.C(n_1648),
.D(n_1606),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1667),
.A2(n_1646),
.B1(n_1577),
.B2(n_1603),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1660),
.B(n_1583),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1659),
.A2(n_1312),
.B1(n_1271),
.B2(n_1241),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1657),
.B(n_1583),
.Y(n_1675)
);

NAND3xp33_ASAP7_75t_SL g1676 ( 
.A(n_1659),
.B(n_1599),
.C(n_1577),
.Y(n_1676)
);

NAND4xp75_ASAP7_75t_L g1677 ( 
.A(n_1661),
.B(n_1596),
.C(n_1605),
.D(n_1607),
.Y(n_1677)
);

NOR3x1_ASAP7_75t_L g1678 ( 
.A(n_1664),
.B(n_1607),
.C(n_1271),
.Y(n_1678)
);

NOR3xp33_ASAP7_75t_L g1679 ( 
.A(n_1674),
.B(n_1665),
.C(n_1662),
.Y(n_1679)
);

AOI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1676),
.A2(n_1668),
.B(n_1593),
.C(n_1587),
.Y(n_1680)
);

OAI211xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1672),
.A2(n_1593),
.B(n_1587),
.C(n_1541),
.Y(n_1681)
);

NOR3xp33_ASAP7_75t_L g1682 ( 
.A(n_1669),
.B(n_1593),
.C(n_1587),
.Y(n_1682)
);

NOR3xp33_ASAP7_75t_L g1683 ( 
.A(n_1677),
.B(n_1675),
.C(n_1673),
.Y(n_1683)
);

AOI221x1_ASAP7_75t_L g1684 ( 
.A1(n_1670),
.A2(n_1541),
.B1(n_1574),
.B2(n_1546),
.C(n_1589),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1682),
.Y(n_1685)
);

NOR2x1_ASAP7_75t_L g1686 ( 
.A(n_1681),
.B(n_1671),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1680),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1683),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1679),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1684),
.Y(n_1690)
);

INVxp33_ASAP7_75t_SL g1691 ( 
.A(n_1689),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1686),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1688),
.A2(n_1678),
.B1(n_1575),
.B2(n_1574),
.C(n_1589),
.Y(n_1693)
);

NAND2x1p5_ASAP7_75t_L g1694 ( 
.A(n_1685),
.B(n_1574),
.Y(n_1694)
);

NOR2x1p5_ASAP7_75t_L g1695 ( 
.A(n_1687),
.B(n_1541),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_L g1696 ( 
.A(n_1695),
.B(n_1687),
.Y(n_1696)
);

NOR3xp33_ASAP7_75t_L g1697 ( 
.A(n_1692),
.B(n_1690),
.C(n_1588),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1694),
.B(n_1575),
.Y(n_1698)
);

XNOR2x1_ASAP7_75t_L g1699 ( 
.A(n_1696),
.B(n_1691),
.Y(n_1699)
);

NOR2x1p5_ASAP7_75t_L g1700 ( 
.A(n_1699),
.B(n_1698),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1700),
.A2(n_1697),
.B1(n_1693),
.B2(n_1574),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1700),
.A2(n_1588),
.B(n_1546),
.Y(n_1702)
);

O2A1O1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1702),
.A2(n_1575),
.B(n_1457),
.C(n_1507),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1701),
.A2(n_1505),
.B1(n_1510),
.B2(n_1504),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1704),
.B(n_1519),
.Y(n_1705)
);

INVxp67_ASAP7_75t_SL g1706 ( 
.A(n_1703),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1706),
.A2(n_1705),
.B(n_1529),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1510),
.B1(n_1504),
.B2(n_1527),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1708),
.A2(n_1527),
.B1(n_1524),
.B2(n_1504),
.C(n_1468),
.Y(n_1709)
);

AOI211xp5_ASAP7_75t_L g1710 ( 
.A1(n_1709),
.A2(n_1236),
.B(n_1323),
.C(n_1253),
.Y(n_1710)
);


endmodule