module fake_jpeg_26388_n_412 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_412);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_412;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_11),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_7),
.B(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_41),
.B(n_42),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_43),
.B(n_50),
.Y(n_120)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_7),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_58),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_55),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx2_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_27),
.B(n_6),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_65),
.Y(n_118)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_72),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_6),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_68),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_31),
.Y(n_70)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx11_ASAP7_75t_SL g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_9),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_40),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_26),
.Y(n_99)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_31),
.B(n_9),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_37),
.B1(n_20),
.B2(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_83),
.A2(n_86),
.B1(n_94),
.B2(n_98),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_37),
.B1(n_23),
.B2(n_30),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_5),
.B(n_13),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_50),
.B(n_58),
.C(n_42),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_37),
.B1(n_30),
.B2(n_18),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_17),
.B1(n_18),
.B2(n_15),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_99),
.B(n_54),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_52),
.A2(n_17),
.B1(n_28),
.B2(n_22),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_107),
.B1(n_59),
.B2(n_76),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_39),
.B1(n_28),
.B2(n_22),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_105),
.A2(n_109),
.B1(n_47),
.B2(n_72),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_28),
.B1(n_22),
.B2(n_15),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_45),
.A2(n_39),
.B1(n_15),
.B2(n_29),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_60),
.B(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_39),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_66),
.A2(n_33),
.B1(n_31),
.B2(n_26),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_71),
.B1(n_57),
.B2(n_44),
.Y(n_152)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

NAND2x1_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_77),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_131),
.B(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_130),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_41),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_141),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_81),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_133),
.B(n_139),
.Y(n_190)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

BUFx2_ASAP7_75t_SL g174 ( 
.A(n_135),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_136),
.B(n_158),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_137),
.Y(n_206)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_26),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_70),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_70),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_156),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_26),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_144),
.Y(n_191)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_148),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_111),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_151),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_63),
.B1(n_33),
.B2(n_2),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_150),
.A2(n_164),
.B1(n_95),
.B2(n_160),
.Y(n_194)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_104),
.B1(n_93),
.B2(n_110),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_111),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_49),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_92),
.A2(n_78),
.B1(n_91),
.B2(n_90),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_165),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_14),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_159),
.B(n_162),
.Y(n_195)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_118),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_163),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_115),
.A2(n_14),
.B1(n_13),
.B2(n_2),
.Y(n_164)
);

OR2x2_ASAP7_75t_SL g166 ( 
.A(n_96),
.B(n_84),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_46),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_96),
.C(n_84),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_178),
.C(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_172),
.B(n_181),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_92),
.B1(n_84),
.B2(n_110),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_176),
.A2(n_161),
.B1(n_131),
.B2(n_102),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_107),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_129),
.B(n_93),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

NAND2xp33_ASAP7_75t_SL g182 ( 
.A(n_127),
.B(n_49),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_182),
.A2(n_183),
.B(n_203),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_100),
.B(n_106),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_46),
.Y(n_221)
);

OAI32xp33_ASAP7_75t_L g186 ( 
.A1(n_129),
.A2(n_106),
.A3(n_100),
.B1(n_90),
.B2(n_95),
.Y(n_186)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_145),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_144),
.B1(n_151),
.B2(n_149),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_49),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_54),
.C(n_126),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_116),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_207),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_46),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_201),
.B(n_207),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_209),
.A2(n_221),
.B(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_157),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_223),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_152),
.B1(n_157),
.B2(n_138),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_213),
.A2(n_217),
.B1(n_226),
.B2(n_228),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_214),
.A2(n_215),
.B1(n_218),
.B2(n_232),
.Y(n_274)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_167),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_222),
.Y(n_252)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_220),
.B(n_241),
.Y(n_276)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_124),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_102),
.B1(n_122),
.B2(n_117),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_225),
.B1(n_236),
.B2(n_169),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_122),
.B1(n_117),
.B2(n_134),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_176),
.A2(n_101),
.B1(n_71),
.B2(n_69),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_227),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_192),
.A2(n_101),
.B1(n_67),
.B2(n_162),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_172),
.A2(n_158),
.B1(n_136),
.B2(n_97),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_169),
.B1(n_197),
.B2(n_170),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_200),
.C(n_202),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_14),
.B(n_13),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_180),
.B(n_54),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_238),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_147),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_235),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_146),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_179),
.A2(n_181),
.B1(n_184),
.B2(n_203),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_239),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_178),
.B(n_0),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_146),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_189),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_243),
.Y(n_270)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

NAND2xp33_ASAP7_75t_SL g244 ( 
.A(n_182),
.B(n_125),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_244),
.A2(n_195),
.B(n_196),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_208),
.C(n_233),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_248),
.A2(n_55),
.B1(n_44),
.B2(n_2),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_227),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_268),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_209),
.A2(n_183),
.B(n_193),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_261),
.B(n_266),
.Y(n_285)
);

OAI21x1_ASAP7_75t_R g255 ( 
.A1(n_215),
.A2(n_173),
.B(n_197),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_255),
.A2(n_262),
.B(n_3),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_212),
.A2(n_239),
.B1(n_211),
.B2(n_210),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_256),
.A2(n_260),
.B1(n_263),
.B2(n_265),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_215),
.B1(n_243),
.B2(n_218),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_212),
.A2(n_193),
.B1(n_168),
.B2(n_170),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_210),
.A2(n_171),
.B(n_135),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_236),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_213),
.A2(n_196),
.B1(n_175),
.B2(n_204),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_221),
.B(n_244),
.Y(n_266)
);

A2O1A1O1Ixp25_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_126),
.B(n_175),
.C(n_56),
.D(n_51),
.Y(n_267)
);

XOR2x1_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_226),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_219),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_237),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_272),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_221),
.A2(n_135),
.B(n_204),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_271),
.A2(n_10),
.B(n_11),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_229),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_275),
.Y(n_290)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_245),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_187),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_279),
.A2(n_282),
.B1(n_303),
.B2(n_305),
.Y(n_312)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_288),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_281),
.A2(n_297),
.B1(n_267),
.B2(n_253),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_258),
.A2(n_217),
.B1(n_230),
.B2(n_242),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

AO22x1_ASAP7_75t_SL g284 ( 
.A1(n_258),
.A2(n_231),
.B1(n_238),
.B2(n_216),
.Y(n_284)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_284),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_289),
.C(n_292),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_208),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_302),
.Y(n_323)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_247),
.B(n_222),
.C(n_232),
.Y(n_289)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_247),
.B(n_125),
.C(n_187),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_254),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_296),
.Y(n_324)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_299),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_55),
.C(n_5),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_264),
.C(n_261),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_260),
.B(n_266),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_246),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_306),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_246),
.A2(n_1),
.B1(n_4),
.B2(n_10),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_294),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_307),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_263),
.B1(n_256),
.B2(n_272),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_313),
.A2(n_318),
.B1(n_319),
.B2(n_296),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_259),
.B1(n_273),
.B2(n_274),
.Y(n_314)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_314),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_291),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_317),
.B(n_330),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_281),
.A2(n_265),
.B1(n_248),
.B2(n_277),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_298),
.A2(n_275),
.B1(n_250),
.B2(n_249),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_300),
.A2(n_259),
.B1(n_257),
.B2(n_253),
.Y(n_320)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_320),
.Y(n_335)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_322),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_297),
.A2(n_270),
.B1(n_276),
.B2(n_249),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_327),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_290),
.A2(n_276),
.B1(n_254),
.B2(n_267),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_315),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_289),
.Y(n_329)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_329),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_287),
.C(n_286),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_331),
.B(n_340),
.C(n_350),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_316),
.A2(n_285),
.B(n_295),
.Y(n_333)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_333),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_334),
.B(n_348),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_323),
.B(n_285),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_341),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_323),
.C(n_292),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_302),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_344),
.Y(n_363)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_309),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_278),
.Y(n_345)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_345),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_303),
.Y(n_347)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_347),
.Y(n_357)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_319),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_284),
.C(n_304),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_332),
.A2(n_316),
.B1(n_338),
.B2(n_342),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_354),
.A2(n_335),
.B1(n_332),
.B2(n_308),
.Y(n_370)
);

AO221x1_ASAP7_75t_L g355 ( 
.A1(n_342),
.A2(n_255),
.B1(n_344),
.B2(n_343),
.C(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

AOI322xp5_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_312),
.A3(n_314),
.B1(n_318),
.B2(n_313),
.C1(n_320),
.C2(n_251),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_338),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_311),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_359),
.A2(n_333),
.B(n_350),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_311),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_365),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_339),
.B(n_301),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_366),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_310),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_339),
.B(n_334),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_341),
.C(n_348),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_369),
.C(n_351),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_364),
.B(n_365),
.C(n_360),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_370),
.A2(n_312),
.B1(n_337),
.B2(n_308),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_363),
.Y(n_371)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_371),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_375),
.C(n_374),
.Y(n_382)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_361),
.B(n_336),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_363),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_378),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_347),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_379),
.B(n_381),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_335),
.C(n_361),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_382),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_368),
.A2(n_351),
.B1(n_359),
.B2(n_310),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_377),
.A2(n_357),
.B1(n_352),
.B2(n_359),
.Y(n_383)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_383),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_356),
.C(n_357),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_385),
.Y(n_396)
);

BUFx24_ASAP7_75t_SL g385 ( 
.A(n_372),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_388),
.A2(n_389),
.B1(n_305),
.B2(n_371),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_384),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_391),
.B(n_393),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_387),
.A2(n_337),
.B(n_372),
.Y(n_392)
);

AOI21xp33_ASAP7_75t_L g402 ( 
.A1(n_392),
.A2(n_325),
.B(n_269),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_375),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_397),
.A2(n_325),
.B(n_251),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_396),
.B(n_386),
.Y(n_398)
);

NOR3xp33_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_399),
.C(n_400),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_395),
.B(n_391),
.Y(n_399)
);

AOI31xp33_ASAP7_75t_L g400 ( 
.A1(n_390),
.A2(n_284),
.A3(n_306),
.B(n_271),
.Y(n_400)
);

OAI31xp33_ASAP7_75t_SL g405 ( 
.A1(n_401),
.A2(n_390),
.A3(n_394),
.B(n_393),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_402),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_405),
.A2(n_403),
.B(n_255),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_407),
.A2(n_408),
.B(n_406),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_404),
.A2(n_268),
.B(n_299),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g410 ( 
.A(n_409),
.Y(n_410)
);

OAI321xp33_ASAP7_75t_L g411 ( 
.A1(n_410),
.A2(n_1),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C(n_408),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_411),
.B(n_10),
.Y(n_412)
);


endmodule